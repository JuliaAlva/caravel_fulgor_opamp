  X �     "�     " user_project_wrapper >A�7KƧ�9D�/��ZT �     "�     " "sky130_fd_pr__pfet_01v8_YT7TV5    �   ,�����������  D  	  D  	����������      A   ,���  N���    `    `  N���  N      A   ,��������������  `����  `�����������      A  , ,���  ����  �  ^  �  ^  ����  �      A  , ,���������  ����L  ����L���������      A  , ,  ����  �  �  ^  �  ^���  ����      A  , ,������g������  ^���  ^���g������g      ^   ,���#  ����#  �  �  �  �  ����#  �      ^   ,���#���}���#���/  ����/  ����}���#���}      ]  , ,���%  r���%    �    �  r���%  r      ]  , ,���%������%  r����  r����������%���      ]  , ,  7���  7  r  �  r  ����  7���      ]  , ,���%�������%���  ����  ��������%����      B   ,���[  ����[  �   �  �   �  ����[  �      B   ,���j  ����j  �   �  �   �  ����j  �      B   ,���[   i���[  �   �  �   �   i���[   i      B   ,���[���M���[����   �����   ����M���[���M      B   ,���j���_���j���M   ����M   ����_���j���_      B   ,���[������[���_   ����_   �������[���      B   ,  /  �  /  �  y  �  y  �  /  �      B   ,  }  �  }  �  �  �  �  �  }  �      B   ,  �  �  �  �    �    �  �  �      B   ,    �    �  c  �  c  �    �      B   ,  g  �  g  �  �  �  �  �  g  �      B   ,  �  �  �  �  �  �  �  �  �  �      B   ,    �    �  M  �  M  �    �      B   ,  �  �  �  �  �  �  �  �  �  �      B   ,  �  �  �  �  �  �  �  �  �  �      B   ,    �    �  2  �  2  �    �      B   ,  T  �  T  �  �  �  �  �  T  �      B   ,  �  �  �  �  	�  �  	�  �  �  �      B   ,  
�  �  
�  �    �    �  
�  �      B   ,  >  �  >  �  j  �  j  �  >  �      B   ,  �  �  �  �  �  �  �  �  �  �      B   ,  �  �  �  �    �    �  �  �      B   ,  (  �  (  �  T  �  T  �  (  �      B   ,  v  �  v  �  �  �  �  �  v  �      B   ,  �  �  �  �  �  �  �  �  �  �      B   ,    �    �  >  �  >  �    �      B   ,  �  �  �  �  A  �  A  �  �  �      B   ,  �   i  �  �  �  �  �   i  �   i      B   ,  �   i  �  �  A  �  A   i  �   i      B   ,  E   i  E  �  �  �  �   i  E   i      B   ,  �   i  �  �  	�  �  	�   i  �   i      B   ,  
�   i  
�  �  +  �  +   i  
�   i      B   ,  /   i  /  �  y  �  y   i  /   i      B   ,  }   i  }  �  �  �  �   i  }   i      B   ,  �   i  �  �    �     i  �   i      B   ,     i    �  c  �  c   i     i      B   ,  g   i  g  �  �  �  �   i  g   i      B   ,  �   i  �  �  �  �  �   i  �   i      B   ,     i    �  M  �  M   i     i      B   ,  E  �  E  �  �  �  �  �  E  �      B   ,  �  �  �  �  	�  �  	�  �  �  �      B   ,  
�  �  
�  �  +  �  +  �  
�  �      B   ,���  ����  �����  �����  ����  �      B   ,����  �����  ����  ����  �����  �      B   ,���#  ����#  ����m  ����m  ����#  �      B   ,���q  ����q  �����  �����  ����q  �      B   ,����  �����  ����	  ����	  �����  �      B   ,���  ����  ����W  ����W  ����  �      B   ,���  ����  �����  �����  ����  �      B   ,����  �����  �����  �����  �����  �      B   ,���   i���  �����  �����   i���   i      B   ,���   i���  ����K  ����K   i���   i      B   ,���O   i���O  ����  ����   i���O   i      B   ,���   i���  �����  �����   i���   i      B   ,����   i����  ����5  ����5   i����   i      B   ,���9   i���9  �����  �����   i���9   i      B   ,���   i���  �����  �����   i���   i      B   ,����   i����  ����  ����   i����   i      B   ,���#   i���#  ����m  ����m   i���#   i      B   ,���q   i���q  �����  �����   i���q   i      B   ,����   i����  ����	  ����	   i����   i      B   ,���   i���  ����W  ����W   i���   i      B   ,���  ����  ����<  ����<  ����  �      B   ,���^  ����^  ����  ����  ����^  �      B   ,���  ����  �����  �����  ����  �      B   ,����  �����  ����&  ����&  �����  �      B   ,���H  ����H  ����t  ����t  ����H  �      B   ,���  ����  �����  �����  ����  �      B   ,����  �����  ����  ����  �����  �      B   ,���2  ����2  ����^  ����^  ����2  �      B   ,����  �����  �����  �����  �����  �      B   ,����  �����  �����  �����  �����  �      B   ,���  ����  ����H  ����H  ����  �      B   ,���  ����  ����K  ����K  ����  �      B   ,���O  ����O  ����  ����  ����O  �      B   ,���  ����  �����  �����  ����  �      B   ,����  �����  ����5  ����5  �����  �      B   ,���9  ����9  �����  �����  ����9  �      B   ,������M����������������������M������M      B   ,�������M�����������5�������5���M�������M      B   ,���9���M���9�������������������M���9���M      B   ,������M����������������������M������M      B   ,�������M���������������������M�������M      B   ,���#���M���#�������m�������m���M���#���M      B   ,���q���M���q�������������������M���q���M      B   ,�������M�����������	�������	���M�������M      B   ,������M����������W�������W���M������M      B   ,������M����������������������M������M      B   ,�������_�������M�������M�������_�������_      B   ,������_������M���<���M���<���_������_      B   ,���^���_���^���M������M������_���^���_      B   ,������_������M�������M�������_������_      B   ,�������_�������M���&���M���&���_�������_      B   ,���H���_���H���M���t���M���t���_���H���_      B   ,������_������M�������M�������_������_      B   ,�������_�������M������M������_�������_      B   ,���2���_���2���M���^���M���^���_���2���_      B   ,�������_�������M�������M�������_�������_      B   ,�������_�������M�������M�������_�������_      B   ,������_������M���H���M���H���_������_      B   ,������M����������K�������K���M������M      B   ,������������_�������_�������������      B   ,������������_���K���_���K���������      B   ,���O������O���_������_���������O���      B   ,������������_�������_�������������      B   ,��������������_���5���_���5����������      B   ,���9������9���_�������_����������9���      B   ,������������_�������_�������������      B   ,��������������_������_�������������      B   ,���#������#���_���m���_���m������#���      B   ,���q������q���_�������_����������q���      B   ,��������������_���	���_���	����������      B   ,������������_���W���_���W���������      B   ,���O���M���O�����������������M���O���M      B   ,  ���_  ���M  2���M  2���_  ���_      B   ,  T���_  T���M  ����M  ����_  T���_      B   ,  ����_  ����M  	����M  	����_  ����_      B   ,  
����_  
����M  ���M  ���_  
����_      B   ,  >���_  >���M  j���M  j���_  >���_      B   ,  ����_  ����M  ����M  ����_  ����_      B   ,  ����_  ����M  ���M  ���_  ����_      B   ,  (���_  (���M  T���M  T���_  (���_      B   ,  v���_  v���M  ����M  ����_  v���_      B   ,  ����_  ����M  ����M  ����_  ����_      B   ,  ���_  ���M  >���M  >���_  ���_      B   ,  ����M  �����  A����  A���M  ����M      B   ,  E���M  E����  �����  ����M  E���M      B   ,  ����M  �����  	�����  	����M  ����M      B   ,  
����M  
�����  +����  +���M  
����M      B   ,  /���M  /����  y����  y���M  /���M      B   ,  }���M  }����  �����  ����M  }���M      B   ,  ����M  �����  ����  ���M  ����M      B   ,  ���M  ����  c����  c���M  ���M      B   ,  g���M  g����  �����  ����M  g���M      B   ,  ����M  �����  �����  ����M  ����M      B   ,  ���M  ����  M����  M���M  ���M      B   ,  ����M  �����  �����  ����M  ����M      B   ,  ����_  ����M  ����M  ����_  ����_      B   ,  ����  ����_  ����_  ����  ����      B   ,  ����  ����_  A���_  A���  ����      B   ,  E���  E���_  ����_  ����  E���      B   ,  ����  ����_  	����_  	����  ����      B   ,  
����  
����_  +���_  +���  
����      B   ,  /���  /���_  y���_  y���  /���      B   ,  }���  }���_  ����_  ����  }���      B   ,  ����  ����_  ���_  ���  ����      B   ,  ���  ���_  c���_  c���  ���      B   ,  g���  g���_  ����_  ����  g���      B   ,  ����  ����_  ����_  ����  ����      B   ,  ���  ���_  M���_  M���  ���      B  , ,����   �����  c   U  c   U   �����   �      B  , ,���������������G   U���G   U������������      B  , ,   �     �  	)  |  	)  |     �        B  , ,          	)  �  	)  �             B  , ,  n    n  	)    	)      n        B  , ,  �    �  	)  f  	)  f    �        B  , ,  

    

  	)  
�  	)  
�    

        B  , ,  X    X  	)    	)      X        B  , ,  �    �  	)  P  	)  P    �        B  , ,  �    �  	)  �  	)  �    �        B  , ,  B    B  	)  �  	)  �    B        B  , ,  �    �  	)  :  	)  :    �        B  , ,  �    �  	)  �  	)  �    �        B  , ,  ,    ,  	)  �  	)  �    ,        B  , ,  z    z  	)  $  	)  $    z        B  , ,  �  M  �  �  ^  �  ^  M  �  M      B  , ,  �  {  �  %  :  %  :  {  �  {      B  , ,  �  {  �  %  �  %  �  {  �  {      B  , ,  ,  {  ,  %  �  %  �  {  ,  {      B  , ,  z  {  z  %  $  %  $  {  z  {      B  , ,  �  I  �  �  ^  �  ^  I  �  I      B  , ,  �  '  �  �  �  �  �  '  �  '      B  , ,  B  '  B  �  �  �  �  '  B  '      B  , ,  �  '  �  �  :  �  :  '  �  '      B  , ,  �  '  �  �  �  �  �  '  �  '      B  , ,  ,  '  ,  �  �  �  �  '  ,  '      B  , ,  z  '  z  �  $  �  $  '  z  '      B  , ,  �  
�  �  �  ^  �  ^  
�  �  
�      B  , ,  �  	�  �  
}  �  
}  �  	�  �  	�      B  , ,  B  	�  B  
}  �  
}  �  	�  B  	�      B  , ,  �  	�  �  
}  :  
}  :  	�  �  	�      B  , ,  �  	�  �  
}  �  
}  �  	�  �  	�      B  , ,  ,  	�  ,  
}  �  
}  �  	�  ,  	�      B  , ,  z  	�  z  
}  $  
}  $  	�  z  	�      B  , ,  �  	�  �  
K  ^  
K  ^  	�  �  	�      B  , ,  E  �  E  �  �  �  �  �  E  �      B  , ,  �  �  �  �  C  �  C  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  A  �  A  �  �  �  �  �  A  �      B  , ,  �  �  �  �  ?  �  ?  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  =  �  =  �  �  �  �  �  =  �      B  , ,  �  �  �  �  ;  �  ;  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  9  �  9  �  �  �  �  �  9  �      B  , ,  �  �  �  �  ^  �  ^  �  �  �      B  , ,  �  �  �  G  ^  G  ^  �  �  �      B  , ,  �  {  �  %  �  %  �  {  �  {      B  , ,  B  {  B  %  �  %  �  {  B  {      B  , ,     {     %  �  %  �  {     {      B  , ,  n  {  n  %    %    {  n  {      B  , ,  �  {  �  %  f  %  f  {  �  {      B  , ,   �  	�   �  
}  |  
}  |  	�   �  	�      B  , ,     	�     
}  �  
}  �  	�     	�      B  , ,  n  	�  n  
}    
}    	�  n  	�      B  , ,  �  	�  �  
}  f  
}  f  	�  �  	�      B  , ,  

  	�  

  
}  
�  
}  
�  	�  

  	�      B  , ,  X  	�  X  
}    
}    	�  X  	�      B  , ,  �  	�  �  
}  P  
}  P  	�  �  	�      B  , ,  

  {  

  %  
�  %  
�  {  

  {      B  , ,  X  {  X  %    %    {  X  {      B  , ,  �  {  �  %  P  %  P  {  �  {      B  , ,  �  �  �  �  O  �  O  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  M  �  M  �  �  �  �  �  M  �      B  , ,  	�  �  	�  �  
K  �  
K  �  	�  �      B  , ,  
�  �  
�  �  �  �  �  �  
�  �      B  , ,  I  �  I  �  �  �  �  �  I  �      B  , ,  �  �  �  �  G  �  G  �  �  �      B  , ,   �  '   �  �  |  �  |  '   �  '      B  , ,     '     �  �  �  �  '     '      B  , ,  n  '  n  �    �    '  n  '      B  , ,  �  '  �  �  f  �  f  '  �  '      B  , ,  

  '  

  �  
�  �  
�  '  

  '      B  , ,  X  '  X  �    �    '  X  '      B  , ,  �  '  �  �  P  �  P  '  �  '      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  Q  �  Q  �  �  �  �  �  Q  �      B  , ,   �  {   �  %  |  %  |  {   �  {      B  , ,   U  �   U  �   �  �   �  �   U  �      B  , ,  �  �  �  �  S  �  S  �  �  �      B  , ,  n  +  n  �    �    +  n  +      B  , ,  �  +  �  �  f  �  f  +  �  +      B  , ,  

  +  

  �  
�  �  
�  +  

  +      B  , ,  X  +  X  �    �    +  X  +      B  , ,  �  +  �  �  P  �  P  +  �  +      B  , ,   �  �   �  �  |  �  |  �   �  �      B  , ,     �     �  �  �  �  �     �      B  , ,  n  �  n  �    �    �  n  �      B  , ,  �  �  �  �  f  �  f  �  �  �      B  , ,  

  �  

  �  
�  �  
�  �  

  �      B  , ,  X  �  X  �    �    �  X  �      B  , ,  �  �  �  �  P  �  P  �  �  �      B  , ,   �  �   �  -  |  -  |  �   �  �      B  , ,     �     -  �  -  �  �     �      B  , ,  n  �  n  -    -    �  n  �      B  , ,  �  �  �  -  f  -  f  �  �  �      B  , ,  

  �  

  -  
�  -  
�  �  

  �      B  , ,  X  �  X  -    -    �  X  �      B  , ,  �  �  �  -  P  -  P  �  �  �      B  , ,   �  /   �  �  |  �  |  /   �  /      B  , ,     /     �  �  �  �  /     /      B  , ,  n  /  n  �    �    /  n  /      B  , ,  �  /  �  �  f  �  f  /  �  /      B  , ,  

  /  

  �  
�  �  
�  /  

  /      B  , ,  X  /  X  �    �    /  X  /      B  , ,  �  /  �  �  P  �  P  /  �  /      B  , ,   �  +   �  �  |  �  |  +   �  +      B  , ,  �   �  �  c  �  c  �   �  �   �      B  , ,  G   �  G  c  �  c  �   �  G   �      B  , ,  �   �  �  c  ?  c  ?   �  �   �      B  , ,  �   �  �  c  	�  c  	�   �  �   �      B  , ,  1   �  1  c  �  c  �   �  1   �      B  , ,     �    c  )  c  )   �     �      B  , ,     +     �  �  �  �  +     +      B  , ,  B  �  B  -  �  -  �  �  B  �      B  , ,  �  �  �  -  :  -  :  �  �  �      B  , ,  �  �  �  -  �  -  �  �  �  �      B  , ,  ,  �  ,  -  �  -  �  �  ,  �      B  , ,  z  �  z  -  $  -  $  �  z  �      B  , ,  �  Q  �  �  ^  �  ^  Q  �  Q      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  B  �  B  �  �  �  �  �  B  �      B  , ,  �  �  �  �  :  �  :  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  ,  �  ,  �  �  �  �  �  ,  �      B  , ,  z  �  z  �  $  �  $  �  z  �      B  , ,  �  �  �  O  ^  O  ^  �  �  �      B  , ,  �  /  �  �  �  �  �  /  �  /      B  , ,  B  /  B  �  �  �  �  /  B  /      B  , ,  �  /  �  �  :  �  :  /  �  /      B  , ,  �  /  �  �  �  �  �  /  �  /      B  , ,  ,  /  ,  �  �  �  �  /  ,  /      B  , ,  z  /  z  �  $  �  $  /  z  /      B  , ,  �  �  �  �  ^  �  ^  �  �  �      B  , ,  �  �  �  S  ^  S  ^  �  �  �      B  , ,  �  +  �  �  �  �  �  +  �  +      B  , ,  B  +  B  �  �  �  �  +  B  +      B  , ,  �  +  �  �  :  �  :  +  �  +      B  , ,  �  +  �  �  �  �  �  +  �  +      B  , ,  ,  +  ,  �  �  �  �  +  ,  +      B  , ,  z  +  z  �  $  �  $  +  z  +      B  , ,  �  �  �  �  ^  �  ^  �  �  �      B  , ,  �   �  �  c  w  c  w   �  �   �      B  , ,     �    c  �  c  �   �     �      B  , ,  i   �  i  c    c     �  i   �      B  , ,  �   �  �  c  a  c  a   �  �   �      B  , ,     �    c  �  c  �   �     �      B  , ,  S   �  S  c  �  c  �   �  S   �      B  , ,  �   U  �   �  ^   �  ^   U  �   U      B  , ,  �  �  �  -  �  -  �  �  �  �      B  , ,���  M���  ����L  ����L  M���  M      B  , ,����  ����  	)���  	)���  ����        B  , ,���*  ���*  	)����  	)����  ���*        B  , ,���x  ���x  	)���"  	)���"  ���x        B  , ,����  ����  	)���p  	)���p  ����        B  , ,���  ���  	)���  	)���  ���        B  , ,���b  ���b  	)���  	)���  ���b        B  , ,���  ���  	)���Z  	)���Z  ���        B  , ,����  ����  	)���  	)���  ����        B  , ,���L  ���L  	)����  	)����  ���L        B  , ,����  ����  	)���D  	)���D  ����        B  , ,����  ����  	)����  	)����  ����        B  , ,���6  ���6  	)����  	)����  ���6        B  , ,����  ����  	)���.  	)���.  ����        B  , ,���Y  ����Y  ����  ����  ����Y  �      B  , ,����  �����  ����W  ����W  �����  �      B  , ,���  ����  �����  �����  ����  �      B  , ,���  	����  
}���Z  
}���Z  	����  	�      B  , ,����  	�����  
}���  
}���  	�����  	�      B  , ,���L  	����L  
}����  
}����  	����L  	�      B  , ,����  	�����  
}���D  
}���D  	�����  	�      B  , ,����  	�����  
}����  
}����  	�����  	�      B  , ,���6  	����6  
}����  
}����  	����6  	�      B  , ,����  	�����  
}���.  
}���.  	�����  	�      B  , ,���  {���  %���Z  %���Z  {���  {      B  , ,����  {����  %���  %���  {����  {      B  , ,���L  {���L  %����  %����  {���L  {      B  , ,����  {����  %���D  %���D  {����  {      B  , ,����  {����  %����  %����  {����  {      B  , ,���6  {���6  %����  %����  {���6  {      B  , ,����  {����  %���.  %���.  {����  {      B  , ,���  ����  ����  ����  ����  �      B  , ,���a  ����a  ����  ����  ����a  �      B  , ,����  �����  ����_  ����_  �����  �      B  , ,���	  ����	  �����  �����  ����	  �      B  , ,���  '���  ����Z  ����Z  '���  '      B  , ,����  '����  ����  ����  '����  '      B  , ,���L  '���L  �����  �����  '���L  '      B  , ,����  '����  ����D  ����D  '����  '      B  , ,����  '����  �����  �����  '����  '      B  , ,���6  '���6  �����  �����  '���6  '      B  , ,����  '����  ����.  ����.  '����  '      B  , ,���]  ����]  ����  ����  ����]  �      B  , ,����  �����  ����[  ����[  �����  �      B  , ,���  ����  �����  �����  ����  �      B  , ,���e  ����e  ����  ����  ����e  �      B  , ,���  ����  ����c  ����c  ����  �      B  , ,���  {���  %���  %���  {���  {      B  , ,���b  {���b  %���  %���  {���b  {      B  , ,���  ����  ����L  ����L  ����  �      B  , ,���  ����  �����  �����  ����  �      B  , ,���  ����  G���L  G���L  ����  �      B  , ,���q  ����q  ����  ����  ����q  �      B  , ,���  I���  ����L  ����L  I���  I      B  , ,����  {����  %���  %���  {����  {      B  , ,���*  {���*  %����  %����  {���*  {      B  , ,����  �����  ����o  ����o  �����  �      B  , ,���  ����  �����  �����  ����  �      B  , ,���m  ����m  ����  ����  ����m  �      B  , ,����  �����  ����k  ����k  �����  �      B  , ,���x  {���x  %���"  %���"  {���x  {      B  , ,���  	����  
K���L  
K���L  	����  	�      B  , ,����  	�����  
}���  
}���  	�����  	�      B  , ,���*  	����*  
}����  
}����  	����*  	�      B  , ,���x  	����x  
}���"  
}���"  	����x  	�      B  , ,����  	�����  
}���p  
}���p  	�����  	�      B  , ,���  	����  
}���  
}���  	����  	�      B  , ,���b  	����b  
}���  
}���  	����b  	�      B  , ,���b  '���b  ����  ����  '���b  '      B  , ,���  
����  ����L  ����L  
����  
�      B  , ,����  '����  ����  ����  '����  '      B  , ,���*  '���*  �����  �����  '���*  '      B  , ,���x  '���x  ����"  ����"  '���x  '      B  , ,����  '����  ����p  ����p  '����  '      B  , ,���  ����  ����  ����  ����  �      B  , ,���i  ����i  ����  ����  ����i  �      B  , ,���  ����  ����g  ����g  ����  �      B  , ,���  ����  ����  ����  ����  �      B  , ,���  '���  ����  ����  '���  '      B  , ,����  {����  %���p  %���p  {����  {      B  , ,���*  ����*  -����  -����  ����*  �      B  , ,���x  ����x  -���"  -���"  ����x  �      B  , ,����  �����  -���p  -���p  �����  �      B  , ,���  ����  -���  -���  ����  �      B  , ,���b  ����b  -���  -���  ����b  �      B  , ,���  ����  ����L  ����L  ����  �      B  , ,����  +����  ����  ����  +����  +      B  , ,���*  +���*  �����  �����  +���*  +      B  , ,���x  +���x  ����"  ����"  +���x  +      B  , ,����  +����  ����p  ����p  +����  +      B  , ,���  +���  ����  ����  +���  +      B  , ,���b  +���b  ����  ����  +���b  +      B  , ,���  ����  S���L  S���L  ����  �      B  , ,���  ����  O���L  O���L  ����  �      B  , ,���   U���   ����L   ����L   U���   U      B  , ,���   ����  c���  c���   ����   �      B  , ,���Q   ����Q  c����  c����   ����Q   �      B  , ,���   ����  c���I  c���I   ����   �      B  , ,����   �����  c���  c���   �����   �      B  , ,���;   ����;  c����  c����   ����;   �      B  , ,���   ����  c���3  c���3   ����   �      B  , ,����  �����  ����  ����  �����  �      B  , ,���*  ����*  �����  �����  ����*  �      B  , ,���x  ����x  ����"  ����"  ����x  �      B  , ,����  �����  ����p  ����p  �����  �      B  , ,���  ����  ����  ����  ����  �      B  , ,���b  ����b  ����  ����  ����b  �      B  , ,���  ����  ����L  ����L  ����  �      B  , ,����  /����  ����  ����  /����  /      B  , ,���*  /���*  �����  �����  /���*  /      B  , ,���x  /���x  ����"  ����"  /���x  /      B  , ,����  /����  ����p  ����p  /����  /      B  , ,���  /���  ����  ����  /���  /      B  , ,���b  /���b  ����  ����  /���b  /      B  , ,���  Q���  ����L  ����L  Q���  Q      B  , ,����  �����  -���  -���  �����  �      B  , ,����  +����  ����D  ����D  +����  +      B  , ,����  +����  �����  �����  +����  +      B  , ,���6  +���6  �����  �����  +���6  +      B  , ,����  +����  ����.  ����.  +����  +      B  , ,���  ����  -���Z  -���Z  ����  �      B  , ,����  �����  -���  -���  �����  �      B  , ,���L  ����L  -����  -����  ����L  �      B  , ,����  �����  -���D  -���D  �����  �      B  , ,����  �����  -����  -����  �����  �      B  , ,���6  ����6  -����  -����  ����6  �      B  , ,����  �����  -���.  -���.  �����  �      B  , ,���  /���  ����Z  ����Z  /���  /      B  , ,����  /����  ����  ����  /����  /      B  , ,����   �����  c���  c���   �����   �      B  , ,���%   ����%  c����  c����   ����%   �      B  , ,���s   ����s  c���  c���   ����s   �      B  , ,����   �����  c���k  c���k   �����   �      B  , ,���   ����  c����  c����   ����   �      B  , ,���]   ����]  c���  c���   ����]   �      B  , ,���L  /���L  �����  �����  /���L  /      B  , ,����  /����  ����D  ����D  /����  /      B  , ,����  /����  �����  �����  /����  /      B  , ,���6  /���6  �����  �����  /���6  /      B  , ,����  /����  ����.  ����.  /����  /      B  , ,���  ����  ����Z  ����Z  ����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,���L  ����L  �����  �����  ����L  �      B  , ,����  �����  ����D  ����D  �����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,���6  ����6  �����  �����  ����6  �      B  , ,����  �����  ����.  ����.  �����  �      B  , ,���  +���  ����Z  ����Z  +���  +      B  , ,����  +����  ����  ����  +����  +      B  , ,���L  +���L  �����  �����  +���L  +      B  , ,������	����������L�������L���	������	      B  , ,��������������������������������������      B  , ,���*�������*�����������������������*����      B  , ,���x�������x�������"�������"�������x����      B  , ,�������������������p�������p������������      B  , ,�����������������������������������      B  , ,���b�������b���������������������b����      B  , ,�����������������Z�������Z�����������      B  , ,��������������������������������������      B  , ,���L�������L�����������������������L����      B  , ,�������������������D�������D������������      B  , ,����������������������������������������      B  , ,���6�������6�����������������������6����      B  , ,�������������������.�������.������������      B  , ,���������������}������}���������������      B  , ,���L�������L���}�������}�����������L����      B  , ,���������������}���D���}���D������������      B  , ,���������������}�������}����������������      B  , ,���6�������6���}�������}�����������6����      B  , ,���������������}���.���}���.������������      B  , ,������������)���Z���)���Z���������      B  , ,��������������)������)�������������      B  , ,���L������L���)�������)����������L���      B  , ,��������������)���D���)���D����������      B  , ,��������������)�������)��������������      B  , ,���6������6���)�������)����������6���      B  , ,��������������)���.���)���.����������      B  , ,������+����������Z�������Z���+������+      B  , ,�������+���������������������+�������+      B  , ,���L���+���L�������������������+���L���+      B  , ,�������+�����������D�������D���+�������+      B  , ,�������+�����������������������+�������+      B  , ,���6���+���6�������������������+���6���+      B  , ,�������+�����������.�������.���+�������+      B  , ,���������������G������G���������������      B  , ,���%�������%���G�������G�����������%����      B  , ,���s�������s���G������G����������s����      B  , ,���������������G���k���G���k������������      B  , ,�������������G�������G���������������      B  , ,���]�������]���G������G����������]����      B  , ,������'����������Z�������Z���'������'      B  , ,�������'���������������������'�������'      B  , ,���L���'���L�������������������'���L���'      B  , ,�������'�����������D�������D���'�������'      B  , ,�������'�����������������������'�������'      B  , ,���6���'���6�������������������'���6���'      B  , ,�������'�����������.�������.���'�������'      B  , ,�������������}���Z���}���Z�����������      B  , ,���b������b���)������)���������b���      B  , ,���b���'���b�����������������'���b���'      B  , ,�������������G������G��������������      B  , ,���Q�������Q���G�������G�����������Q����      B  , ,�������������G���I���G���I�����������      B  , ,���������������G������G���������������      B  , ,���;�������;���G�������G�����������;����      B  , ,�������������G���3���G���3�����������      B  , ,������]���������L������L���]������]      B  , ,�������+���������������������+�������+      B  , ,���*���+���*�������������������+���*���+      B  , ,���x���+���x�������"�������"���+���x���+      B  , ,�������+�����������p�������p���+�������+      B  , ,������+��������������������+������+      B  , ,���b���+���b�����������������+���b���+      B  , ,����������������L�������L���������      B  , ,����������������L�������L���������      B  , ,���������������}������}���������������      B  , ,���*�������*���}�������}�����������*����      B  , ,���x�������x���}���"���}���"�������x����      B  , ,���������������}���p���}���p������������      B  , ,�������������}������}��������������      B  , ,���b�������b���}������}����������b����      B  , ,�������������W���L���W���L�����������      B  , ,������Y���������L������L���Y������Y      B  , ,�������'���������������������'�������'      B  , ,���*���'���*�������������������'���*���'      B  , ,���x���'���x�������"�������"���'���x���'      B  , ,�������'�����������p�������p���'�������'      B  , ,������'��������������������'������'      B  , ,�������������[���L���[���L�����������      B  , ,��������������)������)�������������      B  , ,���*������*���)�������)����������*���      B  , ,���x������x���)���"���)���"������x���      B  , ,��������������)���p���)���p����������      B  , ,������������)������)������������      B  , ,�������������_���L���_���L�����������      B  , ,���������������-������-���������������      B  , ,���*�������*���-�������-�����������*����      B  , ,���x�������x���-���"���-���"�������x����      B  , ,���������������-���p���-���p������������      B  , ,�������������-������-��������������      B  , ,���b�������b���-������-����������b����      B  , ,������a���������L������L���a������a      B  , ,�������/���������������������/�������/      B  , ,���*���/���*�������������������/���*���/      B  , ,���x���/���x�������"�������"���/���x���/      B  , ,�������/�����������p�������p���/�������/      B  , ,������/��������������������/������/      B  , ,���b���/���b�����������������/���b���/      B  , ,���������������L������L���������      B  , ,������������������������������������      B  , ,���*�������*���������������������*����      B  , ,���x�������x������"������"�������x����      B  , ,������������������p������p������������      B  , ,���������������������������������      B  , ,���b�������b�������������������b����      B  , ,������������c���L���c���L���������      B  , ,������e���������L������L���e������e      B  , ,������g��������������������g������g      B  , ,���q���g���q���������������g���q���g      B  , ,�������g����������o������o���g�������g      B  , ,������g��������������������g������g      B  , ,���m���g���m���������������g���m���g      B  , ,�������g����������k������k���g�������g      B  , ,������g������������������g������g      B  , ,���i���g���i���������������g���i���g      B  , ,������g���������g������g���g������g      B  , ,������g������������������g������g      B  , ,���6�������6���-�������-�����������6����      B  , ,���������������-���.���-���.������������      B  , ,����������������Z������Z�����������      B  , ,������������������������������������      B  , ,���L�������L���������������������L����      B  , ,������������������D������D������������      B  , ,��������������������������������������      B  , ,���6�������6���������������������6����      B  , ,������������������.������.������������      B  , ,������/����������Z�������Z���/������/      B  , ,�������/���������������������/�������/      B  , ,���L���/���L�������������������/���L���/      B  , ,�������/�����������D�������D���/�������/      B  , ,�������/�����������������������/�������/      B  , ,���6���/���6�������������������/���6���/      B  , ,�������/�����������.�������.���/�������/      B  , ,�������������-���Z���-���Z�����������      B  , ,���������������-������-���������������      B  , ,���L�������L���-�������-�����������L����      B  , ,���������������-���D���-���D������������      B  , ,���������������-�������-����������������      B  , ,���e���g���e���������������g���e���g      B  , ,������g���������c������c���g������g      B  , ,������g������������������g������g      B  , ,���a���g���a���������������g���a���g      B  , ,�������g����������_������_���g�������g      B  , ,���	���g���	�����������������g���	���g      B  , ,���]���g���]���������������g���]���g      B  , ,�������g����������[������[���g�������g      B  , ,������g��������������������g������g      B  , ,���Y���g���Y���������������g���Y���g      B  , ,�������g����������W������W���g�������g      B  , ,������g��������������������g������g      B  , ,   �����   �����  |����  |����   �����      B  , ,   ����   ����  �����  �����   ����      B  , ,  n����  n����  ����  ����  n����      B  , ,  �����  �����  f����  f����  �����      B  , ,  

����  

����  
�����  
�����  

����      B  , ,  X����  X����  ����  ����  X����      B  , ,  �����  �����  P����  P����  �����      B  , ,  �����  �����  �����  �����  �����      B  , ,  B����  B����  �����  �����  B����      B  , ,  �����  �����  :����  :����  �����      B  , ,  �����  �����  �����  �����  �����      B  , ,  ,����  ,����  �����  �����  ,����      B  , ,  z����  z����  $����  $����  z����      B  , ,  ����	  �����  ^����  ^���	  ����	      B  , ,  z����  z���}  $���}  $����  z����      B  , ,  ����  �����  ^����  ^���  ����      B  , ,  �����  ����}  ����}  �����  �����      B  , ,  ,����  ,���}  ����}  �����  ,����      B  , ,  ����'  �����  �����  ����'  ����'      B  , ,  B���'  B����  �����  ����'  B���'      B  , ,  ����'  �����  :����  :���'  ����'      B  , ,  ����'  �����  �����  ����'  ����'      B  , ,  ,���'  ,����  �����  ����'  ,���'      B  , ,  z���'  z����  $����  $���'  z���'      B  , ,  ����Y  ����  ^���  ^���Y  ����Y      B  , ,  ����  ����)  ����)  ����  ����      B  , ,  B���  B���)  ����)  ����  B���      B  , ,  ����  ����)  :���)  :���  ����      B  , ,  ����  ����)  ����)  ����  ����      B  , ,  ,���  ,���)  ����)  ����  ,���      B  , ,  z���  z���)  $���)  $���  z���      B  , ,  �����  ����[  ^���[  ^����  �����      B  , ,  �����  ����G  w���G  w����  �����      B  , ,  ����  ���G  ����G  �����  ����      B  , ,  i����  i���G  ���G  ����  i����      B  , ,  �����  ����G  a���G  a����  �����      B  , ,  ����  ���G  ����G  �����  ����      B  , ,  S����  S���G  ����G  �����  S����      B  , ,  ����  �����  ^����  ^���  ����      B  , ,  �����  ����W  ^���W  ^����  �����      B  , ,  ����+  �����  �����  ����+  ����+      B  , ,  B���+  B����  �����  ����+  B���+      B  , ,  ����+  �����  :����  :���+  ����+      B  , ,  ����+  �����  �����  ����+  ����+      B  , ,  ,���+  ,����  �����  ����+  ,���+      B  , ,  z���+  z����  $����  $���+  z���+      B  , ,  ����]  ����  ^���  ^���]  ����]      B  , ,  �����  ����}  ����}  �����  �����      B  , ,  B����  B���}  ����}  �����  B����      B  , ,  �����  ����}  :���}  :����  �����      B  , ,  ����  ���G  )���G  )����  ����      B  , ,   ����   ����)  |���)  |���   ����      B  , ,   ���   ���)  ����)  ����   ���      B  , ,  n���  n���)  ���)  ���  n���      B  , ,  ����  ����)  f���)  f���  ����      B  , ,  

���  

���)  
����)  
����  

���      B  , ,  X���  X���)  ���)  ���  X���      B  , ,  ����  ����)  P���)  P���  ����      B  , ,  �����  ����G  ����G  �����  �����      B  , ,   ����'   �����  |����  |���'   ����'      B  , ,   ����+   �����  |����  |���+   ����+      B  , ,   ���+   ����  �����  ����+   ���+      B  , ,  n���+  n����  ����  ���+  n���+      B  , ,  ����+  �����  f����  f���+  ����+      B  , ,  

���+  

����  
�����  
����+  

���+      B  , ,  X���+  X����  ����  ���+  X���+      B  , ,  ����+  �����  P����  P���+  ����+      B  , ,   ���'   ����  �����  ����'   ���'      B  , ,  n���'  n����  ����  ���'  n���'      B  , ,  ����'  �����  f����  f���'  ����'      B  , ,  

���'  

����  
�����  
����'  

���'      B  , ,  X���'  X����  ����  ���'  X���'      B  , ,  ����'  �����  P����  P���'  ����'      B  , ,  G����  G���G  ����G  �����  G����      B  , ,   �����   ����}  |���}  |����   �����      B  , ,   ����   ���}  ����}  �����   ����      B  , ,  n����  n���}  ���}  ����  n����      B  , ,  �����  ����}  f���}  f����  �����      B  , ,  

����  

���}  
����}  
�����  

����      B  , ,  X����  X���}  ���}  ����  X����      B  , ,  �����  ����}  P���}  P����  �����      B  , ,  �����  ����G  ?���G  ?����  �����      B  , ,  �����  ����G  	����G  	�����  �����      B  , ,  1����  1���G  ����G  �����  1����      B  , ,  �����  ����-  f���-  f����  �����      B  , ,  

����  

���-  
����-  
�����  

����      B  , ,  X����  X���-  ���-  ����  X����      B  , ,  �����  ����-  P���-  P����  �����      B  , ,   ����/   �����  |����  |���/   ����/      B  , ,   ���/   ����  �����  ����/   ���/      B  , ,  n���/  n����  ����  ���/  n���/      B  , ,  ����/  �����  f����  f���/  ����/      B  , ,  

���/  

����  
�����  
����/  

���/      B  , ,  X���/  X����  ����  ���/  X���/      B  , ,  ����/  �����  P����  P���/  ����/      B  , ,   �����   ����  |���  |����   �����      B  , ,   ����   ���  ����  �����   ����      B  , ,  n����  n���  ���  ����  n����      B  , ,  �����  ����  f���  f����  �����      B  , ,  

����  

���  
����  
�����  

����      B  , ,  X����  X���  ���  ����  X����      B  , ,  �����  ����  P���  P����  �����      B  , ,   �����   ����-  |���-  |����   �����      B  , ,   ����   ���-  ����-  �����   ����      B  , ,  n����  n���-  ���-  ����  n����      B  , ,   U���g   U���   ����   ����g   U���g      B  , ,  ����g  ����  S���  S���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  Q���g  Q���  ����  ����g  Q���g      B  , ,  ����g  ����  O���  O���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  M���g  M���  ����  ����g  M���g      B  , ,  	����g  	����  
K���  
K���g  	����g      B  , ,  
����g  
����  ����  ����g  
����g      B  , ,  I���g  I���  ����  ����g  I���g      B  , ,  ����g  ����  G���  G���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  �����  ����_  ^���_  ^����  �����      B  , ,  �����  ����  ����  �����  �����      B  , ,  B����  B���  ����  �����  B����      B  , ,  �����  ����  :���  :����  �����      B  , ,  �����  ����  ����  �����  �����      B  , ,  ,����  ,���  ����  �����  ,����      B  , ,  z����  z���  $���  $����  z����      B  , ,  ����  ����  ^���  ^���  ����      B  , ,  ����/  �����  �����  ����/  ����/      B  , ,  ����  ����c  ^���c  ^���  ����      B  , ,  B���/  B����  �����  ����/  B���/      B  , ,  ����e  ����  ^���  ^���e  ����e      B  , ,  ����/  �����  :����  :���/  ����/      B  , ,  ����/  �����  �����  ����/  ����/      B  , ,  ,���/  ,����  �����  ����/  ,���/      B  , ,  z���/  z����  $����  $���/  z���/      B  , ,  ����a  ����  ^���  ^���a  ����a      B  , ,  �����  ����-  ����-  �����  �����      B  , ,  B����  B���-  ����-  �����  B����      B  , ,  �����  ����-  :���-  :����  �����      B  , ,  �����  ����-  ����-  �����  �����      B  , ,  ,����  ,���-  ����-  �����  ,����      B  , ,  z����  z���-  $���-  $����  z����      B  , ,  E���g  E���  ����  ����g  E���g      B  , ,  ����g  ����  C���  C���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  A���g  A���  ����  ����g  A���g      B  , ,  ����g  ����  ?���  ?���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  =���g  =���  ����  ����g  =���g      B  , ,  ����g  ����  ;���  ;���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  9���g  9���  ����  ����g  9���g      _   ,������9���  �  a  �  a���9������9      C   ,���  ����  �  ^  �  ^  ����  �      C   ,���������  ����L  ����L���������      C   ,���[   ����[  c   �  c   �   ����[   �      C   ,���[�������[���G   ����G   ��������[����      C   ,  ����  �  �  ^  �  ^���  ����      C   ,������g������  ^���  ^���g������g      C   ,  

  :  

    
�    
�  :  

  :      C   ,  X  :  X          :  X  :      C   ,  �  :  �    P    P  :  �  :      C   ,  �  :  �    �    �  :  �  :      C   ,  B  :  B    �    �  :  B  :      C   ,  �  :  �    :    :  :  �  :      C   ,  �  :  �    �    �  :  �  :      C   ,  ,  :  ,    �    �  :  ,  :      C   ,  z  :  z    $    $  :  z  :      C   ,   �  :   �    |    |  :   �  :      C   ,  �   �  �  c  �  c  �   �  �   �      C   ,  �   �  �  c  A  c  A   �  �   �      C   ,  E   �  E  c  �  c  �   �  E   �      C   ,  �   �  �  c  	�  c  	�   �  �   �      C   ,  
�   �  
�  c  +  c  +   �  
�   �      C   ,  /   �  /  c  y  c  y   �  /   �      C   ,  }   �  }  c  �  c  �   �  }   �      C   ,  �   �  �  c    c     �  �   �      C   ,     �    c  c  c  c   �     �      C   ,  g   �  g  c  �  c  �   �  g   �      C   ,  �   �  �  c  �  c  �   �  �   �      C   ,     �    c  M  c  M   �     �      C   ,     :       �    �  :     :      C   ,  n  :  n          :  n  :      C   ,  �  :  �    f    f  :  �  :      C   ,���   ����  c����  c����   ����   �      C   ,����   �����  c���5  c���5   �����   �      C   ,���9   ����9  c����  c����   ����9   �      C   ,���   ����  c����  c����   ����   �      C   ,����   �����  c���  c���   �����   �      C   ,���#   ����#  c���m  c���m   ����#   �      C   ,���q   ����q  c����  c����   ����q   �      C   ,����   �����  c���	  c���	   �����   �      C   ,���   ����  c���W  c���W   ����   �      C   ,����  :����  ���  ���  :����  :      C   ,���*  :���*  ����  ����  :���*  :      C   ,���x  :���x  ���"  ���"  :���x  :      C   ,����  :����  ���p  ���p  :����  :      C   ,���  :���  ���  ���  :���  :      C   ,���b  :���b  ���  ���  :���b  :      C   ,���  :���  ���Z  ���Z  :���  :      C   ,����  :����  ���  ���  :����  :      C   ,���L  :���L  ����  ����  :���L  :      C   ,����  :����  ���D  ���D  :����  :      C   ,����  :����  ����  ����  :����  :      C   ,���6  :���6  ����  ����  :���6  :      C   ,����  :����  ���.  ���.  :����  :      C   ,���   ����  c����  c����   ����   �      C   ,���   ����  c���K  c���K   ����   �      C   ,���O   ����O  c���  c���   ����O   �      C   ,�������������G�������G���������������      C   ,���������������G���5���G���5������������      C   ,���9�������9���G�������G�����������9����      C   ,�������������G�������G���������������      C   ,���������������G������G���������������      C   ,���#�������#���G���m���G���m�������#����      C   ,���q�������q���G�������G�����������q����      C   ,���������������G���	���G���	������������      C   ,�������������G���W���G���W�����������      C   ,�������������G�������G���������������      C   ,��������������������������������������      C   ,���*�������*�����������������������*����      C   ,���x�������x�������"�������"�������x����      C   ,�������������������p�������p������������      C   ,�����������������������������������      C   ,���b�������b���������������������b����      C   ,�����������������Z�������Z�����������      C   ,��������������������������������������      C   ,���L�������L�����������������������L����      C   ,�������������������D�������D������������      C   ,����������������������������������������      C   ,���6�������6�����������������������6����      C   ,�������������������.�������.������������      C   ,�������������G���K���G���K�����������      C   ,���O�������O���G������G����������O����      C   ,  �����  ����G  	����G  	�����  �����      C   ,  
�����  
����G  +���G  +����  
�����      C   ,  /����  /���G  y���G  y����  /����      C   ,  }����  }���G  ����G  �����  }����      C   ,  �����  ����G  ���G  ����  �����      C   ,  ����  ���G  c���G  c����  ����      C   ,  g����  g���G  ����G  �����  g����      C   ,  �����  ����G  ����G  �����  �����      C   ,  ����  ���G  M���G  M����  ����      C   ,  �����  ����G  ����G  �����  �����      C   ,   �����   �����  |����  |����   �����      C   ,   ����   ����  �����  �����   ����      C   ,  n����  n����  ����  ����  n����      C   ,  �����  �����  f����  f����  �����      C   ,  

����  

����  
�����  
�����  

����      C   ,  X����  X����  ����  ����  X����      C   ,  �����  �����  P����  P����  �����      C   ,  �����  �����  �����  �����  �����      C   ,  B����  B����  �����  �����  B����      C   ,  �����  �����  :����  :����  �����      C   ,  �����  �����  �����  �����  �����      C   ,  ,����  ,����  �����  �����  ,����      C   ,  z����  z����  $����  $����  z����      C   ,  �����  ����G  A���G  A����  �����      C   ,  E����  E���G  ����G  �����  E����      C  , ,����   �����  c   U  c   U   �����   �      C  , ,���������������G   U���G   U������������      C  , ,  �  �  �  k  P  k  P  �  �  �      C  , ,  �  �  �  k  �  k  �  �  �  �      C  , ,  B  �  B  k  �  k  �  �  B  �      C  , ,  �  �  �  k  :  k  :  �  �  �      C  , ,  �  �  �  k  �  k  �  �  �  �      C  , ,  ,  �  ,  k  �  k  �  �  ,  �      C  , ,  z  �  z  k  $  k  $  �  z  �      C  , ,  �  Y  �    P    P  Y  �  Y      C  , ,  �  Y  �    �    �  Y  �  Y      C  , ,  B  Y  B    �    �  Y  B  Y      C  , ,  �  Y  �    :    :  Y  �  Y      C  , ,  �  Y  �    �    �  Y  �  Y      C  , ,  ,  Y  ,    �    �  Y  ,  Y      C  , ,  z  Y  z    $    $  Y  z  Y      C  , ,  �  	�  �  
�  P  
�  P  	�  �  	�      C  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      C  , ,  B  	�  B  
�  �  
�  �  	�  B  	�      C  , ,  �  	�  �  
�  :  
�  :  	�  �  	�      C  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      C  , ,  ,  	�  ,  
�  �  
�  �  	�  ,  	�      C  , ,  z  	�  z  
�  $  
�  $  	�  z  	�      C  , ,  �  �  �  	3  P  	3  P  �  �  �      C  , ,  �  �  �  	3  �  	3  �  �  �  �      C  , ,  B  �  B  	3  �  	3  �  �  B  �      C  , ,  �  �  �  	3  :  	3  :  �  �  �      C  , ,  �  �  �  	3  �  	3  �  �  �  �      C  , ,  ,  �  ,  	3  �  	3  �  �  ,  �      C  , ,  z  �  z  	3  $  	3  $  �  z  �      C  , ,  �  !  �  �  P  �  P  !  �  !      C  , ,  �  !  �  �  �  �  �  !  �  !      C  , ,  B  !  B  �  �  �  �  !  B  !      C  , ,  �  !  �  �  :  �  :  !  �  !      C  , ,  �  !  �  �  �  �  �  !  �  !      C  , ,  ,  !  ,  �  �  �  �  !  ,  !      C  , ,  z  !  z  �  $  �  $  !  z  !      C  , ,  �  �  �  k  f  k  f  �  �  �      C  , ,  

  �  

  k  
�  k  
�  �  

  �      C  , ,   �  �   �  	3  |  	3  |  �   �  �      C  , ,     �     	3  �  	3  �  �     �      C  , ,  n  �  n  	3    	3    �  n  �      C  , ,  �  �  �  	3  f  	3  f  �  �  �      C  , ,  

  �  

  	3  
�  	3  
�  �  

  �      C  , ,  X  �  X  	3    	3    �  X  �      C  , ,   �  Y   �    |    |  Y   �  Y      C  , ,     Y       �    �  Y     Y      C  , ,  n  Y  n          Y  n  Y      C  , ,   �  	�   �  
�  |  
�  |  	�   �  	�      C  , ,     	�     
�  �  
�  �  	�     	�      C  , ,  n  	�  n  
�    
�    	�  n  	�      C  , ,  �  	�  �  
�  f  
�  f  	�  �  	�      C  , ,   �  !   �  �  |  �  |  !   �  !      C  , ,     !     �  �  �  �  !     !      C  , ,  n  !  n  �    �    !  n  !      C  , ,  �  !  �  �  f  �  f  !  �  !      C  , ,  

  !  

  �  
�  �  
�  !  

  !      C  , ,  X  !  X  �    �    !  X  !      C  , ,  

  	�  

  
�  
�  
�  
�  	�  

  	�      C  , ,  X  	�  X  
�    
�    	�  X  	�      C  , ,  �  Y  �    f    f  Y  �  Y      C  , ,  

  Y  

    
�    
�  Y  

  Y      C  , ,  X  Y  X          Y  X  Y      C  , ,  X  �  X  k    k    �  X  �      C  , ,  n  �  n  k    k    �  n  �      C  , ,   �  �   �  k  |  k  |  �   �  �      C  , ,     �     k  �  k  �  �     �      C  , ,  n  �  n  c    c    �  n  �      C  , ,  �  �  �  c  f  c  f  �  �  �      C  , ,  

  �  

  c  
�  c  
�  �  

  �      C  , ,  X  �  X  c    c    �  X  �      C  , ,   �  Q   �  �  |  �  |  Q   �  Q      C  , ,     Q     �  �  �  �  Q     Q      C  , ,  n  Q  n  �    �    Q  n  Q      C  , ,  �  Q  �  �  f  �  f  Q  �  Q      C  , ,  

  Q  

  �  
�  �  
�  Q  

  Q      C  , ,  X  Q  X  �    �    Q  X  Q      C  , ,   �  �   �  �  |  �  |  �   �  �      C  , ,     �     �  �  �  �  �     �      C  , ,  n  �  n  �    �    �  n  �      C  , ,  �  �  �  �  f  �  f  �  �  �      C  , ,  

  �  

  �  
�  �  
�  �  

  �      C  , ,  X  �  X  �    �    �  X  �      C  , ,   �  �   �  c  |  c  |  �   �  �      C  , ,  �   �  �  c  �  c  �   �  �   �      C  , ,  G   �  G  c  �  c  �   �  G   �      C  , ,  �   �  �  c  ?  c  ?   �  �   �      C  , ,  �   �  �  c  	�  c  	�   �  �   �      C  , ,  1   �  1  c  �  c  �   �  1   �      C  , ,     �    c  )  c  )   �     �      C  , ,     �     c  �  c  �  �     �      C  , ,  z  �  z  c  $  c  $  �  z  �      C  , ,  �  �  �  c  P  c  P  �  �  �      C  , ,  �  �  �  c  �  c  �  �  �  �      C  , ,  B  �  B  c  �  c  �  �  B  �      C  , ,  �  �  �  c  :  c  :  �  �  �      C  , ,  �  �  �  c  �  c  �  �  �  �      C  , ,  �  �  �  �  P  �  P  �  �  �      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,  B  �  B  �  �  �  �  �  B  �      C  , ,  �  �  �  �  :  �  :  �  �  �      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,  ,  �  ,  �  �  �  �  �  ,  �      C  , ,  z  �  z  �  $  �  $  �  z  �      C  , ,  ,  �  ,  c  �  c  �  �  ,  �      C  , ,  �  Q  �  �  P  �  P  Q  �  Q      C  , ,  �  Q  �  �  �  �  �  Q  �  Q      C  , ,  B  Q  B  �  �  �  �  Q  B  Q      C  , ,  �  Q  �  �  :  �  :  Q  �  Q      C  , ,  �  Q  �  �  �  �  �  Q  �  Q      C  , ,  ,  Q  ,  �  �  �  �  Q  ,  Q      C  , ,  �   �  �  c  w  c  w   �  �   �      C  , ,     �    c  �  c  �   �     �      C  , ,  i   �  i  c    c     �  i   �      C  , ,  �   �  �  c  a  c  a   �  �   �      C  , ,     �    c  �  c  �   �     �      C  , ,  S   �  S  c  �  c  �   �  S   �      C  , ,  z  Q  z  �  $  �  $  Q  z  Q      C  , ,����  	�����  
����  
����  	�����  	�      C  , ,���L  	����L  
�����  
�����  	����L  	�      C  , ,����  	�����  
����D  
����D  	�����  	�      C  , ,����  	�����  
�����  
�����  	�����  	�      C  , ,���6  	����6  
�����  
�����  	����6  	�      C  , ,����  	�����  
����.  
����.  	�����  	�      C  , ,����  Y����  ���  ���  Y����  Y      C  , ,���L  Y���L  ����  ����  Y���L  Y      C  , ,����  Y����  ���D  ���D  Y����  Y      C  , ,����  Y����  ����  ����  Y����  Y      C  , ,���6  Y���6  ����  ����  Y���6  Y      C  , ,����  Y����  ���.  ���.  Y����  Y      C  , ,����  �����  	3���  	3���  �����  �      C  , ,���L  ����L  	3����  	3����  ����L  �      C  , ,����  �����  	3���D  	3���D  �����  �      C  , ,����  �����  	3����  	3����  �����  �      C  , ,���6  ����6  	3����  	3����  ����6  �      C  , ,����  �����  	3���.  	3���.  �����  �      C  , ,����  �����  k���  k���  �����  �      C  , ,���L  ����L  k����  k����  ����L  �      C  , ,����  �����  k���D  k���D  �����  �      C  , ,����  �����  k����  k����  �����  �      C  , ,���6  ����6  k����  k����  ����6  �      C  , ,����  �����  k���.  k���.  �����  �      C  , ,����  !����  ����  ����  !����  !      C  , ,���L  !���L  �����  �����  !���L  !      C  , ,����  !����  ����D  ����D  !����  !      C  , ,����  !����  �����  �����  !����  !      C  , ,���6  !���6  �����  �����  !���6  !      C  , ,����  !����  ����.  ����.  !����  !      C  , ,���b  ����b  	3���  	3���  ����b  �      C  , ,���  ����  	3���Z  	3���Z  ����  �      C  , ,����  Y����  ���  ���  Y����  Y      C  , ,���*  Y���*  ����  ����  Y���*  Y      C  , ,���x  Y���x  ���"  ���"  Y���x  Y      C  , ,����  Y����  ���p  ���p  Y����  Y      C  , ,���  Y���  ���  ���  Y���  Y      C  , ,���b  Y���b  ���  ���  Y���b  Y      C  , ,����  �����  k���  k���  �����  �      C  , ,���*  ����*  k����  k����  ����*  �      C  , ,���x  ����x  k���"  k���"  ����x  �      C  , ,����  �����  k���p  k���p  �����  �      C  , ,���  ����  k���  k���  ����  �      C  , ,���b  ����b  k���  k���  ����b  �      C  , ,���  ����  k���Z  k���Z  ����  �      C  , ,���  Y���  ���Z  ���Z  Y���  Y      C  , ,���*  	����*  
�����  
�����  	����*  	�      C  , ,���x  	����x  
����"  
����"  	����x  	�      C  , ,����  	�����  
����p  
����p  	�����  	�      C  , ,���  	����  
����  
����  	����  	�      C  , ,���b  	����b  
����  
����  	����b  	�      C  , ,����  !����  ����  ����  !����  !      C  , ,���*  !���*  �����  �����  !���*  !      C  , ,���x  !���x  ����"  ����"  !���x  !      C  , ,����  !����  ����p  ����p  !����  !      C  , ,���  !���  ����  ����  !���  !      C  , ,���b  !���b  ����  ����  !���b  !      C  , ,���  !���  ����Z  ����Z  !���  !      C  , ,���  	����  
����Z  
����Z  	����  	�      C  , ,����  �����  	3���  	3���  �����  �      C  , ,���*  ����*  	3����  	3����  ����*  �      C  , ,���x  ����x  	3���"  	3���"  ����x  �      C  , ,����  �����  	3���p  	3���p  �����  �      C  , ,���  ����  	3���  	3���  ����  �      C  , ,����  	�����  
����  
����  	�����  	�      C  , ,���  ����  c���  c���  ����  �      C  , ,���b  ����b  c���  c���  ����b  �      C  , ,����  Q����  ����  ����  Q����  Q      C  , ,���*  Q���*  �����  �����  Q���*  Q      C  , ,���x  Q���x  ����"  ����"  Q���x  Q      C  , ,����  Q����  ����p  ����p  Q����  Q      C  , ,���  Q���  ����  ����  Q���  Q      C  , ,���   ����  c���  c���   ����   �      C  , ,���Q   ����Q  c����  c����   ����Q   �      C  , ,���   ����  c���I  c���I   ����   �      C  , ,����   �����  c���  c���   �����   �      C  , ,���;   ����;  c����  c����   ����;   �      C  , ,���   ����  c���3  c���3   ����   �      C  , ,���b  Q���b  ����  ����  Q���b  Q      C  , ,����  �����  ����  ����  �����  �      C  , ,���*  ����*  �����  �����  ����*  �      C  , ,���x  ����x  ����"  ����"  ����x  �      C  , ,����  �����  ����p  ����p  �����  �      C  , ,���  ����  ����  ����  ����  �      C  , ,���b  ����b  ����  ����  ����b  �      C  , ,���  ����  ����Z  ����Z  ����  �      C  , ,���  Q���  ����Z  ����Z  Q���  Q      C  , ,���  ����  c���Z  c���Z  ����  �      C  , ,����  �����  c���  c���  �����  �      C  , ,���*  ����*  c����  c����  ����*  �      C  , ,���x  ����x  c���"  c���"  ����x  �      C  , ,����  �����  c���p  c���p  �����  �      C  , ,����  �����  �����  �����  �����  �      C  , ,���6  ����6  �����  �����  ����6  �      C  , ,����  �����  ����.  ����.  �����  �      C  , ,����  Q����  ����D  ����D  Q����  Q      C  , ,����   �����  c���  c���   �����   �      C  , ,���%   ����%  c����  c����   ����%   �      C  , ,���s   ����s  c���  c���   ����s   �      C  , ,����   �����  c���k  c���k   �����   �      C  , ,���   ����  c����  c����   ����   �      C  , ,���]   ����]  c���  c���   ����]   �      C  , ,����  Q����  �����  �����  Q����  Q      C  , ,���6  Q���6  �����  �����  Q���6  Q      C  , ,����  Q����  ����.  ����.  Q����  Q      C  , ,����  �����  c���D  c���D  �����  �      C  , ,����  �����  c����  c����  �����  �      C  , ,���6  ����6  c����  c����  ����6  �      C  , ,����  �����  c���.  c���.  �����  �      C  , ,����  �����  c���  c���  �����  �      C  , ,���L  ����L  c����  c����  ����L  �      C  , ,����  Q����  ����  ����  Q����  Q      C  , ,���L  Q���L  �����  �����  Q���L  Q      C  , ,����  �����  ����  ����  �����  �      C  , ,���L  ����L  �����  �����  ����L  �      C  , ,����  �����  ����D  ����D  �����  �      C  , ,���������������G������G���������������      C  , ,���%�������%���G�������G�����������%����      C  , ,���s�������s���G������G����������s����      C  , ,���������������G���k���G���k������������      C  , ,�������������G�������G���������������      C  , ,���]�������]���G������G����������]����      C  , ,�������m�������������������m�������m      C  , ,���L���m���L�����������������m���L���m      C  , ,�������m����������D������D���m�������m      C  , ,�������m���������������������m�������m      C  , ,���6���m���6�����������������m���6���m      C  , ,�������m����������.������.���m�������m      C  , ,�����������������������������������      C  , ,���L������L����������������������L���      C  , ,������������������D�������D����������      C  , ,�������������������������������������      C  , ,���6������6����������������������6���      C  , ,������������������.�������.����������      C  , ,���������������G������G���������������      C  , ,���L�������L���G�������G�����������L����      C  , ,���������������G���D���G���D������������      C  , ,���������������G�������G����������������      C  , ,���6�������6���G�������G�����������6����      C  , ,���������������G���.���G���.������������      C  , ,�������������G������G��������������      C  , ,�����������������������������������      C  , ,���*������*����������������������*���      C  , ,���x������x�������"�������"������x���      C  , ,������������������p�������p����������      C  , ,��������������������������������      C  , ,���b������b��������������������b���      C  , ,����������������Z�������Z���������      C  , ,�������m�������������������m�������m      C  , ,���*���m���*�����������������m���*���m      C  , ,���x���m���x������"������"���m���x���m      C  , ,�������m����������p������p���m�������m      C  , ,������m������������������m������m      C  , ,���b���m���b���������������m���b���m      C  , ,���������������G������G���������������      C  , ,���*�������*���G�������G�����������*����      C  , ,���x�������x���G���"���G���"�������x����      C  , ,���������������G���p���G���p������������      C  , ,�������������G������G��������������      C  , ,���b�������b���G������G����������b����      C  , ,�������������G���Z���G���Z�����������      C  , ,������m���������Z������Z���m������m      C  , ,�������������G���I���G���I�����������      C  , ,���������������G������G���������������      C  , ,���;�������;���G�������G�����������;����      C  , ,�������������G���3���G���3�����������      C  , ,���Q�������Q���G�������G�����������Q����      C  , ,�������5���������������������5�������5      C  , ,���*���5���*�������������������5���*���5      C  , ,���x���5���x�������"�������"���5���x���5      C  , ,�������5�����������p�������p���5�������5      C  , ,������5��������������������5������5      C  , ,���b���5���b�����������������5���b���5      C  , ,������5����������Z�������Z���5������5      C  , ,���������������w������w���������������      C  , ,���*�������*���w�������w�����������*����      C  , ,���x�������x���w���"���w���"�������x����      C  , ,���������������w���p���w���p������������      C  , ,�������������w������w��������������      C  , ,���b�������b���w������w����������b����      C  , ,�������������w���Z���w���Z�����������      C  , ,�������e�������������������e�������e      C  , ,���*���e���*�����������������e���*���e      C  , ,���x���e���x������"������"���e���x���e      C  , ,�������e����������p������p���e�������e      C  , ,������e������������������e������e      C  , ,���b���e���b���������������e���b���e      C  , ,������e���������Z������Z���e������e      C  , ,��������������������������������������      C  , ,���*�������*�����������������������*����      C  , ,���x�������x�������"�������"�������x����      C  , ,�������������������p�������p������������      C  , ,�����������������������������������      C  , ,���b�������b���������������������b����      C  , ,�����������������Z�������Z�����������      C  , ,��������������?������?�������������      C  , ,���*������*���?�������?����������*���      C  , ,���x������x���?���"���?���"������x���      C  , ,��������������?���p���?���p����������      C  , ,������������?������?������������      C  , ,���b������b���?������?���������b���      C  , ,������������?���Z���?���Z���������      C  , ,�������e����������D������D���e�������e      C  , ,�������e���������������������e�������e      C  , ,���6���e���6�����������������e���6���e      C  , ,�������e����������.������.���e�������e      C  , ,���L�������L���w�������w�����������L����      C  , ,���������������w���D���w���D������������      C  , ,���������������w�������w����������������      C  , ,���6�������6���w�������w�����������6����      C  , ,���������������w���.���w���.������������      C  , ,���L���5���L�������������������5���L���5      C  , ,�������5�����������D�������D���5�������5      C  , ,��������������������������������������      C  , ,���L�������L�����������������������L����      C  , ,�������������������D�������D������������      C  , ,����������������������������������������      C  , ,���6�������6�����������������������6����      C  , ,�������������������.�������.������������      C  , ,�������5�����������������������5�������5      C  , ,���6���5���6�������������������5���6���5      C  , ,�������5�����������.�������.���5�������5      C  , ,�������5���������������������5�������5      C  , ,���������������w������w���������������      C  , ,�������e�������������������e�������e      C  , ,���L���e���L�����������������e���L���e      C  , ,��������������?������?�������������      C  , ,���L������L���?�������?����������L���      C  , ,��������������?���D���?���D����������      C  , ,��������������?�������?��������������      C  , ,���6������6���?�������?����������6���      C  , ,��������������?���.���?���.����������      C  , ,  ����  �����  P����  P���  ����      C  , ,  ����  �����  �����  ����  ����      C  , ,  B���  B����  �����  ����  B���      C  , ,  ����  �����  :����  :���  ����      C  , ,  ����  �����  �����  ����  ����      C  , ,  ,���  ,����  �����  ����  ,���      C  , ,  z���  z����  $����  $���  z���      C  , ,  ����m  ����  P���  P���m  ����m      C  , ,  ����m  ����  ����  ����m  ����m      C  , ,  B���m  B���  ����  ����m  B���m      C  , ,  ����m  ����  :���  :���m  ����m      C  , ,  ����m  ����  ����  ����m  ����m      C  , ,  ,���m  ,���  ����  ����m  ,���m      C  , ,  z���m  z���  $���  $���m  z���m      C  , ,  �����  ����G  P���G  P����  �����      C  , ,  �����  ����G  ����G  �����  �����      C  , ,  B����  B���G  ����G  �����  B����      C  , ,  �����  ����G  :���G  :����  �����      C  , ,  �����  ����G  ����G  �����  �����      C  , ,  ,����  ,���G  ����G  �����  ,����      C  , ,  z����  z���G  $���G  $����  z����      C  , ,  �����  ����G  w���G  w����  �����      C  , ,  ����  ���G  ����G  �����  ����      C  , ,  i����  i���G  ���G  ����  i����      C  , ,  �����  ����G  a���G  a����  �����      C  , ,  ����  ���G  ����G  �����  ����      C  , ,  S����  S���G  ����G  �����  S����      C  , ,  n����  n���G  ���G  ����  n����      C  , ,  �����  ����G  f���G  f����  �����      C  , ,  

����  

���G  
����G  
�����  

����      C  , ,  X����  X���G  ���G  ����  X����      C  , ,  ����m  ����  f���  f���m  ����m      C  , ,  

���m  

���  
����  
����m  

���m      C  , ,  X���m  X���  ���  ���m  X���m      C  , ,  ����  �����  f����  f���  ����      C  , ,  

���  

����  
�����  
����  

���      C  , ,  X���  X����  ����  ���  X���      C  , ,   ���   ����  �����  ����   ���      C  , ,  �����  ����G  ?���G  ?����  �����      C  , ,  �����  ����G  	����G  	�����  �����      C  , ,  1����  1���G  ����G  �����  1����      C  , ,  ����  ���G  )���G  )����  ����      C  , ,  n���  n����  ����  ���  n���      C  , ,   ���m   ���  ����  ����m   ���m      C  , ,  n���m  n���  ���  ���m  n���m      C  , ,  G����  G���G  ����G  �����  G����      C  , ,   �����   ����G  |���G  |����   �����      C  , ,   ����   ���G  ����G  �����   ����      C  , ,  �����  ����G  ����G  �����  �����      C  , ,   ����m   ����  |���  |���m   ����m      C  , ,   ����   �����  |����  |���   ����      C  , ,  X����  X���w  ���w  ����  X����      C  , ,  

���5  

����  
�����  
����5  

���5      C  , ,  X���5  X����  ����  ���5  X���5      C  , ,   ����e   ����  |���  |���e   ����e      C  , ,   ���e   ���  ����  ����e   ���e      C  , ,   �����   �����  |����  |����   �����      C  , ,   ����   ����  �����  �����   ����      C  , ,  n����  n����  ����  ����  n����      C  , ,  �����  �����  f����  f����  �����      C  , ,  

����  

����  
�����  
�����  

����      C  , ,  X����  X����  ����  ����  X����      C  , ,  n���e  n���  ���  ���e  n���e      C  , ,  ����e  ����  f���  f���e  ����e      C  , ,  

���e  

���  
����  
����e  

���e      C  , ,  X���e  X���  ���  ���e  X���e      C  , ,   ���5   ����  �����  ����5   ���5      C  , ,  n���5  n����  ����  ���5  n���5      C  , ,  ����5  �����  f����  f���5  ����5      C  , ,   �����   ����w  |���w  |����   �����      C  , ,   ����   ���w  ����w  �����   ����      C  , ,  n����  n���w  ���w  ����  n����      C  , ,  �����  ����w  f���w  f����  �����      C  , ,  

����  

���w  
����w  
�����  

����      C  , ,   ����5   �����  |����  |���5   ����5      C  , ,   ����   ����?  |���?  |���   ����      C  , ,   ���   ���?  ����?  ����   ���      C  , ,  n���  n���?  ���?  ���  n���      C  , ,  ����  ����?  f���?  f���  ����      C  , ,  

���  

���?  
����?  
����  

���      C  , ,  X���  X���?  ���?  ���  X���      C  , ,  ����e  ����  :���  :���e  ����e      C  , ,  ����e  ����  ����  ����e  ����e      C  , ,  �����  �����  P����  P����  �����      C  , ,  �����  �����  �����  �����  �����      C  , ,  B����  B����  �����  �����  B����      C  , ,  �����  �����  :����  :����  �����      C  , ,  �����  �����  �����  �����  �����      C  , ,  ,����  ,����  �����  �����  ,����      C  , ,  z����  z����  $����  $����  z����      C  , ,  ,���e  ,���  ����  ����e  ,���e      C  , ,  z���e  z���  $���  $���e  z���e      C  , ,  ����5  �����  :����  :���5  ����5      C  , ,  ����5  �����  �����  ����5  ����5      C  , ,  �����  ����w  P���w  P����  �����      C  , ,  �����  ����w  ����w  �����  �����      C  , ,  B����  B���w  ����w  �����  B����      C  , ,  �����  ����w  :���w  :����  �����      C  , ,  �����  ����w  ����w  �����  �����      C  , ,  ,����  ,���w  ����w  �����  ,����      C  , ,  z����  z���w  $���w  $����  z����      C  , ,  ,���5  ,����  �����  ����5  ,���5      C  , ,  z���5  z����  $����  $���5  z���5      C  , ,  ����5  �����  P����  P���5  ����5      C  , ,  ����5  �����  �����  ����5  ����5      C  , ,  B���5  B����  �����  ����5  B���5      C  , ,  ����e  ����  P���  P���e  ����e      C  , ,  ����e  ����  ����  ����e  ����e      C  , ,  B���e  B���  ����  ����e  B���e      C  , ,  ����  ����?  P���?  P���  ����      C  , ,  ����  ����?  ����?  ����  ����      C  , ,  B���  B���?  ����?  ����  B���      C  , ,  ����  ����?  :���?  :���  ����      C  , ,  ����  ����?  ����?  ����  ����      C  , ,  ,���  ,���?  ����?  ����  ,���      C  , ,  z���  z���?  $���?  $���  z���      D   ,���o   ����o  �   �  �   �   ����o   �      D   ,���o������o���e   ����e   �������o���      D   ,  P  N  P    6    6  N  P  N      D   ,  �  N  �    �    �  N  �  N      D   ,  	�  N  	�    
�    
�  N  	�  N      D   ,  :  N  :            N  :  N      D   ,  �  N  �    n    n  N  �  N      D   ,  �  N  �    �    �  N  �  N      D   ,  $  N  $    
    
  N  $  N      D   ,  r  N  r    X    X  N  r  N      D   ,  �  N  �    �    �  N  �  N      D   ,    N      �    �  N    N      D   ,  \  N  \    B    B  N  \  N      D   ,   �  N   �    �    �  N   �  N      D   ,  �   �  �  �  �  �  �   �  �   �      D   ,     �    �  -  �  -   �     �      D   ,  Y   �  Y  �  {  �  {   �  Y   �      D   ,  �   �  �  �  	�  �  	�   �  �   �      D   ,  
�   �  
�  �    �     �  
�   �      D   ,  C   �  C  �  e  �  e   �  C   �      D   ,  �   �  �  �  �  �  �   �  �   �      D   ,  �   �  �  �    �     �  �   �      D   ,  -   �  -  �  O  �  O   �  -   �      D   ,  {   �  {  �  �  �  �   �  {   �      D   ,  �   �  �  �  �  �  �   �  �   �      D   ,     �    �  9  �  9   �     �      D   ,    N      �    �  N    N      D   ,���   ����  ����7  ����7   ����   �      D   ,���c   ����c  ����  ����   ����c   �      D   ,���   ����  �����  �����   ����   �      D   ,����   �����  ����!  ����!   �����   �      D   ,���M   ����M  ����o  ����o   ����M   �      D   ,���   ����  ����  ����   ����   �      D   ,����   �����  ����  ����   �����   �      D   ,���7   ����7  ����Y  ����Y   ����7   �      D   ,����   �����  �����  �����   �����   �      D   ,����   �����  �����  �����   �����   �      D   ,���!   ����!  ����C  ����C   ����!   �      D   ,���  N���  ���  ���  N���  N      D   ,���  N���  ����  ����  N���  N      D   ,���Z  N���Z  ���@  ���@  N���Z  N      D   ,���  N���  ���  ���  N���  N      D   ,����  N����  ����  ����  N����  N      D   ,���D  N���D  ���*  ���*  N���D  N      D   ,���  N���  ���x  ���x  N���  N      D   ,����  N����  ����  ����  N����  N      D   ,���.  N���.  ���  ���  N���.  N      D   ,���|  N���|  ���b  ���b  N���|  N      D   ,����  N����  ����  ����  N����  N      D   ,���  N���  ����  ����  N���  N      D   ,���f  N���f  ���L  ���L  N���f  N      D   ,����   �����  �����  �����   �����   �      D   ,������������e���7���e���7���������      D   ,���c������c���e������e���������c���      D   ,������������e�������e�������������      D   ,��������������e���!���e���!����������      D   ,���M������M���e���o���e���o������M���      D   ,������������e������e������������      D   ,��������������e������e�������������      D   ,���7������7���e���Y���e���Y������7���      D   ,��������������e�������e��������������      D   ,��������������e�������e��������������      D   ,���!������!���e���C���e���C������!���      D   ,��������������e�������e��������������      D   ,�����������������������������������      D   ,�������������������������������������      D   ,���Z�������Z�������@�������@�������Z����      D   ,�����������������������������������      D   ,����������������������������������������      D   ,���D�������D�������*�������*�������D����      D   ,�����������������x�������x�����������      D   ,����������������������������������������      D   ,���.�������.���������������������.����      D   ,���|�������|�������b�������b�������|����      D   ,����������������������������������������      D   ,�������������������������������������      D   ,���f�������f�������L�������L�������f����      D   ,  ���  ���e  -���e  -���  ���      D   ,  Y���  Y���e  {���e  {���  Y���      D   ,  ����  ����e  	����e  	����  ����      D   ,  
����  
����e  ���e  ���  
����      D   ,  C���  C���e  e���e  e���  C���      D   ,  ����  ����e  ����e  ����  ����      D   ,  ����  ����e  ���e  ���  ����      D   ,  -���  -���e  O���e  O���  -���      D   ,  {���  {���e  ����e  ����  {���      D   ,  ����  ����e  ����e  ����  ����      D   ,  ���  ���e  9���e  9���  ���      D   ,  ����  ����e  ����e  ����  ����      D   ,   �����   �����  �����  �����   �����      D   ,  ����  ����  �����  �����  ����      D   ,  P����  P����  6����  6����  P����      D   ,  �����  �����  �����  �����  �����      D   ,  	�����  	�����  
�����  
�����  	�����      D   ,  :����  :����   ����   ����  :����      D   ,  �����  �����  n����  n����  �����      D   ,  �����  �����  �����  �����  �����      D   ,  $����  $����  
����  
����  $����      D   ,  r����  r����  X����  X����  r����      D   ,  �����  �����  �����  �����  �����      D   ,  ����  ����  �����  �����  ����      D   ,  \����  \����  B����  B����  \����      @   ,�����������  M     M   ����������     �     "�     " "sky130_fd_pr__pfet_01v8_YC9MKB    �   ,���}�������}  	  �  	  ��������}����      A   ,���&���$���&  �  �  �  ����$���&���$      A  , ,���(  ����(  	o  �  	o  �  ����(  �      A  , ,���(���;���(  �����  ��������;���(���;      A  , ,  .���;  .  �  �  �  ����;  .���;      A  , ,���(�������(���;  ����;  ��������(����      ^   ,����������  Y  W  Y  W�����������      ]  , ,���  H���  	�  U  	�  U  H���  H      ]  , ,����������  H���O  H���O�����������      ]  , ,  �����  �  H  U  H  U����  �����      ]  , ,�������������  U����  U���������      B   ,���9  w���9  �����  �����  w���9  w      B   ,���  w���  �����  �����  w���  w      B   ,����  w����  ����  ����  w����  w      B   ,���#  w���#  ����m  ����m  w���#  w      B   ,���q  w���q  �����  �����  w���q  w      B   ,����  w����  ����	  ����	  w����  w      B   ,���  w���  ����W  ����W  w���  w      B   ,���[  w���[  �   �  �   �  w���[  w      B   ,  �  w  �  �  �  �  �  w  �  w      B   ,  �  w  �  �  A  �  A  w  �  w      B   ,  E  w  E  �  �  �  �  w  E  w      B   ,  �  w  �  �  	�  �  	�  w  �  w      B   ,  
�  w  
�  �  +  �  +  w  
�  w      B   ,  /  w  /  �  y  �  y  w  /  w      B   ,  }  w  }  �  �  �  �  w  }  w      B   ,���H�������H  w���t  w���t�������H����      B   ,����������  w����  w���������������      B   ,������������  w���  w���������������      B   ,���2�������2  w���^  w���^�������2����      B   ,������������  w����  w����������������      B   ,������������  w����  w����������������      B   ,����������  w���H  w���H�����������      B   ,���j�������j  w   �  w   ��������j����      B   ,  �����  �  w  �  w  �����  �����      B   ,  ����    w  2  w  2����  ����      B   ,  T����  T  w  �  w  �����  T����      B   ,  �����  �  w  	�  w  	�����  �����      B   ,  
�����  
�  w    w  ����  
�����      B   ,  >����  >  w  j  w  j����  >����      B   ,  �����  �  w  �  w  �����  �����      B   ,���9���?���9�������������������?���9���?      B   ,������?����������������������?������?      B   ,�������?���������������������?�������?      B   ,���#���?���#�������m�������m���?���#���?      B   ,���q���?���q�������������������?���q���?      B   ,�������?�����������	�������	���?�������?      B   ,������?����������W�������W���?������?      B   ,���[���?���[����   �����   ����?���[���?      B   ,  ����?  �����  �����  ����?  ����?      B   ,  ����?  �����  A����  A���?  ����?      B   ,  E���?  E����  �����  ����?  E���?      B   ,  ����?  �����  	�����  	����?  ����?      B   ,  
����?  
�����  +����  +���?  
����?      B   ,  /���?  /����  y����  y���?  /���?      B   ,  }���?  }����  �����  ����?  }���?      B  , ,����  �����  	o   U  	o   U  �����  �      B  , ,����  �����  q   U  q   U  �����  �      B  , ,���(�������(   U����   U�����������(����      B  , ,  .����  .   U  �   U  �����  .����      B  , ,���������������9   U���9   U������������      B  , ,���������������;   U���;   U������������      B  , ,  �  �  �  	o  M  	o  M  �  �  �      B  , ,  �  �  �  	o  	�  	o  	�  �  �  �      B  , ,  
K  �  
K  	o  
�  	o  
�  �  
K  �      B  , ,  �  �  �  	o  I  	o  I  �  �  �      B  , ,  �  �  �  	o  �  	o  �  �  �  �      B  , ,  G  �  G  	o  �  	o  �  �  G  �      B  , ,  �  �  �  	o  E  	o  E  �  �  �      B  , ,  �  �  �  	o  �  	o  �  �  �  �      B  , ,   �  �   �  	o  �  	o  �  �   �  �      B  , ,  �  �  �  q  �  q  �  �  �  �      B  , ,  G  �  G  q  �  q  �  �  G  �      B  , ,  �  �  �  q  ?  q  ?  �  �  �      B  , ,  �  �  �  q  	�  q  	�  �  �  �      B  , ,  1  �  1  q  �  q  �  �  1  �      B  , ,    �    q  )  q  )  �    �      B  , ,  �  �  �  q  w  q  w  �  �  �      B  , ,  .  O  .  �  �  �  �  O  .  O      B  , ,  .  �  .  �  �  �  �  �  .  �      B  , ,   �  Q   �  �  |  �  |  Q   �  Q      B  , ,     Q     �  �  �  �  Q     Q      B  , ,  n  Q  n  �    �    Q  n  Q      B  , ,  �  Q  �  �  f  �  f  Q  �  Q      B  , ,  

  Q  

  �  
�  �  
�  Q  

  Q      B  , ,  X  Q  X  �    �    Q  X  Q      B  , ,  �  Q  �  �  P  �  P  Q  �  Q      B  , ,  �  Q  �  �  �  �  �  Q  �  Q      B  , ,  .  �  .  Q  �  Q  �  �  .  �      B  , ,   �  �   �  �  |  �  |  �   �  �      B  , ,     �     �  �  �  �  �     �      B  , ,  n  �  n  �    �    �  n  �      B  , ,  �  �  �  �  f  �  f  �  �  �      B  , ,  

  �  

  �  
�  �  
�  �  

  �      B  , ,  X  �  X  �    �    �  X  �      B  , ,  �  �  �  �  P  �  P  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  .  S  .  �  �  �  �  S  .  S      B  , ,   �  �   �  S  |  S  |  �   �  �      B  , ,     �     S  �  S  �  �     �      B  , ,  n  �  n  S    S    �  n  �      B  , ,  �  �  �  S  f  S  f  �  �  �      B  , ,  

  �  

  S  
�  S  
�  �  

  �      B  , ,  X  �  X  S    S    �  X  �      B  , ,  �  �  �  S  P  S  P  �  �  �      B  , ,  �  �  �  S  �  S  �  �  �  �      B  , ,  .   �  .  �  �  �  �   �  .   �      B  , ,   �   U   �   �  |   �  |   U   �   U      B  , ,      U      �  �   �  �   U      U      B  , ,  n   U  n   �     �     U  n   U      B  , ,  �   U  �   �  f   �  f   U  �   U      B  , ,  

   U  

   �  
�   �  
�   U  

   U      B  , ,  X   U  X   �     �     U  X   U      B  , ,  �   U  �   �  P   �  P   U  �   U      B  , ,  �   U  �   �  �   �  �   U  �   U      B  , ,  S  �  S  	o  �  	o  �  �  S  �      B  , ,  �  �  �  	o  Q  	o  Q  �  �  �      B  , ,  �  �  �  	o  �  	o  �  �  �  �      B  , ,  O  �  O  	o  �  	o  �  �  O  �      B  , ,����  �����  q���k  q���k  �����  �      B  , ,���b  ����b  ����  ����  ����b  �      B  , ,���  ����  ����Z  ����Z  ����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,���L  ����L  �����  �����  ����L  �      B  , ,����  �����  ����D  ����D  �����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,���6  ����6  �����  �����  ����6  �      B  , ,����  �����  ����.  ����.  �����  �      B  , ,���  ����  q����  q����  ����  �      B  , ,���]  ����]  q���  q���  ����]  �      B  , ,���  ����  	o���e  	o���e  ����  �      B  , ,���  ����  	o���  	o���  ����  �      B  , ,���c  ����c  	o���  	o���  ����c  �      B  , ,���  ����  	o���a  	o���a  ����  �      B  , ,���  ����  	o����  	o����  ����  �      B  , ,���_  ����_  	o���	  	o���	  ����_  �      B  , ,���(  S���(  �����  �����  S���(  S      B  , ,����  �����  	o���]  	o���]  �����  �      B  , ,���b  ����b  S���  S���  ����b  �      B  , ,���  ����  S���Z  S���Z  ����  �      B  , ,����  �����  S���  S���  �����  �      B  , ,���L  ����L  S����  S����  ����L  �      B  , ,����  �����  S���D  S���D  �����  �      B  , ,����  �����  S����  S����  �����  �      B  , ,���6  ����6  S����  S����  ����6  �      B  , ,����  �����  S���.  S���.  �����  �      B  , ,���  ����  	o����  	o����  ����  �      B  , ,���[  ����[  	o���  	o���  ����[  �      B  , ,���(  ����(  �����  �����  ����(  �      B  , ,����  �����  	o���Y  	o���Y  �����  �      B  , ,���b  Q���b  ����  ����  Q���b  Q      B  , ,���  Q���  ����Z  ����Z  Q���  Q      B  , ,����  Q����  ����  ����  Q����  Q      B  , ,���L  Q���L  �����  �����  Q���L  Q      B  , ,���(   ����(  �����  �����   ����(   �      B  , ,����  Q����  ����D  ����D  Q����  Q      B  , ,���b   U���b   ����   ����   U���b   U      B  , ,���   U���   ����Z   ����Z   U���   U      B  , ,����   U����   ����   ����   U����   U      B  , ,���L   U���L   �����   �����   U���L   U      B  , ,����   U����   ����D   ����D   U����   U      B  , ,����   U����   �����   �����   U����   U      B  , ,���6   U���6   �����   �����   U���6   U      B  , ,����   U����   ����.   ����.   U����   U      B  , ,����  Q����  �����  �����  Q����  Q      B  , ,���6  Q���6  �����  �����  Q���6  Q      B  , ,����  Q����  ����.  ����.  Q����  Q      B  , ,���  ����  	o����  	o����  ����  �      B  , ,���W  ����W  	o���  	o���  ����W  �      B  , ,���g  ����g  	o���  	o���  ����g  �      B  , ,���(  O���(  �����  �����  O���(  O      B  , ,���  ����  q���3  q���3  ����  �      B  , ,����  �����  q���  q���  �����  �      B  , ,���%  ����%  q����  q����  ����%  �      B  , ,���s  ����s  q���  q���  ����s  �      B  , ,���(  ����(  Q����  Q����  ����(  �      B  , ,�����������������������������������      B  , ,���L������L����������������������L���      B  , ,������������������D�������D����������      B  , ,�������������������������������������      B  , ,���6������6����������������������6���      B  , ,������������������.�������.����������      B  , ,���(���W���(�����������������W���(���W      B  , ,���b�������b���W������W����������b����      B  , ,�������������W���Z���W���Z�����������      B  , ,���������������W������W���������������      B  , ,���L�������L���W�������W�����������L����      B  , ,���������������W���D���W���D������������      B  , ,���������������W�������W����������������      B  , ,���6�������6���W�������W�����������6����      B  , ,���������������W���.���W���.������������      B  , ,���(������(����������������������(���      B  , ,���b���Y���b���������������Y���b���Y      B  , ,������Y���������Z������Z���Y������Y      B  , ,�������Y�������������������Y�������Y      B  , ,���L���Y���L�����������������Y���L���Y      B  , ,�������Y����������D������D���Y�������Y      B  , ,�������Y���������������������Y�������Y      B  , ,���6���Y���6�����������������Y���6���Y      B  , ,�������Y����������.������.���Y�������Y      B  , ,���(�������(���Y�������Y�����������(����      B  , ,���b������b��������������������b���      B  , ,����������������Z�������Z���������      B  , ,�����������������������������������      B  , ,���L������L����������������������L���      B  , ,������������������D�������D����������      B  , ,�������������������������������������      B  , ,���6������6����������������������6���      B  , ,������������������.�������.����������      B  , ,���(���[���(�����������������[���(���[      B  , ,���(������(����������������������(���      B  , ,�������������9���3���9���3�����������      B  , ,���������������9������9���������������      B  , ,���%�������%���9�������9�����������%����      B  , ,���s�������s���9������9����������s����      B  , ,���������������9���k���9���k������������      B  , ,�������������9�������9���������������      B  , ,���]�������]���9������9����������]����      B  , ,���b������b��������������������b���      B  , ,���g�������g���;������;����������g����      B  , ,�������������;���e���;���e�����������      B  , ,�������������;������;��������������      B  , ,���c�������c���;������;����������c����      B  , ,�������������;���a���;���a�����������      B  , ,�������������;�������;���������������      B  , ,���_�������_���;���	���;���	�������_����      B  , ,���������������;���]���;���]������������      B  , ,�������������;�������;���������������      B  , ,���[�������[���;������;����������[����      B  , ,���������������;���Y���;���Y������������      B  , ,�������������;�������;���������������      B  , ,���W�������W���;������;����������W����      B  , ,����������������Z�������Z���������      B  , ,  �����  ����W  P���W  P����  �����      B  , ,  �����  ����W  ����W  �����  �����      B  , ,  .���W  .���  ����  ����W  .���W      B  , ,   ����   �����  |����  |���   ����      B  , ,   ���   ����  �����  ����   ���      B  , ,  n���  n����  ����  ���  n���      B  , ,  ����  �����  f����  f���  ����      B  , ,  

���  

����  
�����  
����  

���      B  , ,  X���  X����  ����  ���  X���      B  , ,  ����  �����  P����  P���  ����      B  , ,  ����  �����  �����  ����  ����      B  , ,  .���  .����  �����  ����  .���      B  , ,  .���[  .���  ����  ����[  .���[      B  , ,   ���   ����  �����  ����   ���      B  , ,  n���  n����  ����  ���  n���      B  , ,  ����  �����  f����  f���  ����      B  , ,  

���  

����  
�����  
����  

���      B  , ,  X���  X����  ����  ���  X���      B  , ,  ����  �����  P����  P���  ����      B  , ,  ����  �����  �����  ����  ����      B  , ,   ����   �����  |����  |���   ����      B  , ,   ����Y   ����  |���  |���Y   ����Y      B  , ,  �����  ����9  ����9  �����  �����      B  , ,  G����  G���9  ����9  �����  G����      B  , ,  �����  ����9  ?���9  ?����  �����      B  , ,  �����  ����9  	����9  	�����  �����      B  , ,  1����  1���9  ����9  �����  1����      B  , ,  ����  ���9  )���9  )����  ����      B  , ,  �����  ����9  w���9  w����  �����      B  , ,  .���  .����  �����  ����  .���      B  , ,   ���Y   ���  ����  ����Y   ���Y      B  , ,  n���Y  n���  ���  ���Y  n���Y      B  , ,  ����Y  ����  f���  f���Y  ����Y      B  , ,  

���Y  

���  
����  
����Y  

���Y      B  , ,  X���Y  X���  ���  ���Y  X���Y      B  , ,  ����Y  ����  P���  P���Y  ����Y      B  , ,  ����Y  ����  ����  ����Y  ����Y      B  , ,   �����   ����W  |���W  |����   �����      B  , ,  .����  .���Y  ����Y  �����  .����      B  , ,   ����   ���W  ����W  �����   ����      B  , ,  n����  n���W  ���W  ����  n����      B  , ,  �����  ����W  f���W  f����  �����      B  , ,  

����  

���W  
����W  
�����  

����      B  , ,  X����  X���W  ���W  ����  X����      B  , ,   �����   ����;  ����;  �����   �����      B  , ,  S����  S���;  ����;  �����  S����      B  , ,  �����  ����;  Q���;  Q����  �����      B  , ,  �����  ����;  ����;  �����  �����      B  , ,  O����  O���;  ����;  �����  O����      B  , ,  �����  ����;  M���;  M����  �����      B  , ,  �����  ����;  	����;  	�����  �����      B  , ,  
K����  
K���;  
����;  
�����  
K����      B  , ,  �����  ����;  I���;  I����  �����      B  , ,  �����  ����;  ����;  �����  �����      B  , ,  G����  G���;  ����;  �����  G����      B  , ,  �����  ����;  E���;  E����  �����      B  , ,  �����  ����;  ����;  �����  �����      _   ,���%  c���%  �  �  �  �  c���%  c      _   ,���%���+���%����  �����  ����+���%���+      C   ,���(  ����(  	o  �  	o  �  ����(  �      C   ,���(���;���(  �����  ��������;���(���;      C   ,���9  ����9  q����  q����  ����9  �      C   ,���  ����  q����  q����  ����  �      C   ,����  �����  q���  q���  �����  �      C   ,���#  ����#  q���m  q���m  ����#  �      C   ,���q  ����q  q����  q����  ����q  �      C   ,����  �����  q���	  q���	  �����  �      C   ,���  ����  q���W  q���W  ����  �      C   ,���[  ����[  q   �  q   �  ����[  �      C   ,  �  �  �  q  �  q  �  �  �  �      C   ,  �  �  �  q  A  q  A  �  �  �      C   ,  E  �  E  q  �  q  �  �  E  �      C   ,  �  �  �  q  	�  q  	�  �  �  �      C   ,  
�  �  
�  q  +  q  +  �  
�  �      C   ,  /  �  /  q  y  q  y  �  /  �      C   ,  }  �  }  q  �  q  �  �  }  �      C   ,���b������b  ����  ����������b���      C   ,���������  ����Z  ����Z���������      C   ,�����������  ����  ��������������      C   ,���L������L  �����  �����������L���      C   ,�����������  ����D  ����D����������      C   ,�����������  �����  ���������������      C   ,���6������6  �����  �����������6���      C   ,�����������  ����.  ����.����������      C   ,   ����   �  �  |  �  |���   ����      C   ,   ���     �  �  �  ����   ���      C   ,  n���  n  �    �  ���  n���      C   ,  ����  �  �  f  �  f���  ����      C   ,  

���  

  �  
�  �  
����  

���      C   ,  X���  X  �    �  ���  X���      C   ,  ����  �  �  P  �  P���  ����      C   ,  ����  �  �  �  �  ����  ����      C   ,���9�������9���9�������9�����������9����      C   ,�������������9�������9���������������      C   ,���������������9������9���������������      C   ,���#�������#���9���m���9���m�������#����      C   ,���q�������q���9�������9�����������q����      C   ,���������������9���	���9���	������������      C   ,�������������9���W���9���W�����������      C   ,���[�������[���9   ����9   ��������[����      C   ,  �����  ����9  ����9  �����  �����      C   ,  �����  ����9  A���9  A����  �����      C   ,  E����  E���9  ����9  �����  E����      C   ,  �����  ����9  	����9  	�����  �����      C   ,  
�����  
����9  +���9  +����  
�����      C   ,  /����  /���9  y���9  y����  /����      C   ,  }����  }���9  ����9  �����  }����      C   ,  .���;  .  �  �  �  ����;  .���;      C   ,���(�������(���;  ����;  ��������(����      C  , ,����  �����  q   U  q   U  �����  �      C  , ,���������������9   U���9   U������������      C  , ,  G  �  G  q  �  q  �  �  G  �      C  , ,  �  �  �  q  ?  q  ?  �  �  �      C  , ,  �  �  �  q  	�  q  	�  �  �  �      C  , ,  1  �  1  q  �  q  �  �  1  �      C  , ,    �    q  )  q  )  �    �      C  , ,  �  �  �  q  w  q  w  �  �  �      C  , ,   �  �   �  A  |  A  |  �   �  �      C  , ,     �     A  �  A  �  �     �      C  , ,  n  �  n  A    A    �  n  �      C  , ,  �  �  �  A  f  A  f  �  �  �      C  , ,  

  �  

  A  
�  A  
�  �  

  �      C  , ,  X  �  X  A    A    �  X  �      C  , ,  �  �  �  A  P  A  P  �  �  �      C  , ,  �  �  �  A  �  A  �  �  �  �      C  , ,   �  /   �  �  |  �  |  /   �  /      C  , ,     /     �  �  �  �  /     /      C  , ,  n  /  n  �    �    /  n  /      C  , ,  �  /  �  �  f  �  f  /  �  /      C  , ,  

  /  

  �  
�  �  
�  /  

  /      C  , ,  X  /  X  �    �    /  X  /      C  , ,  �  /  �  �  P  �  P  /  �  /      C  , ,  �  /  �  �  �  �  �  /  �  /      C  , ,   �  �   �  q  |  q  |  �   �  �      C  , ,     �     q  �  q  �  �     �      C  , ,  n  �  n  q    q    �  n  �      C  , ,  �  �  �  q  f  q  f  �  �  �      C  , ,  

  �  

  q  
�  q  
�  �  

  �      C  , ,  X  �  X  q    q    �  X  �      C  , ,  �  �  �  q  P  q  P  �  �  �      C  , ,  �  �  �  q  �  q  �  �  �  �      C  , ,   �   _   �  	  |  	  |   _   �   _      C  , ,      _     	  �  	  �   _      _      C  , ,  n   _  n  	    	     _  n   _      C  , ,  �   _  �  	  f  	  f   _  �   _      C  , ,  

   _  

  	  
�  	  
�   _  

   _      C  , ,  X   _  X  	    	     _  X   _      C  , ,  �   _  �  	  P  	  P   _  �   _      C  , ,  �   _  �  	  �  	  �   _  �   _      C  , ,  �  �  �  q  �  q  �  �  �  �      C  , ,���L  ����L  A����  A����  ����L  �      C  , ,����  �����  A���D  A���D  �����  �      C  , ,����  �����  A����  A����  �����  �      C  , ,���6  ����6  A����  A����  ����6  �      C  , ,����  �����  A���.  A���.  �����  �      C  , ,����  �����  q���  q���  �����  �      C  , ,���b  ����b  q���  q���  ����b  �      C  , ,���  ����  q���Z  q���Z  ����  �      C  , ,����  �����  q���  q���  �����  �      C  , ,���L  ����L  q����  q����  ����L  �      C  , ,����  �����  q���D  q���D  �����  �      C  , ,����  �����  q����  q����  �����  �      C  , ,���6  ����6  q����  q����  ����6  �      C  , ,����  �����  q���.  q���.  �����  �      C  , ,���%  ����%  q����  q����  ����%  �      C  , ,���s  ����s  q���  q���  ����s  �      C  , ,����  �����  q���k  q���k  �����  �      C  , ,���  ����  q����  q����  ����  �      C  , ,���]  ����]  q���  q���  ����]  �      C  , ,���  ����  q���3  q���3  ����  �      C  , ,���b  ����b  A���  A���  ����b  �      C  , ,���b  /���b  ����  ����  /���b  /      C  , ,���b   _���b  	���  	���   _���b   _      C  , ,���   _���  	���Z  	���Z   _���   _      C  , ,����   _����  	���  	���   _����   _      C  , ,���L   _���L  	����  	����   _���L   _      C  , ,����   _����  	���D  	���D   _����   _      C  , ,����   _����  	����  	����   _����   _      C  , ,���6   _���6  	����  	����   _���6   _      C  , ,����   _����  	���.  	���.   _����   _      C  , ,���  /���  ����Z  ����Z  /���  /      C  , ,����  /����  ����  ����  /����  /      C  , ,���L  /���L  �����  �����  /���L  /      C  , ,����  /����  ����D  ����D  /����  /      C  , ,����  /����  �����  �����  /����  /      C  , ,���6  /���6  �����  �����  /���6  /      C  , ,����  /����  ����.  ����.  /����  /      C  , ,���  ����  A���Z  A���Z  ����  �      C  , ,����  �����  A���  A���  �����  �      C  , ,�����������������Z�������Z�����������      C  , ,��������������������������������������      C  , ,���L�������L�����������������������L����      C  , ,�������������������D�������D������������      C  , ,����������������������������������������      C  , ,���6�������6�����������������������6����      C  , ,�������������������.�������.������������      C  , ,���b�������b���9������9����������b����      C  , ,�������������9���Z���9���Z�����������      C  , ,���������������9������9���������������      C  , ,���L�������L���9�������9�����������L����      C  , ,���������������9���D���9���D������������      C  , ,���������������9�������9����������������      C  , ,���6�������6���9�������9�����������6����      C  , ,���������������9���.���9���.������������      C  , ,���b���'���b�����������������'���b���'      C  , ,������'����������Z�������Z���'������'      C  , ,�������'���������������������'�������'      C  , ,���L���'���L�������������������'���L���'      C  , ,�������'�����������D�������D���'�������'      C  , ,�������'�����������������������'�������'      C  , ,���6���'���6�������������������'���6���'      C  , ,�������'�����������.�������.���'�������'      C  , ,���b�������b���i������i����������b����      C  , ,�������������i���Z���i���Z�����������      C  , ,���������������i������i���������������      C  , ,���L�������L���i�������i�����������L����      C  , ,���������������i���D���i���D������������      C  , ,���������������i�������i����������������      C  , ,���6�������6���i�������i�����������6����      C  , ,���������������i���.���i���.������������      C  , ,�������������9���3���9���3�����������      C  , ,���������������9������9���������������      C  , ,���%�������%���9�������9�����������%����      C  , ,���s�������s���9������9����������s����      C  , ,���������������9���k���9���k������������      C  , ,�������������9�������9���������������      C  , ,���]�������]���9������9����������]����      C  , ,���b�������b���������������������b����      C  , ,   ����'   �����  |����  |���'   ����'      C  , ,   ���'   ����  �����  ����'   ���'      C  , ,  n���'  n����  ����  ���'  n���'      C  , ,  ����'  �����  f����  f���'  ����'      C  , ,  

���'  

����  
�����  
����'  

���'      C  , ,  X���'  X����  ����  ���'  X���'      C  , ,  ����'  �����  P����  P���'  ����'      C  , ,  ����'  �����  �����  ����'  ����'      C  , ,   �����   ����9  |���9  |����   �����      C  , ,   ����   ���9  ����9  �����   ����      C  , ,  n����  n���9  ���9  ����  n����      C  , ,  �����  ����9  f���9  f����  �����      C  , ,  

����  

���9  
����9  
�����  

����      C  , ,  X����  X���9  ���9  ����  X����      C  , ,  �����  ����9  P���9  P����  �����      C  , ,  �����  ����9  ����9  �����  �����      C  , ,   �����   ����i  |���i  |����   �����      C  , ,   ����   ���i  ����i  �����   ����      C  , ,  n����  n���i  ���i  ����  n����      C  , ,  �����  ����i  f���i  f����  �����      C  , ,  

����  

���i  
����i  
�����  

����      C  , ,  X����  X���i  ���i  ����  X����      C  , ,  �����  ����i  P���i  P����  �����      C  , ,  �����  ����i  ����i  �����  �����      C  , ,   �����   �����  |����  |����   �����      C  , ,   ����   ����  �����  �����   ����      C  , ,  n����  n����  ����  ����  n����      C  , ,  �����  �����  f����  f����  �����      C  , ,  

����  

����  
�����  
�����  

����      C  , ,  X����  X����  ����  ����  X����      C  , ,  �����  �����  P����  P����  �����      C  , ,  �����  �����  �����  �����  �����      C  , ,  �����  ����9  ����9  �����  �����      C  , ,  G����  G���9  ����9  �����  G����      C  , ,  �����  ����9  ?���9  ?����  �����      C  , ,  �����  ����9  	����9  	�����  �����      C  , ,  1����  1���9  ����9  �����  1����      C  , ,  ����  ���9  )���9  )����  ����      C  , ,  �����  ����9  w���9  w����  �����      D   ,���M  ����M  ����o  ����o  ����M  �      D   ,���  ����  ����  ����  ����  �      D   ,����  �����  ����  ����  �����  �      D   ,���7  ����7  ����Y  ����Y  ����7  �      D   ,����  �����  �����  �����  �����  �      D   ,����  �����  �����  �����  �����  �      D   ,���!  ����!  ����C  ����C  ����!  �      D   ,���o  ����o  �   �  �   �  ����o  �      D   ,  �  �  �  �  �  �  �  �  �  �      D   ,    �    �  -  �  -  �    �      D   ,  Y  �  Y  �  {  �  {  �  Y  �      D   ,  �  �  �  �  	�  �  	�  �  �  �      D   ,  
�  �  
�  �    �    �  
�  �      D   ,  C  �  C  �  e  �  e  �  C  �      D   ,  �  �  �  �  �  �  �  �  �  �      D   ,���D���$���D  ����*  ����*���$���D���$      D   ,������$���  ����x  ����x���$������$      D   ,�������$����  �����  ��������$�������$      D   ,���.���$���.  ����  �������$���.���$      D   ,���|���$���|  ����b  ����b���$���|���$      D   ,�������$����  �����  ��������$�������$      D   ,������$���  �����  ��������$������$      D   ,���f���$���f  ����L  ����L���$���f���$      D   ,   ����$   �  �  �  �  ����$   ����$      D   ,  ���$    �  �  �  ����$  ���$      D   ,  P���$  P  �  6  �  6���$  P���$      D   ,  ����$  �  �  �  �  ����$  ����$      D   ,  	����$  	�  �  
�  �  
����$  	����$      D   ,  :���$  :  �     �   ���$  :���$      D   ,  ����$  �  �  n  �  n���$  ����$      D   ,  ����$  �  �  �  �  ����$  ����$      D   ,���M���q���M���W���o���W���o���q���M���q      D   ,������q������W������W������q������q      D   ,�������q�������W������W������q�������q      D   ,���7���q���7���W���Y���W���Y���q���7���q      D   ,�������q�������W�������W�������q�������q      D   ,�������q�������W�������W�������q�������q      D   ,���!���q���!���W���C���W���C���q���!���q      D   ,���o���q���o���W   ����W   ����q���o���q      D   ,  ����q  ����W  ����W  ����q  ����q      D   ,  ���q  ���W  -���W  -���q  ���q      D   ,  Y���q  Y���W  {���W  {���q  Y���q      D   ,  ����q  ����W  	����W  	����q  ����q      D   ,  
����q  
����W  ���W  ���q  
����q      D   ,  C���q  C���W  e���W  e���q  C���q      D   ,  ����q  ����W  ����W  ����q  ����q      @   ,���t�������t  
#  �  
#  ��������t����     �     "�     " "sky130_fd_pr__nfet_01v8_8JUMX6    �   ,���`���:���`  �  n�  �  n����:���`���:      A   ,���	  !���	  �  l�  �  l�  !���	  !      A   ,���	���K���	����  l�����  l����K���	���K      A  , ,���  q���    n�    n�  q���  q      A  , ,���������  q����  q�������������      A  , ,  nK���  nK  q  n�  q  n����  nK���      A  , ,�������������  n����  n������������      ^   ,����  �����  �  or  �  or  �����  �      ^   ,�����������  ����2  ����2����������      ^   ,  m����  m�  �  or  �  or���  m����      ^   ,�������h�������  or���  or���h�������h      ]  , ,����  �����  2  mt  2  mt  �����  �      ]  , ,���������������\  mt���\  mt������������      B   ,���   i���  m   �  m   �   i���   i      B   ,�������������   �����   ����������      B   ,  �   i  �  m  �  m  �   i  �   i      B   ,  �   i  �  m  	�  m  	�   i  �   i      B   ,  
�   i  
�  m  q  m  q   i  
�   i      B   ,  �   i  �  m  U  m  U   i  �   i      B   ,  w   i  w  m  9  m  9   i  w   i      B   ,  [   i  [  m    m     i  [   i      B   ,  ?   i  ?  m    m     i  ?   i      B   ,  #   i  #  m  �  m  �   i  #   i      B   ,     i    m  �  m  �   i     i      B   ,  �   i  �  m   �  m   �   i  �   i      B   ,  !�   i  !�  m  #�  m  #�   i  !�   i      B   ,  $�   i  $�  m  &u  m  &u   i  $�   i      B   ,  '�   i  '�  m  )Y  m  )Y   i  '�   i      B   ,  *{   i  *{  m  ,=  m  ,=   i  *{   i      B   ,  -_   i  -_  m  /!  m  /!   i  -_   i      B   ,  0C   i  0C  m  2  m  2   i  0C   i      B   ,  3'   i  3'  m  4�  m  4�   i  3'   i      B   ,  6   i  6  m  7�  m  7�   i  6   i      B   ,  8�   i  8�  m  :�  m  :�   i  8�   i      B   ,  ;�   i  ;�  m  =�  m  =�   i  ;�   i      B   ,  >�   i  >�  m  @y  m  @y   i  >�   i      B   ,  A�   i  A�  m  C]  m  C]   i  A�   i      B   ,  D   i  D  m  FA  m  FA   i  D   i      B   ,  Gc   i  Gc  m  I%  m  I%   i  Gc   i      B   ,  JG   i  JG  m  L	  m  L	   i  JG   i      B   ,  M+   i  M+  m  N�  m  N�   i  M+   i      B   ,  P   i  P  m  Q�  m  Q�   i  P   i      B   ,  R�   i  R�  m  T�  m  T�   i  R�   i      B   ,  U�   i  U�  m  W�  m  W�   i  U�   i      B   ,  X�   i  X�  m  Z}  m  Z}   i  X�   i      B   ,  [�   i  [�  m  ]a  m  ]a   i  [�   i      B   ,  ^�   i  ^�  m  `E  m  `E   i  ^�   i      B   ,  ag   i  ag  m  c)  m  c)   i  ag   i      B   ,  dK   i  dK  m  f  m  f   i  dK   i      B   ,  g/   i  g/  m  h�  m  h�   i  g/   i      B   ,  j   i  j  m  k�  m  k�   i  j   i      B   ,     i    m  �  m  �   i     i      B   ,����   i����  m����  m����   i����   i      B   ,����   i����  m����  m����   i����   i      B   ,����   i����  m���}  m���}   i����   i      B   ,����   i����  m���a  m���a   i����   i      B   ,����   i����  m���E  m���E   i����   i      B   ,���g   i���g  m���)  m���)   i���g   i      B   ,���K   i���K  m���  m���   i���K   i      B   ,���/   i���/  m����  m����   i���/   i      B   ,���   i���  m����  m����   i���   i      B   ,����   i����  m����  m����   i����   i      B   ,����   i����  m����  m����   i����   i      B   ,����   i����  m����  m����   i����   i      B   ,����   i����  m���e  m���e   i����   i      B   ,����   i����  m���I  m���I   i����   i      B   ,���k   i���k  m���-  m���-   i���k   i      B   ,���O   i���O  m���  m���   i���O   i      B   ,���3   i���3  m����  m����   i���3   i      B   ,���   i���  m����  m����   i���   i      B   ,����   i����  m��Ͻ  m��Ͻ   i����   i      B   ,����   i����  m��ҡ  m��ҡ   i����   i      B   ,����   i����  m��Յ  m��Յ   i����   i      B   ,��֧   i��֧  m���i  m���i   i��֧   i      B   ,��ً   i��ً  m���M  m���M   i��ً   i      B   ,���o   i���o  m���1  m���1   i���o   i      B   ,���S   i���S  m���  m���   i���S   i      B   ,���7   i���7  m����  m����   i���7   i      B   ,���   i���  m����  m����   i���   i      B   ,����   i����  m����  m����   i����   i      B   ,����   i����  m���  m���   i����   i      B   ,����   i����  m���  m���   i����   i      B   ,���   i���  m���m  m���m   i���   i      B   ,���   i���  m���Q  m���Q   i���   i      B   ,���s   i���s  m���5  m���5   i���s   i      B   ,���W   i���W  m���  m���   i���W   i      B   ,���;   i���;  m����  m����   i���;   i      B   ,���+   i���+  m����  m����   i���+   i      B   ,���   i���  m����  m����   i���   i      B   ,����������������������������������      B   ,�������������������������������������      B   ,�������������������������������������      B   ,������������������}�������}����������      B   ,������������������a�������a����������      B   ,������������������E�������E����������      B   ,���g������g�������)�������)������g���      B   ,���K������K��������������������K���      B   ,���/������/����������������������/���      B   ,����������������������������������      B   ,�������������������������������������      B   ,�������������������������������������      B   ,�������������������������������������      B   ,������������������e�������e����������      B   ,������������������I�������I����������      B   ,���k������k�������-�������-������k���      B   ,���O������O��������������������O���      B   ,���3������3����������������������3���      B   ,����������������������������������      B   ,�����������������Ͻ������Ͻ����������      B   ,�����������������ҡ������ҡ����������      B   ,�����������������Յ������Յ����������      B   ,��֧�����֧�������i�������i�����֧���      B   ,��ً�����ً�������M�������M�����ً���      B   ,���o������o�������1�������1������o���      B   ,���S������S��������������������S���      B   ,���7������7����������������������7���      B   ,����������������������������������      B   ,�������������������������������������      B   ,�����������������������������������      B   ,�����������������������������������      B   ,����������������m�������m���������      B   ,����������������Q�������Q���������      B   ,���s������s�������5�������5������s���      B   ,���W������W��������������������W���      B   ,���;������;����������������������;���      B   ,���+������+����������������������+���      B   ,  ���  ����  �����  ����  ���      B   ,  ����  �����  �����  ����  ����      B   ,  ����  �����  	�����  	����  ����      B   ,  
����  
�����  q����  q���  
����      B   ,  ����  �����  U����  U���  ����      B   ,  w���  w����  9����  9���  w���      B   ,  [���  [����  ����  ���  [���      B   ,  ?���  ?����  ����  ���  ?���      B   ,  #���  #����  �����  ����  #���      B   ,  ���  ����  �����  ����  ���      B   ,  ����  �����   �����   ����  ����      B   ,  !����  !�����  #�����  #����  !����      B   ,  $����  $�����  &u����  &u���  $����      B   ,  '����  '�����  )Y����  )Y���  '����      B   ,  *{���  *{����  ,=����  ,=���  *{���      B   ,  -_���  -_����  /!����  /!���  -_���      B   ,  0C���  0C����  2����  2���  0C���      B   ,  3'���  3'����  4�����  4����  3'���      B   ,  6���  6����  7�����  7����  6���      B   ,  8����  8�����  :�����  :����  8����      B   ,  ;����  ;�����  =�����  =����  ;����      B   ,  >����  >�����  @y����  @y���  >����      B   ,  A����  A�����  C]����  C]���  A����      B   ,  D���  D����  FA����  FA���  D���      B   ,  Gc���  Gc����  I%����  I%���  Gc���      B   ,  JG���  JG����  L	����  L	���  JG���      B   ,  M+���  M+����  N�����  N����  M+���      B   ,  P���  P����  Q�����  Q����  P���      B   ,  R����  R�����  T�����  T����  R����      B   ,  U����  U�����  W�����  W����  U����      B   ,  X����  X�����  Z}����  Z}���  X����      B   ,  [����  [�����  ]a����  ]a���  [����      B   ,  ^����  ^�����  `E����  `E���  ^����      B   ,  ag���  ag����  c)����  c)���  ag���      B   ,  dK���  dK����  f����  f���  dK���      B   ,  g/���  g/����  h�����  h����  g/���      B   ,  j���  j����  k�����  k����  j���      B  , ,����  s����     U     U  s����  s      B  , ,����   �����  c   U  c   U   �����   �      B  , ,���������������G   U���G   U������������      B  , ,���������������   U���   U������������      B  , ,  nK  
�  nK  �  n�  �  n�  
�  nK  
�      B  , ,  R�  q  R�    SW    SW  q  R�  q      B  , ,  8	  :  8	  �  8�  �  8�  :  8	  :      B  , ,  :�  :  :�  �  ;�  �  ;�  :  :�  :      B  , ,  =�  :  =�  �  >{  �  >{  :  =�  :      B  , ,  @�  :  @�  �  A_  �  A_  :  @�  :      B  , ,  C�  :  C�  �  DC  �  DC  :  C�  :      B  , ,  F}  :  F}  �  G'  �  G'  :  F}  :      B  , ,  Ia  :  Ia  �  J  �  J  :  Ia  :      B  , ,  LE  :  LE  �  L�  �  L�  :  LE  :      B  , ,  O)  :  O)  �  O�  �  O�  :  O)  :      B  , ,  R  :  R  �  R�  �  R�  :  R  :      B  , ,  T�  :  T�  �  U�  �  U�  :  T�  :      B  , ,  W�  :  W�  �  X  �  X  :  W�  :      B  , ,  Z�  :  Z�  �  [c  �  [c  :  Z�  :      B  , ,  ]�  :  ]�  �  ^G  �  ^G  :  ]�  :      B  , ,  `�  :  `�  �  a+  �  a+  :  `�  :      B  , ,  ce  :  ce  �  d  �  d  :  ce  :      B  , ,  fI  :  fI  �  f�  �  f�  :  fI  :      B  , ,  i-  :  i-  �  i�  �  i�  :  i-  :      B  , ,  l  :  l  �  l�  �  l�  :  l  :      B  , ,  S  s  S    T)    T)  s  S  s      B  , ,  Vc  s  Vc    W    W  s  Vc  s      B  , ,  YG  s  YG    Y�    Y�  s  YG  s      B  , ,  \+  s  \+    \�    \�  s  \+  s      B  , ,  _  s  _    _�    _�  s  _  s      B  , ,  a�  s  a�    b�    b�  s  a�  s      B  , ,  d�  s  d�    e�    e�  s  d�  s      B  , ,  g�  s  g�    he    he  s  g�  s      B  , ,  j�  s  j�    kI    kI  s  j�  s      B  , ,  nK  A  nK  �  n�  �  n�  A  nK  A      B  , ,  T�  �  T�  8  U�  8  U�  �  T�  �      B  , ,  W�  �  W�  8  X  8  X  �  W�  �      B  , ,  Z�  �  Z�  8  [c  8  [c  �  Z�  �      B  , ,  ]�  �  ]�  8  ^G  8  ^G  �  ]�  �      B  , ,  `�  �  `�  8  a+  8  a+  �  `�  �      B  , ,  ce  �  ce  8  d  8  d  �  ce  �      B  , ,  fI  �  fI  8  f�  8  f�  �  fI  �      B  , ,  i-  �  i-  8  i�  8  i�  �  i-  �      B  , ,  l  �  l  8  l�  8  l�  �  l  �      B  , ,  nK  �  nK  �  n�  �  n�  �  nK  �      B  , ,  T  q  T    T�    T�  q  T  q      B  , ,  UU  q  UU    U�    U�  q  UU  q      B  , ,  V�  q  V�    WS    WS  q  V�  q      B  , ,  W�  q  W�    X�    X�  q  W�  q      B  , ,  YQ  q  YQ    Y�    Y�  q  YQ  q      B  , ,  Z�  q  Z�    [O    [O  q  Z�  q      B  , ,  [�  q  [�    \�    \�  q  [�  q      B  , ,  ]M  q  ]M    ]�    ]�  q  ]M  q      B  , ,  ^�  q  ^�    _K    _K  q  ^�  q      B  , ,  _�  q  _�    `�    `�  q  _�  q      B  , ,  aI  q  aI    a�    a�  q  aI  q      B  , ,  b�  q  b�    cG    cG  q  b�  q      B  , ,  c�  q  c�    d�    d�  q  c�  q      B  , ,  eE  q  eE    e�    e�  q  eE  q      B  , ,  f�  q  f�    gC    gC  q  f�  q      B  , ,  g�  q  g�    h�    h�  q  g�  q      B  , ,  iA  q  iA    i�    i�  q  iA  q      B  , ,  j�  q  j�    k?    k?  q  j�  q      B  , ,  k�  q  k�    l�    l�  q  k�  q      B  , ,  nK  �  nK  C  n�  C  n�  �  nK  �      B  , ,  =�  �  =�  8  >{  8  >{  �  =�  �      B  , ,  @�  �  @�  8  A_  8  A_  �  @�  �      B  , ,  C�  �  C�  8  DC  8  DC  �  C�  �      B  , ,  F}  �  F}  8  G'  8  G'  �  F}  �      B  , ,  Ia  �  Ia  8  J  8  J  �  Ia  �      B  , ,  LE  �  LE  8  L�  8  L�  �  LE  �      B  , ,  O)  �  O)  8  O�  8  O�  �  O)  �      B  , ,  R  �  R  8  R�  8  R�  �  R  �      B  , ,  H  q  H    H�    H�  q  H  q      B  , ,  Ia  q  Ia    J    J  q  Ia  q      B  , ,  J�  q  J�    K_    K_  q  J�  q      B  , ,  L	  q  L	    L�    L�  q  L	  q      B  , ,  M]  q  M]    N    N  q  M]  q      B  , ,  N�  q  N�    O[    O[  q  N�  q      B  , ,  P  q  P    P�    P�  q  P  q      B  , ,  QY  q  QY    R    R  q  QY  q      B  , ,  9q  q  9q    :    :  q  9q  q      B  , ,  9{  s  9{    :%    :%  s  9{  s      B  , ,  <_  s  <_    =	    =	  s  <_  s      B  , ,  ?C  s  ?C    ?�    ?�  s  ?C  s      B  , ,  B'  s  B'    B�    B�  s  B'  s      B  , ,  E  s  E    E�    E�  s  E  s      B  , ,  G�  s  G�    H�    H�  s  G�  s      B  , ,  J�  s  J�    K}    K}  s  J�  s      B  , ,  M�  s  M�    Na    Na  s  M�  s      B  , ,  P�  s  P�    QE    QE  s  P�  s      B  , ,  :�  q  :�    ;o    ;o  q  :�  q      B  , ,  <  q  <    <�    <�  q  <  q      B  , ,  =m  q  =m    >    >  q  =m  q      B  , ,  >�  q  >�    ?k    ?k  q  >�  q      B  , ,  @  q  @    @�    @�  q  @  q      B  , ,  Ai  q  Ai    B    B  q  Ai  q      B  , ,  B�  q  B�    Cg    Cg  q  B�  q      B  , ,  D  q  D    D�    D�  q  D  q      B  , ,  Ee  q  Ee    F    F  q  Ee  q      B  , ,  F�  q  F�    Gc    Gc  q  F�  q      B  , ,  8	  �  8	  8  8�  8  8�  �  8	  �      B  , ,  :�  �  :�  8  ;�  8  ;�  �  :�  �      B  , ,  8  q  8    8�    8�  q  8  q      B  , ,  :�  �  :�  �  ;�  �  ;�  �  :�  �      B  , ,  =�  �  =�  �  >{  �  >{  �  =�  �      B  , ,  @�  �  @�  �  A_  �  A_  �  @�  �      B  , ,  C�  �  C�  �  DC  �  DC  �  C�  �      B  , ,  F}  �  F}  �  G'  �  G'  �  F}  �      B  , ,  Ia  �  Ia  �  J  �  J  �  Ia  �      B  , ,  LE  �  LE  �  L�  �  L�  �  LE  �      B  , ,  O)  �  O)  �  O�  �  O�  �  O)  �      B  , ,  R  �  R  �  R�  �  R�  �  R  �      B  , ,  8	  �  8	  <  8�  <  8�  �  8	  �      B  , ,  :�  �  :�  <  ;�  <  ;�  �  :�  �      B  , ,  =�  �  =�  <  >{  <  >{  �  =�  �      B  , ,  @�  �  @�  <  A_  <  A_  �  @�  �      B  , ,  C�  �  C�  <  DC  <  DC  �  C�  �      B  , ,  F}  �  F}  <  G'  <  G'  �  F}  �      B  , ,  Ia  �  Ia  <  J  <  J  �  Ia  �      B  , ,  LE  �  LE  <  L�  <  L�  �  LE  �      B  , ,  O)  �  O)  <  O�  <  O�  �  O)  �      B  , ,  R  �  R  <  R�  <  R�  �  R  �      B  , ,  8	  >  8	  �  8�  �  8�  >  8	  >      B  , ,  :�  >  :�  �  ;�  �  ;�  >  :�  >      B  , ,  =�  >  =�  �  >{  �  >{  >  =�  >      B  , ,  @�  >  @�  �  A_  �  A_  >  @�  >      B  , ,  C�  >  C�  �  DC  �  DC  >  C�  >      B  , ,  F}  >  F}  �  G'  �  G'  >  F}  >      B  , ,  Ia  >  Ia  �  J  �  J  >  Ia  >      B  , ,  LE  >  LE  �  L�  �  L�  >  LE  >      B  , ,  O)  >  O)  �  O�  �  O�  >  O)  >      B  , ,  R  >  R  �  R�  �  R�  >  R  >      B  , ,  8	  �  8	  �  8�  �  8�  �  8	  �      B  , ,  :�  �  :�  �  ;�  �  ;�  �  :�  �      B  , ,  =�  �  =�  �  >{  �  >{  �  =�  �      B  , ,  @�  �  @�  �  A_  �  A_  �  @�  �      B  , ,  C�  �  C�  �  DC  �  DC  �  C�  �      B  , ,  F}  �  F}  �  G'  �  G'  �  F}  �      B  , ,  Ia  �  Ia  �  J  �  J  �  Ia  �      B  , ,  LE  �  LE  �  L�  �  L�  �  LE  �      B  , ,  O)  �  O)  �  O�  �  O�  �  O)  �      B  , ,  R  �  R  �  R�  �  R�  �  R  �      B  , ,  8	  �  8	  �  8�  �  8�  �  8	  �      B  , ,  W�  �  W�  �  X  �  X  �  W�  �      B  , ,  Z�  �  Z�  �  [c  �  [c  �  Z�  �      B  , ,  ]�  �  ]�  �  ^G  �  ^G  �  ]�  �      B  , ,  `�  �  `�  �  a+  �  a+  �  `�  �      B  , ,  ce  �  ce  �  d  �  d  �  ce  �      B  , ,  fI  �  fI  �  f�  �  f�  �  fI  �      B  , ,  i-  �  i-  �  i�  �  i�  �  i-  �      B  , ,  l  �  l  �  l�  �  l�  �  l  �      B  , ,  nK  E  nK  �  n�  �  n�  E  nK  E      B  , ,  T�  >  T�  �  U�  �  U�  >  T�  >      B  , ,  W�  >  W�  �  X  �  X  >  W�  >      B  , ,  Z�  >  Z�  �  [c  �  [c  >  Z�  >      B  , ,  ]�  >  ]�  �  ^G  �  ^G  >  ]�  >      B  , ,  `�  >  `�  �  a+  �  a+  >  `�  >      B  , ,  ce  >  ce  �  d  �  d  >  ce  >      B  , ,  fI  >  fI  �  f�  �  f�  >  fI  >      B  , ,  i-  >  i-  �  i�  �  i�  >  i-  >      B  , ,  l  >  l  �  l�  �  l�  >  l  >      B  , ,  nK  �  nK  G  n�  G  n�  �  nK  �      B  , ,  T�  �  T�  <  U�  <  U�  �  T�  �      B  , ,  W�  �  W�  <  X  <  X  �  W�  �      B  , ,  Z�  �  Z�  <  [c  <  [c  �  Z�  �      B  , ,  ]�  �  ]�  <  ^G  <  ^G  �  ]�  �      B  , ,  `�  �  `�  <  a+  <  a+  �  `�  �      B  , ,  ce  �  ce  <  d  <  d  �  ce  �      B  , ,  fI  �  fI  <  f�  <  f�  �  fI  �      B  , ,  i-  �  i-  <  i�  <  i�  �  i-  �      B  , ,  l  �  l  <  l�  <  l�  �  l  �      B  , ,  nK  �  nK  �  n�  �  n�  �  nK  �      B  , ,  T�  �  T�  �  U�  �  U�  �  T�  �      B  , ,  W�  �  W�  �  X  �  X  �  W�  �      B  , ,  Z�  �  Z�  �  [c  �  [c  �  Z�  �      B  , ,  ]�  �  ]�  �  ^G  �  ^G  �  ]�  �      B  , ,  `�  �  `�  �  a+  �  a+  �  `�  �      B  , ,  ce  �  ce  �  d  �  d  �  ce  �      B  , ,  fI  �  fI  �  f�  �  f�  �  fI  �      B  , ,  i-  �  i-  �  i�  �  i�  �  i-  �      B  , ,  l  �  l  �  l�  �  l�  �  l  �      B  , ,  nK  I  nK  �  n�  �  n�  I  nK  I      B  , ,  T�  �  T�  �  U�  �  U�  �  T�  �      B  , ,  !  �  !  �  �  �  �  �  !  �      B  , ,  !  �  !  <  �  <  �  �  !  �      B  , ,  !  �  !  8  �  8  �  �  !  �      B  , ,  !  >  !  �  �  �  �  >  !  >      B  , ,    :    �  �  �  �  :    :      B  , ,    :    �  �  �  �  :    :      B  , ,  �  :  �  �  �  �  �  :  �  :      B  , ,  !  �  !  �  �  �  �  �  !  �      B  , ,  	�  :  	�  �  
s  �  
s  :  	�  :      B  , ,  �  :  �  �  W  �  W  :  �  :      B  , ,  �  :  �  �  ;  �  ;  :  �  :      B  , ,  u  :  u  �    �    :  u  :      B  , ,  Y  :  Y  �    �    :  Y  :      B  , ,  =  :  =  �  �  �  �  :  =  :      B  , ,  !  :  !  �  �  �  �  :  !  :      B  , ,    :    �  �  �  �  :    :      B  , ,   �  :   �  �  !�  �  !�  :   �  :      B  , ,  #�  :  #�  �  $w  �  $w  :  #�  :      B  , ,  &�  :  &�  �  '[  �  '[  :  &�  :      B  , ,  )�  :  )�  �  *?  �  *?  :  )�  :      B  , ,  ,y  :  ,y  �  -#  �  -#  :  ,y  :      B  , ,  /]  :  /]  �  0  �  0  :  /]  :      B  , ,  2A  :  2A  �  2�  �  2�  :  2A  :      B  , ,  5%  :  5%  �  5�  �  5�  :  5%  :      B  , ,  2A  �  2A  8  2�  8  2�  �  2A  �      B  , ,  5%  �  5%  8  5�  8  5�  �  5%  �      B  , ,  !�  q  !�    "3    "3  q  !�  q      B  , ,  "�  q  "�    #�    #�  q  "�  q      B  , ,  $1  q  $1    $�    $�  q  $1  q      B  , ,  %?  s  %?    %�    %�  s  %?  s      B  , ,  %�  q  %�    &/    &/  q  %�  q      B  , ,  &�  q  &�    '�    '�  q  &�  q      B  , ,  (-  q  (-    (�    (�  q  (-  q      B  , ,  )�  q  )�    *+    *+  q  )�  q      B  , ,  *�  q  *�    +    +  q  *�  q      B  , ,  ,)  q  ,)    ,�    ,�  q  ,)  q      B  , ,  -}  q  -}    .'    .'  q  -}  q      B  , ,  .�  q  .�    /{    /{  q  .�  q      B  , ,  0%  q  0%    0�    0�  q  0%  q      B  , ,  1y  q  1y    2#    2#  q  1y  q      B  , ,  2�  q  2�    3w    3w  q  2�  q      B  , ,  4!  q  4!    4�    4�  q  4!  q      B  , ,  5u  q  5u    6    6  q  5u  q      B  , ,  6�  q  6�    7s    7s  q  6�  q      B  , ,  (#  s  (#    (�    (�  s  (#  s      B  , ,  +  s  +    +�    +�  s  +  s      B  , ,  -�  s  -�    .�    .�  s  -�  s      B  , ,  0�  s  0�    1y    1y  s  0�  s      B  , ,  3�  s  3�    4]    4]  s  3�  s      B  , ,  6�  s  6�    7A    7A  s  6�  s      B  , ,  �  s  �    =    =  s  �  s      B  , ,  9  q  9    �    �  q  9  q      B  , ,  �  q  �    7    7  q  �  q      B  , ,  �  q  �    �    �  q  �  q      B  , ,   5  q   5     �     �  q   5  q      B  , ,  w  s  w     !     !  s  w  s      B  , ,  "[  s  "[    #    #  s  "[  s      B  , ,    �    8  �  8  �  �    �      B  , ,   �  �   �  8  !�  8  !�  �   �  �      B  , ,  #�  �  #�  8  $w  8  $w  �  #�  �      B  , ,  &�  �  &�  8  '[  8  '[  �  &�  �      B  , ,  )�  �  )�  8  *?  8  *?  �  )�  �      B  , ,  ,y  �  ,y  8  -#  8  -#  �  ,y  �      B  , ,  /]  �  /]  8  0  8  0  �  /]  �      B  , ,  �  s  �    u    u  s  �  s      B  , ,  �  �  �  8  �  8  �  �  �  �      B  , ,  	�  �  	�  8  
s  8  
s  �  	�  �      B  , ,  �  �  �  8  W  8  W  �  �  �      B  , ,  �  �  �  8  ;  8  ;  �  �  �      B  , ,  u  �  u  8    8    �  u  �      B  , ,  Y  �  Y  8    8    �  Y  �      B  , ,  =  �  =  8  �  8  �  �  =  �      B  , ,  �  q  �    O    O  q  �  q      B  , ,  �  q  �    �    �  q  �  q      B  , ,   U  q   U     �     �  q   U  q      B  , ,  	�  q  	�    
K    
K  q  	�  q      B  , ,  
�  q  
�    �    �  q  
�  q      B  , ,  I  q  I    �    �  q  I  q      B  , ,  �  q  �    G    G  q  �  q      B  , ,  �  q  �    �    �  q  �  q      B  , ,  E  q  E    �    �  q  E  q      B  , ,  �  q  �    C    C  q  �  q      B  , ,  �  q  �    �    �  q  �  q      B  , ,  A  q  A    �    �  q  A  q      B  , ,  �  q  �    ?    ?  q  �  q      B  , ,  �  q  �    �    �  q  �  q      B  , ,  =  q  =    �    �  q  =  q      B  , ,  �  q  �    ;    ;  q  �  q      B  , ,  �  q  �    �    �  q  �  q      B  , ,  �  s  �    Y    Y  s  �  s      B  , ,    s      �    �  s    s      B  , ,  �  s  �    �    �  s  �  s      B  , ,  M  q  M    �    �  q  M  q      B  , ,    �    8  �  8  �  �    �      B  , ,    �    8  �  8  �  �    �      B  , ,  �  s  �    9    9  s  �  s      B  , ,  s  s  s          s  s  s      B  , ,  W  s  W    	    	  s  W  s      B  , ,  ;  s  ;    �    �  s  ;  s      B  , ,    s      �    �  s    s      B  , ,  �  q  �    S    S  q  �  q      B  , ,  �  q  �    �    �  q  �  q      B  , ,  Q  q  Q    �    �  q  Q  q      B  , ,    >    �  �  �  �  >    >      B  , ,  �  >  �  �  �  �  �  >  �  >      B  , ,    �    �  �  �  �  �    �      B  , ,    �    �  �  �  �  �    �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  	�  �  	�  �  
s  �  
s  �  	�  �      B  , ,  �  �  �  �  W  �  W  �  �  �      B  , ,  �  �  �  �  ;  �  ;  �  �  �      B  , ,  u  �  u  �    �    �  u  �      B  , ,  Y  �  Y  �    �    �  Y  �      B  , ,  =  �  =  �  �  �  �  �  =  �      B  , ,  	�  >  	�  �  
s  �  
s  >  	�  >      B  , ,  �  >  �  �  W  �  W  >  �  >      B  , ,  �  >  �  �  ;  �  ;  >  �  >      B  , ,  u  >  u  �    �    >  u  >      B  , ,  Y  >  Y  �    �    >  Y  >      B  , ,  =  >  =  �  �  �  �  >  =  >      B  , ,  u  �  u  �    �    �  u  �      B  , ,  Y  �  Y  �    �    �  Y  �      B  , ,  =  �  =  �  �  �  �  �  =  �      B  , ,    �    �  �  �  �  �    �      B  , ,    �    �  �  �  �  �    �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,    �    <  �  <  �  �    �      B  , ,    �    <  �  <  �  �    �      B  , ,  �  �  �  <  �  <  �  �  �  �      B  , ,  	�  �  	�  <  
s  <  
s  �  	�  �      B  , ,  �  �  �  <  W  <  W  �  �  �      B  , ,  �  �  �  <  ;  <  ;  �  �  �      B  , ,  u  �  u  <    <    �  u  �      B  , ,  Y  �  Y  <    <    �  Y  �      B  , ,  =  �  =  <  �  <  �  �  =  �      B  , ,  	�  �  	�  �  
s  �  
s  �  	�  �      B  , ,  �  �  �  �  W  �  W  �  �  �      B  , ,  �  �  �  �  ;  �  ;  �  �  �      B  , ,    >    �  �  �  �  >    >      B  , ,  &�  �  &�  <  '[  <  '[  �  &�  �      B  , ,  )�  �  )�  <  *?  <  *?  �  )�  �      B  , ,  ,y  �  ,y  <  -#  <  -#  �  ,y  �      B  , ,    �    �  �  �  �  �    �      B  , ,   �  �   �  �  !�  �  !�  �   �  �      B  , ,  #�  �  #�  �  $w  �  $w  �  #�  �      B  , ,  &�  �  &�  �  '[  �  '[  �  &�  �      B  , ,  )�  �  )�  �  *?  �  *?  �  )�  �      B  , ,  ,y  �  ,y  �  -#  �  -#  �  ,y  �      B  , ,  /]  �  /]  �  0  �  0  �  /]  �      B  , ,  2A  �  2A  �  2�  �  2�  �  2A  �      B  , ,  5%  �  5%  �  5�  �  5�  �  5%  �      B  , ,  /]  �  /]  <  0  <  0  �  /]  �      B  , ,  2A  �  2A  <  2�  <  2�  �  2A  �      B  , ,  5%  �  5%  <  5�  <  5�  �  5%  �      B  , ,  &�  �  &�  �  '[  �  '[  �  &�  �      B  , ,  )�  �  )�  �  *?  �  *?  �  )�  �      B  , ,  ,y  �  ,y  �  -#  �  -#  �  ,y  �      B  , ,  /]  �  /]  �  0  �  0  �  /]  �      B  , ,  2A  �  2A  �  2�  �  2�  �  2A  �      B  , ,  5%  �  5%  �  5�  �  5�  �  5%  �      B  , ,    �    �  �  �  �  �    �      B  , ,   �  �   �  �  !�  �  !�  �   �  �      B  , ,  #�  �  #�  �  $w  �  $w  �  #�  �      B  , ,    �    <  �  <  �  �    �      B  , ,   �  �   �  <  !�  <  !�  �   �  �      B  , ,  #�  �  #�  <  $w  <  $w  �  #�  �      B  , ,    >    �  �  �  �  >    >      B  , ,   �  >   �  �  !�  �  !�  >   �  >      B  , ,  #�  >  #�  �  $w  �  $w  >  #�  >      B  , ,  &�  >  &�  �  '[  �  '[  >  &�  >      B  , ,  )�  >  )�  �  *?  �  *?  >  )�  >      B  , ,  ,y  >  ,y  �  -#  �  -#  >  ,y  >      B  , ,  /]  >  /]  �  0  �  0  >  /]  >      B  , ,  2A  >  2A  �  2�  �  2�  >  2A  >      B  , ,  5%  >  5%  �  5�  �  5�  >  5%  >      B  , ,  !  
�  !  @  �  @  �  
�  !  
�      B  , ,  !  	B  !  	�  �  	�  �  	B  !  	B      B  , ,  !  �  !  �  �  �  �  �  !  �      B  , ,  !  �  !  D  �  D  �  �  !  �      B  , ,    F    �  �  �  �  F    F      B  , ,    F    �  �  �  �  F    F      B  , ,  �  F  �  �  �  �  �  F  �  F      B  , ,  	�  F  	�  �  
s  �  
s  F  	�  F      B  , ,  �  F  �  �  W  �  W  F  �  F      B  , ,  �  F  �  �  ;  �  ;  F  �  F      B  , ,  u  F  u  �    �    F  u  F      B  , ,  Y  F  Y  �    �    F  Y  F      B  , ,  =  F  =  �  �  �  �  F  =  F      B  , ,  !  F  !  �  �  �  �  F  !  F      B  , ,    F    �  �  �  �  F    F      B  , ,   �  F   �  �  !�  �  !�  F   �  F      B  , ,  #�  F  #�  �  $w  �  $w  F  #�  F      B  , ,  &�  F  &�  �  '[  �  '[  F  &�  F      B  , ,  )�  F  )�  �  *?  �  *?  F  )�  F      B  , ,  ,y  F  ,y  �  -#  �  -#  F  ,y  F      B  , ,  /]  F  /]  �  0  �  0  F  /]  F      B  , ,  2A  F  2A  �  2�  �  2�  F  2A  F      B  , ,  5%  F  5%  �  5�  �  5�  F  5%  F      B  , ,  !  �  !  �  �  �  �  �  !  �      B  , ,  !  �  !  H  �  H  �  �  !  �      B  , ,  )�  �  )�  �  *?  �  *?  �  )�  �      B  , ,  ,y  �  ,y  �  -#  �  -#  �  ,y  �      B  , ,  /]  �  /]  �  0  �  0  �  /]  �      B  , ,  2A  �  2A  �  2�  �  2�  �  2A  �      B  , ,  5%  �  5%  �  5�  �  5�  �  5%  �      B  , ,  #�  
�  #�  @  $w  @  $w  
�  #�  
�      B  , ,    �    D  �  D  �  �    �      B  , ,   �  �   �  D  !�  D  !�  �   �  �      B  , ,  #�  �  #�  D  $w  D  $w  �  #�  �      B  , ,  &�  �  &�  D  '[  D  '[  �  &�  �      B  , ,  )�  �  )�  D  *?  D  *?  �  )�  �      B  , ,  ,y  �  ,y  D  -#  D  -#  �  ,y  �      B  , ,  /]  �  /]  D  0  D  0  �  /]  �      B  , ,  2A  �  2A  D  2�  D  2�  �  2A  �      B  , ,  5%  �  5%  D  5�  D  5�  �  5%  �      B  , ,  &�  
�  &�  @  '[  @  '[  
�  &�  
�      B  , ,  )�  
�  )�  @  *?  @  *?  
�  )�  
�      B  , ,  ,y  
�  ,y  @  -#  @  -#  
�  ,y  
�      B  , ,  /]  
�  /]  @  0  @  0  
�  /]  
�      B  , ,  2A  
�  2A  @  2�  @  2�  
�  2A  
�      B  , ,  5%  
�  5%  @  5�  @  5�  
�  5%  
�      B  , ,    
�    @  �  @  �  
�    
�      B  , ,    	B    	�  �  	�  �  	B    	B      B  , ,   �  	B   �  	�  !�  	�  !�  	B   �  	B      B  , ,  #�  	B  #�  	�  $w  	�  $w  	B  #�  	B      B  , ,  &�  	B  &�  	�  '[  	�  '[  	B  &�  	B      B  , ,  )�  	B  )�  	�  *?  	�  *?  	B  )�  	B      B  , ,  ,y  	B  ,y  	�  -#  	�  -#  	B  ,y  	B      B  , ,  /]  	B  /]  	�  0  	�  0  	B  /]  	B      B  , ,  2A  	B  2A  	�  2�  	�  2�  	B  2A  	B      B  , ,  5%  	B  5%  	�  5�  	�  5�  	B  5%  	B      B  , ,   �  
�   �  @  !�  @  !�  
�   �  
�      B  , ,    �    �  �  �  �  �    �      B  , ,   �  �   �  �  !�  �  !�  �   �  �      B  , ,  #�  �  #�  �  $w  �  $w  �  #�  �      B  , ,  &�  �  &�  �  '[  �  '[  �  &�  �      B  , ,  Y  �  Y  D    D    �  Y  �      B  , ,  =  �  =  D  �  D  �  �  =  �      B  , ,    
�    @  �  @  �  
�    
�      B  , ,    	B    	�  �  	�  �  	B    	B      B  , ,    	B    	�  �  	�  �  	B    	B      B  , ,  �  	B  �  	�  �  	�  �  	B  �  	B      B  , ,  	�  	B  	�  	�  
s  	�  
s  	B  	�  	B      B  , ,    �    �  �  �  �  �    �      B  , ,    �    �  �  �  �  �    �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  	�  �  	�  �  
s  �  
s  �  	�  �      B  , ,  �  �  �  �  W  �  W  �  �  �      B  , ,  �  �  �  �  ;  �  ;  �  �  �      B  , ,  u  �  u  �    �    �  u  �      B  , ,  Y  �  Y  �    �    �  Y  �      B  , ,  =  �  =  �  �  �  �  �  =  �      B  , ,  �  	B  �  	�  W  	�  W  	B  �  	B      B  , ,  �  	B  �  	�  ;  	�  ;  	B  �  	B      B  , ,  u  	B  u  	�    	�    	B  u  	B      B  , ,  Y  	B  Y  	�    	�    	B  Y  	B      B  , ,  =  	B  =  	�  �  	�  �  	B  =  	B      B  , ,  �  
�  �  @  W  @  W  
�  �  
�      B  , ,  �  
�  �  @  ;  @  ;  
�  �  
�      B  , ,  u  
�  u  @    @    
�  u  
�      B  , ,  Y  
�  Y  @    @    
�  Y  
�      B  , ,  =  
�  =  @  �  @  �  
�  =  
�      B  , ,    �    D  �  D  �  �    �      B  , ,    �    D  �  D  �  �    �      B  , ,  �  �  �  D  �  D  �  �  �  �      B  , ,  	�  �  	�  D  
s  D  
s  �  	�  �      B  , ,  �  �  �  D  W  D  W  �  �  �      B  , ,  �  �  �  D  ;  D  ;  �  �  �      B  , ,  u  �  u  D    D    �  u  �      B  , ,    
�    @  �  @  �  
�    
�      B  , ,  �  
�  �  @  �  @  �  
�  �  
�      B  , ,  	�  
�  	�  @  
s  @  
s  
�  	�  
�      B  , ,  �  �  �  �  ;  �  ;  �  �  �      B  , ,  u  �  u  �    �    �  u  �      B  , ,  Y  �  Y  �    �    �  Y  �      B  , ,  =  �  =  �  �  �  �  �  =  �      B  , ,    �    �  �  �  �  �    �      B  , ,    �    H  �  H  �  �    �      B  , ,    �    H  �  H  �  �    �      B  , ,  �  �  �  H  �  H  �  �  �  �      B  , ,  	�  �  	�  H  
s  H  
s  �  	�  �      B  , ,  �  �  �  H  W  H  W  �  �  �      B  , ,  �  �  �  H  ;  H  ;  �  �  �      B  , ,  u  �  u  H    H    �  u  �      B  , ,  Y  �  Y  H    H    �  Y  �      B  , ,  =  �  =  H  �  H  �  �  =  �      B  , ,    �    �  �  �  �  �    �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �   �  �  c  9  c  9   �  �   �      B  , ,  s   �  s  c    c     �  s   �      B  , ,  W   �  W  c  	  c  	   �  W   �      B  , ,  ;   �  ;  c  �  c  �   �  ;   �      B  , ,     �    c  �  c  �   �     �      B  , ,     �    c  �  c  �   �     �      B  , ,  �   �  �  c  �  c  �   �  �   �      B  , ,  �   �  �  c  u  c  u   �  �   �      B  , ,  �   �  �  c  Y  c  Y   �  �   �      B  , ,  	�  �  	�  �  
s  �  
s  �  	�  �      B  , ,  �  �  �  �  W  �  W  �  �  �      B  , ,  &�  �  &�  H  '[  H  '[  �  &�  �      B  , ,  )�  �  )�  H  *?  H  *?  �  )�  �      B  , ,  ,y  �  ,y  H  -#  H  -#  �  ,y  �      B  , ,  /]  �  /]  H  0  H  0  �  /]  �      B  , ,  2A  �  2A  H  2�  H  2�  �  2A  �      B  , ,  5%  �  5%  H  5�  H  5�  �  5%  �      B  , ,   �  �   �  �  !�  �  !�  �   �  �      B  , ,  #�  �  #�  �  $w  �  $w  �  #�  �      B  , ,  &�  �  &�  �  '[  �  '[  �  &�  �      B  , ,  )�  �  )�  �  *?  �  *?  �  )�  �      B  , ,  ,y  �  ,y  �  -#  �  -#  �  ,y  �      B  , ,  /]  �  /]  �  0  �  0  �  /]  �      B  , ,  2A  �  2A  �  2�  �  2�  �  2A  �      B  , ,  5%  �  5%  �  5�  �  5�  �  5%  �      B  , ,    �    �  �  �  �  �    �      B  , ,    �    H  �  H  �  �    �      B  , ,  �   �  �  c  =  c  =   �  �   �      B  , ,  w   �  w  c   !  c   !   �  w   �      B  , ,  "[   �  "[  c  #  c  #   �  "[   �      B  , ,  %?   �  %?  c  %�  c  %�   �  %?   �      B  , ,  (#   �  (#  c  (�  c  (�   �  (#   �      B  , ,  +   �  +  c  +�  c  +�   �  +   �      B  , ,  -�   �  -�  c  .�  c  .�   �  -�   �      B  , ,  0�   �  0�  c  1y  c  1y   �  0�   �      B  , ,  3�   �  3�  c  4]  c  4]   �  3�   �      B  , ,  6�   �  6�  c  7A  c  7A   �  6�   �      B  , ,   �  �   �  H  !�  H  !�  �   �  �      B  , ,  #�  �  #�  H  $w  H  $w  �  #�  �      B  , ,  8	  F  8	  �  8�  �  8�  F  8	  F      B  , ,  :�  F  :�  �  ;�  �  ;�  F  :�  F      B  , ,  =�  F  =�  �  >{  �  >{  F  =�  F      B  , ,  @�  F  @�  �  A_  �  A_  F  @�  F      B  , ,  C�  F  C�  �  DC  �  DC  F  C�  F      B  , ,  F}  F  F}  �  G'  �  G'  F  F}  F      B  , ,  Ia  F  Ia  �  J  �  J  F  Ia  F      B  , ,  LE  F  LE  �  L�  �  L�  F  LE  F      B  , ,  O)  F  O)  �  O�  �  O�  F  O)  F      B  , ,  R  F  R  �  R�  �  R�  F  R  F      B  , ,  T�  F  T�  �  U�  �  U�  F  T�  F      B  , ,  W�  F  W�  �  X  �  X  F  W�  F      B  , ,  Z�  F  Z�  �  [c  �  [c  F  Z�  F      B  , ,  ]�  F  ]�  �  ^G  �  ^G  F  ]�  F      B  , ,  `�  F  `�  �  a+  �  a+  F  `�  F      B  , ,  ce  F  ce  �  d  �  d  F  ce  F      B  , ,  fI  F  fI  �  f�  �  f�  F  fI  F      B  , ,  i-  F  i-  �  i�  �  i�  F  i-  F      B  , ,  l  F  l  �  l�  �  l�  F  l  F      B  , ,  nK  �  nK  O  n�  O  n�  �  nK  �      B  , ,  nK  	�  nK  
K  n�  
K  n�  	�  nK  	�      B  , ,  T�  
�  T�  @  U�  @  U�  
�  T�  
�      B  , ,  W�  
�  W�  @  X  @  X  
�  W�  
�      B  , ,  Z�  
�  Z�  @  [c  @  [c  
�  Z�  
�      B  , ,  ]�  
�  ]�  @  ^G  @  ^G  
�  ]�  
�      B  , ,  `�  
�  `�  @  a+  @  a+  
�  `�  
�      B  , ,  ce  
�  ce  @  d  @  d  
�  ce  
�      B  , ,  fI  
�  fI  @  f�  @  f�  
�  fI  
�      B  , ,  i-  
�  i-  @  i�  @  i�  
�  i-  
�      B  , ,  l  
�  l  @  l�  @  l�  
�  l  
�      B  , ,  T�  �  T�  �  U�  �  U�  �  T�  �      B  , ,  W�  �  W�  �  X  �  X  �  W�  �      B  , ,  Z�  �  Z�  �  [c  �  [c  �  Z�  �      B  , ,  ]�  �  ]�  �  ^G  �  ^G  �  ]�  �      B  , ,  `�  �  `�  �  a+  �  a+  �  `�  �      B  , ,  ce  �  ce  �  d  �  d  �  ce  �      B  , ,  fI  �  fI  �  f�  �  f�  �  fI  �      B  , ,  i-  �  i-  �  i�  �  i�  �  i-  �      B  , ,  l  �  l  �  l�  �  l�  �  l  �      B  , ,  nK  M  nK  �  n�  �  n�  M  nK  M      B  , ,  T�  	B  T�  	�  U�  	�  U�  	B  T�  	B      B  , ,  W�  	B  W�  	�  X  	�  X  	B  W�  	B      B  , ,  Z�  	B  Z�  	�  [c  	�  [c  	B  Z�  	B      B  , ,  ]�  	B  ]�  	�  ^G  	�  ^G  	B  ]�  	B      B  , ,  `�  	B  `�  	�  a+  	�  a+  	B  `�  	B      B  , ,  ce  	B  ce  	�  d  	�  d  	B  ce  	B      B  , ,  fI  	B  fI  	�  f�  	�  f�  	B  fI  	B      B  , ,  i-  	B  i-  	�  i�  	�  i�  	B  i-  	B      B  , ,  l  	B  l  	�  l�  	�  l�  	B  l  	B      B  , ,  T�  �  T�  D  U�  D  U�  �  T�  �      B  , ,  W�  �  W�  D  X  D  X  �  W�  �      B  , ,  Z�  �  Z�  D  [c  D  [c  �  Z�  �      B  , ,  ]�  �  ]�  D  ^G  D  ^G  �  ]�  �      B  , ,  `�  �  `�  D  a+  D  a+  �  `�  �      B  , ,  ce  �  ce  D  d  D  d  �  ce  �      B  , ,  fI  �  fI  D  f�  D  f�  �  fI  �      B  , ,  i-  �  i-  D  i�  D  i�  �  i-  �      B  , ,  l  �  l  D  l�  D  l�  �  l  �      B  , ,  nK  �  nK  �  n�  �  n�  �  nK  �      B  , ,  8	  
�  8	  @  8�  @  8�  
�  8	  
�      B  , ,  8	  	B  8	  	�  8�  	�  8�  	B  8	  	B      B  , ,  :�  	B  :�  	�  ;�  	�  ;�  	B  :�  	B      B  , ,  =�  	B  =�  	�  >{  	�  >{  	B  =�  	B      B  , ,  @�  	B  @�  	�  A_  	�  A_  	B  @�  	B      B  , ,  C�  	B  C�  	�  DC  	�  DC  	B  C�  	B      B  , ,  F}  	B  F}  	�  G'  	�  G'  	B  F}  	B      B  , ,  Ia  	B  Ia  	�  J  	�  J  	B  Ia  	B      B  , ,  LE  	B  LE  	�  L�  	�  L�  	B  LE  	B      B  , ,  O)  	B  O)  	�  O�  	�  O�  	B  O)  	B      B  , ,  R  	B  R  	�  R�  	�  R�  	B  R  	B      B  , ,  8	  �  8	  �  8�  �  8�  �  8	  �      B  , ,  :�  �  :�  �  ;�  �  ;�  �  :�  �      B  , ,  =�  �  =�  �  >{  �  >{  �  =�  �      B  , ,  @�  �  @�  �  A_  �  A_  �  @�  �      B  , ,  C�  �  C�  �  DC  �  DC  �  C�  �      B  , ,  F}  �  F}  �  G'  �  G'  �  F}  �      B  , ,  Ia  �  Ia  �  J  �  J  �  Ia  �      B  , ,  LE  �  LE  �  L�  �  L�  �  LE  �      B  , ,  O)  �  O)  �  O�  �  O�  �  O)  �      B  , ,  8	  �  8	  D  8�  D  8�  �  8	  �      B  , ,  :�  �  :�  D  ;�  D  ;�  �  :�  �      B  , ,  =�  �  =�  D  >{  D  >{  �  =�  �      B  , ,  @�  �  @�  D  A_  D  A_  �  @�  �      B  , ,  C�  �  C�  D  DC  D  DC  �  C�  �      B  , ,  F}  �  F}  D  G'  D  G'  �  F}  �      B  , ,  Ia  �  Ia  D  J  D  J  �  Ia  �      B  , ,  LE  �  LE  D  L�  D  L�  �  LE  �      B  , ,  O)  �  O)  D  O�  D  O�  �  O)  �      B  , ,  R  �  R  D  R�  D  R�  �  R  �      B  , ,  R  �  R  �  R�  �  R�  �  R  �      B  , ,  @�  
�  @�  @  A_  @  A_  
�  @�  
�      B  , ,  C�  
�  C�  @  DC  @  DC  
�  C�  
�      B  , ,  F}  
�  F}  @  G'  @  G'  
�  F}  
�      B  , ,  Ia  
�  Ia  @  J  @  J  
�  Ia  
�      B  , ,  LE  
�  LE  @  L�  @  L�  
�  LE  
�      B  , ,  O)  
�  O)  @  O�  @  O�  
�  O)  
�      B  , ,  R  
�  R  @  R�  @  R�  
�  R  
�      B  , ,  :�  
�  :�  @  ;�  @  ;�  
�  :�  
�      B  , ,  =�  
�  =�  @  >{  @  >{  
�  =�  
�      B  , ,  :�  �  :�  �  ;�  �  ;�  �  :�  �      B  , ,  =�  �  =�  �  >{  �  >{  �  =�  �      B  , ,  @�  �  @�  �  A_  �  A_  �  @�  �      B  , ,  C�  �  C�  �  DC  �  DC  �  C�  �      B  , ,  F}  �  F}  �  G'  �  G'  �  F}  �      B  , ,  Ia  �  Ia  �  J  �  J  �  Ia  �      B  , ,  LE  �  LE  �  L�  �  L�  �  LE  �      B  , ,  O)  �  O)  �  O�  �  O�  �  O)  �      B  , ,  8	  �  8	  H  8�  H  8�  �  8	  �      B  , ,  :�  �  :�  H  ;�  H  ;�  �  :�  �      B  , ,  =�  �  =�  H  >{  H  >{  �  =�  �      B  , ,  @�  �  @�  H  A_  H  A_  �  @�  �      B  , ,  C�  �  C�  H  DC  H  DC  �  C�  �      B  , ,  F}  �  F}  H  G'  H  G'  �  F}  �      B  , ,  Ia  �  Ia  H  J  H  J  �  Ia  �      B  , ,  LE  �  LE  H  L�  H  L�  �  LE  �      B  , ,  O)  �  O)  H  O�  H  O�  �  O)  �      B  , ,  R  �  R  H  R�  H  R�  �  R  �      B  , ,  9{   �  9{  c  :%  c  :%   �  9{   �      B  , ,  <_   �  <_  c  =	  c  =	   �  <_   �      B  , ,  ?C   �  ?C  c  ?�  c  ?�   �  ?C   �      B  , ,  B'   �  B'  c  B�  c  B�   �  B'   �      B  , ,  E   �  E  c  E�  c  E�   �  E   �      B  , ,  G�   �  G�  c  H�  c  H�   �  G�   �      B  , ,  J�   �  J�  c  K}  c  K}   �  J�   �      B  , ,  M�   �  M�  c  Na  c  Na   �  M�   �      B  , ,  P�   �  P�  c  QE  c  QE   �  P�   �      B  , ,  R  �  R  �  R�  �  R�  �  R  �      B  , ,  8	  �  8	  �  8�  �  8�  �  8	  �      B  , ,  T�  �  T�  H  U�  H  U�  �  T�  �      B  , ,  W�  �  W�  H  X  H  X  �  W�  �      B  , ,  Z�  �  Z�  H  [c  H  [c  �  Z�  �      B  , ,  ]�  �  ]�  H  ^G  H  ^G  �  ]�  �      B  , ,  `�  �  `�  H  a+  H  a+  �  `�  �      B  , ,  ce  �  ce  H  d  H  d  �  ce  �      B  , ,  fI  �  fI  H  f�  H  f�  �  fI  �      B  , ,  i-  �  i-  H  i�  H  i�  �  i-  �      B  , ,  l  �  l  H  l�  H  l�  �  l  �      B  , ,  nK  �  nK  �  n�  �  n�  �  nK  �      B  , ,  nK  �  nK  S  n�  S  n�  �  nK  �      B  , ,  nK  Q  nK  �  n�  �  n�  Q  nK  Q      B  , ,  T�  �  T�  �  U�  �  U�  �  T�  �      B  , ,  W�  �  W�  �  X  �  X  �  W�  �      B  , ,  Z�  �  Z�  �  [c  �  [c  �  Z�  �      B  , ,  ]�  �  ]�  �  ^G  �  ^G  �  ]�  �      B  , ,  `�  �  `�  �  a+  �  a+  �  `�  �      B  , ,  ce  �  ce  �  d  �  d  �  ce  �      B  , ,  fI  �  fI  �  f�  �  f�  �  fI  �      B  , ,  S   �  S  c  T)  c  T)   �  S   �      B  , ,  Vc   �  Vc  c  W  c  W   �  Vc   �      B  , ,  YG   �  YG  c  Y�  c  Y�   �  YG   �      B  , ,  \+   �  \+  c  \�  c  \�   �  \+   �      B  , ,  _   �  _  c  _�  c  _�   �  _   �      B  , ,  a�   �  a�  c  b�  c  b�   �  a�   �      B  , ,  d�   �  d�  c  e�  c  e�   �  d�   �      B  , ,  g�   �  g�  c  he  c  he   �  g�   �      B  , ,  j�   �  j�  c  kI  c  kI   �  j�   �      B  , ,  nK   U  nK   �  n�   �  n�   U  nK   U      B  , ,  i-  �  i-  �  i�  �  i�  �  i-  �      B  , ,  l  �  l  �  l�  �  l�  �  l  �      B  , ,���  
����  �����  �����  
����  
�      B  , ,���1  :���1  �����  �����  :���1  :      B  , ,���  :���  ���Ϳ  ���Ϳ  :���  :      B  , ,����  :����  ���У  ���У  :����  :      B  , ,����  :����  ���Ӈ  ���Ӈ  :����  :      B  , ,����  :����  ����k  ����k  :����  :      B  , ,��إ  :��إ  ����O  ����O  :��إ  :      B  , ,��ۉ  :��ۉ  ����3  ����3  :��ۉ  :      B  , ,���m  :���m  ����  ����  :���m  :      B  , ,���Q  :���Q  �����  �����  :���Q  :      B  , ,���5  :���5  �����  �����  :���5  :      B  , ,���  :���  �����  �����  :���  :      B  , ,����  :����  ����  ����  :����  :      B  , ,����  :����  ����  ����  :����  :      B  , ,����  :����  ����o  ����o  :����  :      B  , ,���  :���  ����S  ����S  :���  :      B  , ,����  :����  ����7  ����7  :����  :      B  , ,���q  :���q  ����  ����  :���q  :      B  , ,���U  :���U  �����  �����  :���U  :      B  , ,���9  :���9  �����  �����  :���9  :      B  , ,���5  ����5  �����  �����  ����5  �      B  , ,���5  ����5  <����  <����  ����5  �      B  , ,���5  ����5  8����  8����  ����5  �      B  , ,���5  >���5  �����  �����  >���5  >      B  , ,���5  ����5  �����  �����  ����5  �      B  , ,����  q����  ���W  ���W  q����  q      B  , ,���  q���  ����  ����  q���  q      B  , ,���  s���  ���Q  ���Q  s���  s      B  , ,���  s���  ���5  ���5  s���  s      B  , ,���o  s���o  ���  ���  s���o  s      B  , ,���S  s���S  ����  ����  s���S  s      B  , ,���7  s���7  ����  ����  s���7  s      B  , ,���  s���  ����  ����  s���  s      B  , ,���]  q���]  ���  ���  q���]  q      B  , ,����  s����  ����  ����  s����  s      B  , ,����  s����  ����  ����  s����  s      B  , ,����  s����  ���q  ���q  s����  s      B  , ,����  q����  ���[  ���[  q����  q      B  , ,���	  q���	  ����  ����  q���	  q      B  , ,���  ����  8����  8����  ����  �      B  , ,����  �����  8���  8���  �����  �      B  , ,����  �����  8���  8���  �����  �      B  , ,����  �����  8���o  8���o  �����  �      B  , ,���  ����  8���S  8���S  ����  �      B  , ,����  �����  8���7  8���7  �����  �      B  , ,���  q���  ����  ����  q���  q      B  , ,���q  ����q  8���  8���  ����q  �      B  , ,���U  ����U  8����  8����  ����U  �      B  , ,���9  ����9  8����  8����  ����9  �      B  , ,���q  q���q  ���  ���  q���q  q      B  , ,����  q����  ���o  ���o  q����  q      B  , ,���  q���  ����  ����  q���  q      B  , ,���m  q���m  ���  ���  q���m  q      B  , ,����  q����  ���k  ���k  q����  q      B  , ,���  q���  ���  ���  q���  q      B  , ,���i  q���i  ���  ���  q���i  q      B  , ,���  q���  ���g  ���g  q���  q      B  , ,���  q���  ���  ���  q���  q      B  , ,���e  q���e  ���  ���  q���e  q      B  , ,���  q���  ���c  ���c  q���  q      B  , ,���  q���  ���  ���  q���  q      B  , ,���a  q���a  ���  ���  q���a  q      B  , ,����  q����  ���_  ���_  q����  q      B  , ,���Y  q���Y  ���  ���  q���Y  q      B  , ,����  s����  ����  ����  s����  s      B  , ,����  s����  ���m  ���m  s����  s      B  , ,��ȿ  s��ȿ  ���i  ���i  s��ȿ  s      B  , ,���1  ����1  8����  8����  ����1  �      B  , ,��ȍ  q��ȍ  ���7  ���7  q��ȍ  q      B  , ,����  q����  ��ʋ  ��ʋ  q����  q      B  , ,���5  q���5  ����  ����  q���5  q      B  , ,��̉  q��̉  ���3  ���3  q��̉  q      B  , ,����  q����  ��·  ��·  q����  q      B  , ,���1  q���1  ����  ����  q���1  q      B  , ,��Ѕ  q��Ѕ  ���/  ���/  q��Ѕ  q      B  , ,����  q����  ��҃  ��҃  q����  q      B  , ,���-  q���-  ����  ����  q���-  q      B  , ,��ԁ  q��ԁ  ���+  ���+  q��ԁ  q      B  , ,����  q����  ���  ���  q����  q      B  , ,���)  q���)  ����  ����  q���)  q      B  , ,���}  q���}  ���'  ���'  q���}  q      B  , ,����  q����  ���{  ���{  q����  q      B  , ,���%  q���%  ����  ����  q���%  q      B  , ,���y  q���y  ���#  ���#  q���y  q      B  , ,����  q����  ���w  ���w  q����  q      B  , ,���!  q���!  ����  ����  q���!  q      B  , ,���u  q���u  ���  ���  q���u  q      B  , ,����  q����  ���s  ���s  q����  q      B  , ,���  q���  ����  ����  q���  q      B  , ,���  ����  8��Ϳ  8��Ϳ  ����  �      B  , ,����  �����  8��У  8��У  �����  �      B  , ,����  �����  8��Ӈ  8��Ӈ  �����  �      B  , ,����  �����  8���k  8���k  �����  �      B  , ,��إ  ���إ  8���O  8���O  ���إ  �      B  , ,��ۉ  ���ۉ  8���3  8���3  ���ۉ  �      B  , ,���m  ����m  8���  8���  ����m  �      B  , ,���Q  ����Q  8����  8����  ����Q  �      B  , ,��ˣ  s��ˣ  ���M  ���M  s��ˣ  s      B  , ,��·  s��·  ���1  ���1  s��·  s      B  , ,���k  s���k  ���  ���  s���k  s      B  , ,���O  s���O  ����  ����  s���O  s      B  , ,���3  s���3  ����  ����  s���3  s      B  , ,���  s���  ����  ����  s���  s      B  , ,����  s����  ��ݥ  ��ݥ  s����  s      B  , ,����  �����  <��Ӈ  <��Ӈ  �����  �      B  , ,����  �����  <���k  <���k  �����  �      B  , ,��إ  ���إ  <���O  <���O  ���إ  �      B  , ,��ۉ  ���ۉ  <���3  <���3  ���ۉ  �      B  , ,���m  ����m  <���  <���  ����m  �      B  , ,���1  >���1  �����  �����  >���1  >      B  , ,���  >���  ���Ϳ  ���Ϳ  >���  >      B  , ,����  >����  ���У  ���У  >����  >      B  , ,����  >����  ���Ӈ  ���Ӈ  >����  >      B  , ,����  >����  ����k  ����k  >����  >      B  , ,��إ  >��إ  ����O  ����O  >��إ  >      B  , ,��ۉ  >��ۉ  ����3  ����3  >��ۉ  >      B  , ,���m  >���m  ����  ����  >���m  >      B  , ,���Q  >���Q  �����  �����  >���Q  >      B  , ,���Q  ����Q  <����  <����  ����Q  �      B  , ,����  �����  ����k  ����k  �����  �      B  , ,��إ  ���إ  ����O  ����O  ���إ  �      B  , ,��ۉ  ���ۉ  ����3  ����3  ���ۉ  �      B  , ,���m  ����m  ����  ����  ����m  �      B  , ,���Q  ����Q  �����  �����  ����Q  �      B  , ,���1  ����1  �����  �����  ����1  �      B  , ,���  ����  ���Ϳ  ���Ϳ  ����  �      B  , ,����  �����  ���У  ���У  �����  �      B  , ,����  �����  ���Ӈ  ���Ӈ  �����  �      B  , ,���1  ����1  <����  <����  ����1  �      B  , ,���  ����  <��Ϳ  <��Ϳ  ����  �      B  , ,���1  ����1  �����  �����  ����1  �      B  , ,���  ����  ���Ϳ  ���Ϳ  ����  �      B  , ,����  �����  ���У  ���У  �����  �      B  , ,����  �����  ���Ӈ  ���Ӈ  �����  �      B  , ,����  �����  ����k  ����k  �����  �      B  , ,��إ  ���إ  ����O  ����O  ���إ  �      B  , ,��ۉ  ���ۉ  ����3  ����3  ���ۉ  �      B  , ,���m  ����m  ����  ����  ����m  �      B  , ,���Q  ����Q  �����  �����  ����Q  �      B  , ,����  �����  <��У  <��У  �����  �      B  , ,����  >����  ����o  ����o  >����  >      B  , ,���  >���  ����S  ����S  >���  >      B  , ,����  >����  ����7  ����7  >����  >      B  , ,���q  >���q  ����  ����  >���q  >      B  , ,���U  >���U  �����  �����  >���U  >      B  , ,���9  >���9  �����  �����  >���9  >      B  , ,����  �����  ����o  ����o  �����  �      B  , ,���  ����  <����  <����  ����  �      B  , ,����  �����  <���  <���  �����  �      B  , ,����  �����  <���  <���  �����  �      B  , ,����  �����  <���o  <���o  �����  �      B  , ,���  ����  <���S  <���S  ����  �      B  , ,����  �����  <���7  <���7  �����  �      B  , ,���q  ����q  <���  <���  ����q  �      B  , ,���U  ����U  <����  <����  ����U  �      B  , ,���9  ����9  <����  <����  ����9  �      B  , ,���  ����  ����S  ����S  ����  �      B  , ,����  �����  ����7  ����7  �����  �      B  , ,���q  ����q  ����  ����  ����q  �      B  , ,���U  ����U  �����  �����  ����U  �      B  , ,���9  ����9  �����  �����  ����9  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,���  >���  �����  �����  >���  >      B  , ,����  >����  ����  ����  >����  >      B  , ,����  >����  ����  ����  >����  >      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,����  �����  ����o  ����o  �����  �      B  , ,���  ����  ����S  ����S  ����  �      B  , ,����  �����  ����7  ����7  �����  �      B  , ,���q  ����q  ����  ����  ����q  �      B  , ,���U  ����U  �����  �����  ����U  �      B  , ,���9  ����9  �����  �����  ����9  �      B  , ,����  :����  �����  �����  :����  :      B  , ,����  :����  ����  ����  :����  :      B  , ,����  :����  ����c  ����c  :����  :      B  , ,����  :����  ����G  ����G  :����  :      B  , ,����  :����  ����+  ����+  :����  :      B  , ,���e  :���e  ����  ����  :���e  :      B  , ,���I  :���I  �����  �����  :���I  :      B  , ,���-  :���-  �����  �����  :���-  :      B  , ,���  :���  �����  �����  :���  :      B  , ,����  :����  �����  �����  :����  :      B  , ,����  :����  �����  �����  :����  :      B  , ,����  :����  ����g  ����g  :����  :      B  , ,����  :����  ����K  ����K  :����  :      B  , ,����  :����  ����/  ����/  :����  :      B  , ,���i  :���i  ����  ����  :���i  :      B  , ,���M  :���M  �����  �����  :���M  :      B  , ,���E  :���E  �����  �����  :���E  :      B  , ,���)  :���)  �����  �����  :���)  :      B  , ,���  :���  �����  �����  :���  :      B  , ,����  q����  ���S  ���S  q����  q      B  , ,���I  ����I  8����  8����  ����I  �      B  , ,���-  ����-  8����  8����  ����-  �      B  , ,���  ����  8����  8����  ����  �      B  , ,����  �����  8����  8����  �����  �      B  , ,����  �����  8����  8����  �����  �      B  , ,����  �����  8���g  8���g  �����  �      B  , ,����  �����  8���K  8���K  �����  �      B  , ,����  �����  8���/  8���/  �����  �      B  , ,���i  ����i  8���  8���  ����i  �      B  , ,���M  ����M  8����  8����  ����M  �      B  , ,����  s����  ��ƅ  ��ƅ  s����  s      B  , ,���=  q���=  ����  ����  q���=  q      B  , ,��đ  q��đ  ���;  ���;  q��đ  q      B  , ,����  s����  ���e  ���e  s����  s      B  , ,����  s����  ���I  ���I  s����  s      B  , ,����  s����  ���-  ���-  s����  s      B  , ,���g  s���g  ���  ���  s���g  s      B  , ,���K  s���K  ����  ����  s���K  s      B  , ,���/  s���/  ����  ����  s���/  s      B  , ,���9  q���9  ����  ����  q���9  q      B  , ,���  s���  ����  ����  s���  s      B  , ,����  s����  ��á  ��á  s����  s      B  , ,����  q����  ��Ə  ��Ə  q����  q      B  , ,����  q����  ����  ����  q����  q      B  , ,���Q  q���Q  ����  ����  q���Q  q      B  , ,����  q����  ���O  ���O  q����  q      B  , ,����  q����  ����  ����  q����  q      B  , ,���M  q���M  ����  ����  q���M  q      B  , ,����  q����  ���K  ���K  q����  q      B  , ,����  q����  ����  ����  q����  q      B  , ,���I  q���I  ����  ����  q���I  q      B  , ,����  q����  ���G  ���G  q����  q      B  , ,����  q����  ����  ����  q����  q      B  , ,���E  q���E  ����  ����  q���E  q      B  , ,����  q����  ���C  ���C  q����  q      B  , ,����  q����  ����  ����  q����  q      B  , ,���A  q���A  ����  ����  q���A  q      B  , ,����  q����  ���?  ���?  q����  q      B  , ,����  q����  ��  ��  q����  q      B  , ,����  �����  8���+  8���+  �����  �      B  , ,���e  ����e  8���  8���  ����e  �      B  , ,���  ����  C����  C����  ����  �      B  , ,���  ����  �����  �����  ����  �      B  , ,���m  q���m  ���  ���  q���m  q      B  , ,����  q����  ���k  ���k  q����  q      B  , ,���  q���  ����  ����  q���  q      B  , ,���i  q���i  ���  ���  q���i  q      B  , ,����  q����  ���g  ���g  q����  q      B  , ,���  q���  ����  ����  q���  q      B  , ,���e  q���e  ���  ���  q���e  q      B  , ,����  q����  ���c  ���c  q����  q      B  , ,���  q���  ����  ����  q���  q      B  , ,���a  q���a  ���  ���  q���a  q      B  , ,����  q����  ���_  ���_  q����  q      B  , ,���	  q���	  ����  ����  q���	  q      B  , ,���]  q���]  ���  ���  q���]  q      B  , ,����  q����  ���[  ���[  q����  q      B  , ,���  q���  ����  ����  q���  q      B  , ,���Y  q���Y  ���  ���  q���Y  q      B  , ,����  q����  ���W  ���W  q����  q      B  , ,���  q���  ����  ����  q���  q      B  , ,���U  q���U  ����  ����  q���U  q      B  , ,���E  ����E  8����  8����  ����E  �      B  , ,���)  ����)  8����  8����  ����)  �      B  , ,���  A���  �����  �����  A���  A      B  , ,����  s����  ���a  ���a  s����  s      B  , ,����  s����  ���E  ���E  s����  s      B  , ,���  s���  ���)  ���)  s���  s      B  , ,���c  s���c  ���  ���  s���c  s      B  , ,���G  s���G  ����  ����  s���G  s      B  , ,���+  s���+  ����  ����  s���+  s      B  , ,���  s���  ����  ����  s���  s      B  , ,����  s����  ����  ����  s����  s      B  , ,����  s����  ����  ����  s����  s      B  , ,���  ����  8����  8����  ����  �      B  , ,����  �����  8����  8����  �����  �      B  , ,����  �����  8���  8���  �����  �      B  , ,����  �����  8���c  8���c  �����  �      B  , ,����  �����  8���G  8���G  �����  �      B  , ,���e  >���e  ����  ����  >���e  >      B  , ,���E  ����E  �����  �����  ����E  �      B  , ,���  E���  �����  �����  E���  E      B  , ,���)  ����)  �����  �����  ����)  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,����  �����  ����c  ����c  �����  �      B  , ,����  �����  ����G  ����G  �����  �      B  , ,����  �����  ����+  ����+  �����  �      B  , ,���e  ����e  ����  ����  ����e  �      B  , ,���  ����  G����  G����  ����  �      B  , ,���E  >���E  �����  �����  >���E  >      B  , ,���)  >���)  �����  �����  >���)  >      B  , ,���  >���  �����  �����  >���  >      B  , ,����  >����  �����  �����  >����  >      B  , ,����  >����  ����  ����  >����  >      B  , ,���  I���  �����  �����  I���  I      B  , ,���E  ����E  �����  �����  ����E  �      B  , ,���)  ����)  �����  �����  ����)  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,����  �����  ����c  ����c  �����  �      B  , ,����  �����  ����G  ����G  �����  �      B  , ,����  �����  ����+  ����+  �����  �      B  , ,���e  ����e  ����  ����  ����e  �      B  , ,����  >����  ����c  ����c  >����  >      B  , ,����  >����  ����G  ����G  >����  >      B  , ,����  >����  ����+  ����+  >����  >      B  , ,���  ����  �����  �����  ����  �      B  , ,���E  ����E  <����  <����  ����E  �      B  , ,���)  ����)  <����  <����  ����)  �      B  , ,���  ����  <����  <����  ����  �      B  , ,����  �����  <����  <����  �����  �      B  , ,����  �����  <���  <���  �����  �      B  , ,����  �����  <���c  <���c  �����  �      B  , ,����  �����  <���G  <���G  �����  �      B  , ,����  �����  <���+  <���+  �����  �      B  , ,���e  ����e  <���  <���  ����e  �      B  , ,���-  ����-  �����  �����  ����-  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  ����g  ����g  �����  �      B  , ,���I  >���I  �����  �����  >���I  >      B  , ,���-  >���-  �����  �����  >���-  >      B  , ,���  >���  �����  �����  >���  >      B  , ,����  >����  �����  �����  >����  >      B  , ,����  >����  �����  �����  >����  >      B  , ,����  >����  ����g  ����g  >����  >      B  , ,���I  ����I  �����  �����  ����I  �      B  , ,���-  ����-  �����  �����  ����-  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  ����g  ����g  �����  �      B  , ,����  �����  ����K  ����K  �����  �      B  , ,����  �����  ����/  ����/  �����  �      B  , ,���i  ����i  ����  ����  ����i  �      B  , ,���M  ����M  �����  �����  ����M  �      B  , ,����  >����  ����K  ����K  >����  >      B  , ,����  >����  ����/  ����/  >����  >      B  , ,���i  >���i  ����  ����  >���i  >      B  , ,���M  >���M  �����  �����  >���M  >      B  , ,���i  ����i  ����  ����  ����i  �      B  , ,���M  ����M  �����  �����  ����M  �      B  , ,����  �����  ����K  ����K  �����  �      B  , ,����  �����  ����/  ����/  �����  �      B  , ,���i  ����i  <���  <���  ����i  �      B  , ,���M  ����M  <����  <����  ����M  �      B  , ,����  �����  <���K  <���K  �����  �      B  , ,����  �����  <���/  <���/  �����  �      B  , ,���I  ����I  �����  �����  ����I  �      B  , ,���I  ����I  <����  <����  ����I  �      B  , ,���-  ����-  <����  <����  ����-  �      B  , ,���  ����  <����  <����  ����  �      B  , ,����  �����  <����  <����  �����  �      B  , ,����  �����  <����  <����  �����  �      B  , ,����  �����  <���g  <���g  �����  �      B  , ,���  ����  O����  O����  ����  �      B  , ,���E  F���E  �����  �����  F���E  F      B  , ,���)  F���)  �����  �����  F���)  F      B  , ,���  F���  �����  �����  F���  F      B  , ,����  F����  �����  �����  F����  F      B  , ,����  F����  ����  ����  F����  F      B  , ,����  F����  ����c  ����c  F����  F      B  , ,����  F����  ����G  ����G  F����  F      B  , ,����  F����  ����+  ����+  F����  F      B  , ,���e  F���e  ����  ����  F���e  F      B  , ,���I  F���I  �����  �����  F���I  F      B  , ,���-  F���-  �����  �����  F���-  F      B  , ,���  F���  �����  �����  F���  F      B  , ,����  F����  �����  �����  F����  F      B  , ,����  F����  �����  �����  F����  F      B  , ,����  F����  ����g  ����g  F����  F      B  , ,����  F����  ����K  ����K  F����  F      B  , ,����  F����  ����/  ����/  F����  F      B  , ,���i  F���i  ����  ����  F���i  F      B  , ,���M  F���M  �����  �����  F���M  F      B  , ,���I  ����I  �����  �����  ����I  �      B  , ,���-  ����-  �����  �����  ����-  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  ����g  ����g  �����  �      B  , ,����  �����  ����K  ����K  �����  �      B  , ,����  �����  ����/  ����/  �����  �      B  , ,���i  ����i  ����  ����  ����i  �      B  , ,���M  ����M  �����  �����  ����M  �      B  , ,���I  
����I  @����  @����  
����I  
�      B  , ,���-  
����-  @����  @����  
����-  
�      B  , ,���  
����  @����  @����  
����  
�      B  , ,����  
�����  @����  @����  
�����  
�      B  , ,����  
�����  @����  @����  
�����  
�      B  , ,����  
�����  @���g  @���g  
�����  
�      B  , ,����  
�����  @���K  @���K  
�����  
�      B  , ,����  
�����  @���/  @���/  
�����  
�      B  , ,���i  
����i  @���  @���  
����i  
�      B  , ,���M  
����M  @����  @����  
����M  
�      B  , ,���I  	B���I  	�����  	�����  	B���I  	B      B  , ,���-  	B���-  	�����  	�����  	B���-  	B      B  , ,���  	B���  	�����  	�����  	B���  	B      B  , ,����  	B����  	�����  	�����  	B����  	B      B  , ,����  	B����  	�����  	�����  	B����  	B      B  , ,����  	B����  	����g  	����g  	B����  	B      B  , ,����  	B����  	����K  	����K  	B����  	B      B  , ,����  	B����  	����/  	����/  	B����  	B      B  , ,���i  	B���i  	����  	����  	B���i  	B      B  , ,���M  	B���M  	�����  	�����  	B���M  	B      B  , ,���I  ����I  D����  D����  ����I  �      B  , ,���-  ����-  D����  D����  ����-  �      B  , ,���  ����  D����  D����  ����  �      B  , ,����  �����  D����  D����  �����  �      B  , ,����  �����  D����  D����  �����  �      B  , ,����  �����  D���g  D���g  �����  �      B  , ,����  �����  D���K  D���K  �����  �      B  , ,����  �����  D���/  D���/  �����  �      B  , ,���i  ����i  D���  D���  ����i  �      B  , ,���M  ����M  D����  D����  ����M  �      B  , ,���E  	B���E  	�����  	�����  	B���E  	B      B  , ,���)  	B���)  	�����  	�����  	B���)  	B      B  , ,���  	B���  	�����  	�����  	B���  	B      B  , ,����  	B����  	�����  	�����  	B����  	B      B  , ,����  	B����  	����  	����  	B����  	B      B  , ,����  	B����  	����c  	����c  	B����  	B      B  , ,����  	B����  	����G  	����G  	B����  	B      B  , ,����  	B����  	����+  	����+  	B����  	B      B  , ,���e  	B���e  	����  	����  	B���e  	B      B  , ,���  
����  @����  @����  
����  
�      B  , ,����  
�����  @����  @����  
�����  
�      B  , ,����  
�����  @���  @���  
�����  
�      B  , ,����  
�����  @���c  @���c  
�����  
�      B  , ,����  
�����  @���G  @���G  
�����  
�      B  , ,����  
�����  @���+  @���+  
�����  
�      B  , ,���e  
����e  @���  @���  
����e  
�      B  , ,���  M���  �����  �����  M���  M      B  , ,���E  ����E  �����  �����  ����E  �      B  , ,���)  ����)  �����  �����  ����)  �      B  , ,���  ����  �����  �����  ����  �      B  , ,���E  ����E  D����  D����  ����E  �      B  , ,���)  ����)  D����  D����  ����)  �      B  , ,���  ����  D����  D����  ����  �      B  , ,����  �����  D����  D����  �����  �      B  , ,����  �����  D���  D���  �����  �      B  , ,����  �����  D���c  D���c  �����  �      B  , ,����  �����  D���G  D���G  �����  �      B  , ,����  �����  D���+  D���+  �����  �      B  , ,���e  ����e  D���  D���  ����e  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,����  �����  ����c  ����c  �����  �      B  , ,����  �����  ����G  ����G  �����  �      B  , ,����  �����  ����+  ����+  �����  �      B  , ,���e  ����e  ����  ����  ����e  �      B  , ,���E  
����E  @����  @����  
����E  
�      B  , ,���)  
����)  @����  @����  
����)  
�      B  , ,���  	����  
K����  
K����  	����  	�      B  , ,���  ����  �����  �����  ����  �      B  , ,���E  ����E  H����  H����  ����E  �      B  , ,���)  ����)  H����  H����  ����)  �      B  , ,���  ����  H����  H����  ����  �      B  , ,����  �����  H����  H����  �����  �      B  , ,����  �����  H���  H���  �����  �      B  , ,����  �����  H���c  H���c  �����  �      B  , ,����  �����  H���G  H���G  �����  �      B  , ,����  �����  H���+  H���+  �����  �      B  , ,���  ����  S����  S����  ����  �      B  , ,���e  ����e  H���  H���  ����e  �      B  , ,���   U���   �����   �����   U���   U      B  , ,����   �����  c���a  c���a   �����   �      B  , ,����   �����  c���E  c���E   �����   �      B  , ,���   ����  c���)  c���)   ����   �      B  , ,���c   ����c  c���  c���   ����c   �      B  , ,���G   ����G  c����  c����   ����G   �      B  , ,���+   ����+  c����  c����   ����+   �      B  , ,���   ����  c����  c����   ����   �      B  , ,����   �����  c����  c����   �����   �      B  , ,���  Q���  �����  �����  Q���  Q      B  , ,���E  ����E  �����  �����  ����E  �      B  , ,���)  ����)  �����  �����  ����)  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,����  �����  ����c  ����c  �����  �      B  , ,����  �����  ����G  ����G  �����  �      B  , ,����  �����  ����+  ����+  �����  �      B  , ,���e  ����e  ����  ����  ����e  �      B  , ,����   �����  c����  c����   �����   �      B  , ,����   �����  c���-  c���-   �����   �      B  , ,���g   ����g  c���  c���   ����g   �      B  , ,���K   ����K  c����  c����   ����K   �      B  , ,���/   ����/  c����  c����   ����/   �      B  , ,���   ����  c����  c����   ����   �      B  , ,����   �����  c��á  c��á   �����   �      B  , ,����   �����  c��ƅ  c��ƅ   �����   �      B  , ,���-  ����-  H����  H����  ����-  �      B  , ,���  ����  H����  H����  ����  �      B  , ,����  �����  H����  H����  �����  �      B  , ,����  �����  H����  H����  �����  �      B  , ,����  �����  H���g  H���g  �����  �      B  , ,����  �����  H���K  H���K  �����  �      B  , ,����  �����  H���/  H���/  �����  �      B  , ,���i  ����i  H���  H���  ����i  �      B  , ,���M  ����M  H����  H����  ����M  �      B  , ,���I  ����I  H����  H����  ����I  �      B  , ,����   �����  c���e  c���e   �����   �      B  , ,���I  ����I  �����  �����  ����I  �      B  , ,���-  ����-  �����  �����  ����-  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,����  �����  ����g  ����g  �����  �      B  , ,����  �����  ����K  ����K  �����  �      B  , ,����  �����  ����/  ����/  �����  �      B  , ,���i  ����i  ����  ����  ����i  �      B  , ,���M  ����M  �����  �����  ����M  �      B  , ,����   �����  c���I  c���I   �����   �      B  , ,���5  	B���5  	�����  	�����  	B���5  	B      B  , ,���5  ����5  H����  H����  ����5  �      B  , ,���5  
����5  @����  @����  
����5  
�      B  , ,���5  ����5  �����  �����  ����5  �      B  , ,���5  ����5  �����  �����  ����5  �      B  , ,���1  F���1  �����  �����  F���1  F      B  , ,���  F���  ���Ϳ  ���Ϳ  F���  F      B  , ,����  F����  ���У  ���У  F����  F      B  , ,����  F����  ���Ӈ  ���Ӈ  F����  F      B  , ,����  F����  ����k  ����k  F����  F      B  , ,��إ  F��إ  ����O  ����O  F��إ  F      B  , ,��ۉ  F��ۉ  ����3  ����3  F��ۉ  F      B  , ,���m  F���m  ����  ����  F���m  F      B  , ,���Q  F���Q  �����  �����  F���Q  F      B  , ,���5  F���5  �����  �����  F���5  F      B  , ,���  F���  �����  �����  F���  F      B  , ,����  F����  ����  ����  F����  F      B  , ,����  F����  ����  ����  F����  F      B  , ,����  F����  ����o  ����o  F����  F      B  , ,���  F���  ����S  ����S  F���  F      B  , ,����  F����  ����7  ����7  F����  F      B  , ,���q  F���q  ����  ����  F���q  F      B  , ,���U  F���U  �����  �����  F���U  F      B  , ,���9  F���9  �����  �����  F���9  F      B  , ,���5  ����5  D����  D����  ����5  �      B  , ,���q  
����q  @���  @���  
����q  
�      B  , ,���U  
����U  @����  @����  
����U  
�      B  , ,���9  
����9  @����  @����  
����9  
�      B  , ,����  �����  D���7  D���7  �����  �      B  , ,���q  ����q  D���  D���  ����q  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,����  �����  ����o  ����o  �����  �      B  , ,���  ����  ����S  ����S  ����  �      B  , ,����  �����  ����7  ����7  �����  �      B  , ,���q  ����q  ����  ����  ����q  �      B  , ,���U  ����U  �����  �����  ����U  �      B  , ,���9  ����9  �����  �����  ����9  �      B  , ,���U  ����U  D����  D����  ����U  �      B  , ,���9  ����9  D����  D����  ����9  �      B  , ,����  �����  D���  D���  �����  �      B  , ,����  �����  D���o  D���o  �����  �      B  , ,���  	B���  	�����  	�����  	B���  	B      B  , ,����  	B����  	����  	����  	B����  	B      B  , ,����  	B����  	����  	����  	B����  	B      B  , ,����  	B����  	����o  	����o  	B����  	B      B  , ,���  	B���  	����S  	����S  	B���  	B      B  , ,����  	B����  	����7  	����7  	B����  	B      B  , ,���q  	B���q  	����  	����  	B���q  	B      B  , ,���U  	B���U  	�����  	�����  	B���U  	B      B  , ,���9  	B���9  	�����  	�����  	B���9  	B      B  , ,���  ����  D���S  D���S  ����  �      B  , ,���  
����  @����  @����  
����  
�      B  , ,����  
�����  @���  @���  
�����  
�      B  , ,����  
�����  @���  @���  
�����  
�      B  , ,����  
�����  @���o  @���o  
�����  
�      B  , ,���  
����  @���S  @���S  
����  
�      B  , ,����  
�����  @���7  @���7  
�����  
�      B  , ,���  ����  D����  D����  ����  �      B  , ,����  �����  D���  D���  �����  �      B  , ,����  
�����  @��Ӈ  @��Ӈ  
�����  
�      B  , ,����  
�����  @���k  @���k  
�����  
�      B  , ,��إ  
���إ  @���O  @���O  
���إ  
�      B  , ,����  	B����  	���У  	���У  	B����  	B      B  , ,����  	B����  	���Ӈ  	���Ӈ  	B����  	B      B  , ,���1  ����1  D����  D����  ����1  �      B  , ,���  ����  D��Ϳ  D��Ϳ  ����  �      B  , ,��ۉ  
���ۉ  @���3  @���3  
���ۉ  
�      B  , ,���1  
����1  @����  @����  
����1  
�      B  , ,���  
����  @��Ϳ  @��Ϳ  
����  
�      B  , ,���1  	B���1  	�����  	�����  	B���1  	B      B  , ,���  	B���  	���Ϳ  	���Ϳ  	B���  	B      B  , ,���1  ����1  �����  �����  ����1  �      B  , ,���  ����  ���Ϳ  ���Ϳ  ����  �      B  , ,����  �����  ���У  ���У  �����  �      B  , ,����  �����  ���Ӈ  ���Ӈ  �����  �      B  , ,����  �����  ����k  ����k  �����  �      B  , ,��إ  ���إ  ����O  ����O  ���إ  �      B  , ,���m  
����m  @���  @���  
����m  
�      B  , ,��ۉ  ���ۉ  ����3  ����3  ���ۉ  �      B  , ,���m  ����m  ����  ����  ����m  �      B  , ,���Q  ����Q  �����  �����  ����Q  �      B  , ,���Q  
����Q  @����  @����  
����Q  
�      B  , ,��إ  	B��إ  	����O  	����O  	B��إ  	B      B  , ,��ۉ  	B��ۉ  	����3  	����3  	B��ۉ  	B      B  , ,���m  	B���m  	����  	����  	B���m  	B      B  , ,����  �����  D��У  D��У  �����  �      B  , ,����  �����  D��Ӈ  D��Ӈ  �����  �      B  , ,����  �����  D���k  D���k  �����  �      B  , ,��إ  ���إ  D���O  D���O  ���إ  �      B  , ,��ۉ  ���ۉ  D���3  D���3  ���ۉ  �      B  , ,���m  ����m  D���  D���  ����m  �      B  , ,���Q  ����Q  D����  D����  ����Q  �      B  , ,���Q  	B���Q  	�����  	�����  	B���Q  	B      B  , ,����  	B����  	����k  	����k  	B����  	B      B  , ,����  
�����  @��У  @��У  
�����  
�      B  , ,����  �����  H��У  H��У  �����  �      B  , ,����  �����  H��Ӈ  H��Ӈ  �����  �      B  , ,����  �����  H���k  H���k  �����  �      B  , ,��إ  ���إ  H���O  H���O  ���إ  �      B  , ,��ۉ  ���ۉ  H���3  H���3  ���ۉ  �      B  , ,��ȿ   ���ȿ  c���i  c���i   ���ȿ   �      B  , ,��ˣ   ���ˣ  c���M  c���M   ���ˣ   �      B  , ,��·   ���·  c���1  c���1   ���·   �      B  , ,���k   ����k  c���  c���   ����k   �      B  , ,���O   ����O  c����  c����   ����O   �      B  , ,���3   ����3  c����  c����   ����3   �      B  , ,���   ����  c����  c����   ����   �      B  , ,����   �����  c��ݥ  c��ݥ   �����   �      B  , ,����   �����  c����  c����   �����   �      B  , ,����   �����  c���m  c���m   �����   �      B  , ,���m  ����m  H���  H���  ����m  �      B  , ,���Q  ����Q  H����  H����  ����Q  �      B  , ,���1  ����1  H����  H����  ����1  �      B  , ,���1  ����1  �����  �����  ����1  �      B  , ,���  ����  ���Ϳ  ���Ϳ  ����  �      B  , ,����  �����  ���У  ���У  �����  �      B  , ,����  �����  ���Ӈ  ���Ӈ  �����  �      B  , ,����  �����  ����k  ����k  �����  �      B  , ,��إ  ���إ  ����O  ����O  ���إ  �      B  , ,��ۉ  ���ۉ  ����3  ����3  ���ۉ  �      B  , ,���m  ����m  ����  ����  ����m  �      B  , ,���Q  ����Q  �����  �����  ����Q  �      B  , ,���  ����  H��Ϳ  H��Ϳ  ����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,����  �����  ����o  ����o  �����  �      B  , ,���  ����  ����S  ����S  ����  �      B  , ,����  �����  ����7  ����7  �����  �      B  , ,���   ����  c���Q  c���Q   ����   �      B  , ,���   ����  c���5  c���5   ����   �      B  , ,���o   ����o  c���  c���   ����o   �      B  , ,���S   ����S  c����  c����   ����S   �      B  , ,���7   ����7  c����  c����   ����7   �      B  , ,���   ����  c����  c����   ����   �      B  , ,����   �����  c����  c����   �����   �      B  , ,����   �����  c����  c����   �����   �      B  , ,����   �����  c���q  c���q   �����   �      B  , ,���q  ����q  ����  ����  ����q  �      B  , ,���U  ����U  �����  �����  ����U  �      B  , ,���9  ����9  �����  �����  ����9  �      B  , ,����  �����  H���  H���  �����  �      B  , ,����  �����  H���  H���  �����  �      B  , ,����  �����  H���o  H���o  �����  �      B  , ,���  ����  H���S  H���S  ����  �      B  , ,����  �����  H���7  H���7  �����  �      B  , ,���q  ����q  H���  H���  ����q  �      B  , ,���U  ����U  H����  H����  ����U  �      B  , ,���9  ����9  H����  H����  ����9  �      B  , ,���  ����  H����  H����  ����  �      B  , ,���  ����  �����  �����  ����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,������a��������������������a������a      B  , ,���5�������5���b�������b�����������5����      B  , ,���5���d���5�����������������d���5���d      B  , ,���1������1����������������������1���      B  , ,���������������Ϳ������Ϳ���������      B  , ,�����������������У������У����������      B  , ,�����������������Ӈ������Ӈ����������      B  , ,������������������k�������k����������      B  , ,��إ�����إ�������O�������O�����إ���      B  , ,��ۉ�����ۉ�������3�������3�����ۉ���      B  , ,���m������m��������������������m���      B  , ,���Q������Q����������������������Q���      B  , ,���5������5����������������������5���      B  , ,����������������������������������      B  , ,�����������������������������������      B  , ,�����������������������������������      B  , ,������������������o�������o����������      B  , ,����������������S�������S���������      B  , ,������������������7�������7����������      B  , ,���q������q��������������������q���      B  , ,���U������U����������������������U���      B  , ,���9������9����������������������9���      B  , ,���5�������5���f�������f�����������5����      B  , ,���5���h���5�����������������h���5���h      B  , ,���5������5����������������������5���      B  , ,���5�������5���j�������j�����������5����      B  , ,�������d����������7������7���d�������d      B  , ,���q���d���q���������������d���q���d      B  , ,���U���d���U�����������������d���U���d      B  , ,���9���d���9�����������������d���9���d      B  , ,���o�������o���G������G����������o����      B  , ,���S�������S���G�������G�����������S����      B  , ,���7�������7���G�������G�����������7����      B  , ,�������������G�������G���������������      B  , ,���������������G�������G����������������      B  , ,���������������G�������G����������������      B  , ,���������������G���q���G���q������������      B  , ,�������������G���Q���G���Q�����������      B  , ,�������������b�������b���������������      B  , ,���������������b������b���������������      B  , ,���������������b������b���������������      B  , ,���������������b���o���b���o������������      B  , ,�������������b���S���b���S�����������      B  , ,���������������b���7���b���7������������      B  , ,���q�������q���b������b����������q����      B  , ,���U�������U���b�������b�����������U����      B  , ,���9�������9���b�������b�����������9����      B  , ,�������������G���5���G���5�����������      B  , ,������d��������������������d������d      B  , ,�������d�������������������d�������d      B  , ,�������d�������������������d�������d      B  , ,�������d����������o������o���d�������d      B  , ,������d���������S������S���d������d      B  , ,���m�������m���b������b����������m����      B  , ,���Q�������Q���b�������b�����������Q����      B  , ,��ˣ������ˣ���G���M���G���M������ˣ����      B  , ,��·������·���G���1���G���1������·����      B  , ,���k�������k���G������G����������k����      B  , ,���O�������O���G�������G�����������O����      B  , ,���3�������3���G�������G�����������3����      B  , ,�������������G�������G���������������      B  , ,���������������G��ݥ���G��ݥ������������      B  , ,���������������G�������G����������������      B  , ,���������������G���m���G���m������������      B  , ,���1�������1���b�������b�����������1����      B  , ,���1���d���1�����������������d���1���d      B  , ,������d��������Ϳ�����Ϳ���d������d      B  , ,�������d���������У�����У���d�������d      B  , ,�������d���������Ӈ�����Ӈ���d�������d      B  , ,�������d����������k������k���d�������d      B  , ,��إ���d��إ������O������O���d��إ���d      B  , ,��ۉ���d��ۉ������3������3���d��ۉ���d      B  , ,���m���d���m���������������d���m���d      B  , ,���Q���d���Q�����������������d���Q���d      B  , ,�������������b��Ϳ���b��Ϳ�����������      B  , ,���������������b��У���b��У������������      B  , ,���������������b��Ӈ���b��Ӈ������������      B  , ,���������������b���k���b���k������������      B  , ,��إ������إ���b���O���b���O������إ����      B  , ,��ȿ������ȿ���G���i���G���i������ȿ����      B  , ,��ۉ������ۉ���b���3���b���3������ۉ����      B  , ,��إ������إ���f���O���f���O������إ����      B  , ,��ۉ������ۉ���f���3���f���3������ۉ����      B  , ,���m�������m���f������f����������m����      B  , ,���Q�������Q���f�������f�����������Q����      B  , ,���1�������1���f�������f�����������1����      B  , ,���1���h���1�����������������h���1���h      B  , ,������h��������Ϳ�����Ϳ���h������h      B  , ,�������h���������У�����У���h�������h      B  , ,�������h���������Ӈ�����Ӈ���h�������h      B  , ,�������h����������k������k���h�������h      B  , ,��إ���h��إ������O������O���h��إ���h      B  , ,��ۉ���h��ۉ������3������3���h��ۉ���h      B  , ,���m���h���m���������������h���m���h      B  , ,���Q���h���Q�����������������h���Q���h      B  , ,�������������f��Ϳ���f��Ϳ�����������      B  , ,���1������1����������������������1���      B  , ,���������������Ϳ������Ϳ���������      B  , ,�����������������У������У����������      B  , ,�����������������Ӈ������Ӈ����������      B  , ,������������������k�������k����������      B  , ,��إ�����إ�������O�������O�����إ���      B  , ,��ۉ�����ۉ�������3�������3�����ۉ���      B  , ,���m������m��������������������m���      B  , ,���Q������Q����������������������Q���      B  , ,���������������f��У���f��У������������      B  , ,���������������f��Ӈ���f��Ӈ������������      B  , ,���1�������1���j�������j�����������1����      B  , ,�������������j��Ϳ���j��Ϳ�����������      B  , ,���������������j��У���j��У������������      B  , ,���������������j��Ӈ���j��Ӈ������������      B  , ,���������������j���k���j���k������������      B  , ,��إ������إ���j���O���j���O������إ����      B  , ,��ۉ������ۉ���j���3���j���3������ۉ����      B  , ,���m�������m���j������j����������m����      B  , ,���Q�������Q���j�������j�����������Q����      B  , ,���������������f���k���f���k������������      B  , ,�������������f���S���f���S�����������      B  , ,���������������f���7���f���7������������      B  , ,���q�������q���f������f����������q����      B  , ,���U�������U���f�������f�����������U����      B  , ,���9�������9���f�������f�����������9����      B  , ,�������������f�������f���������������      B  , ,������h��������������������h������h      B  , ,����������������������������������      B  , ,�����������������������������������      B  , ,�����������������������������������      B  , ,������������������o�������o����������      B  , ,����������������S�������S���������      B  , ,������������������7�������7����������      B  , ,���q������q��������������������q���      B  , ,���U������U����������������������U���      B  , ,���9������9����������������������9���      B  , ,�������h�������������������h�������h      B  , ,�������h�������������������h�������h      B  , ,�������h����������o������o���h�������h      B  , ,������h���������S������S���h������h      B  , ,�������h����������7������7���h�������h      B  , ,���q���h���q���������������h���q���h      B  , ,���U���h���U�����������������h���U���h      B  , ,���9���h���9�����������������h���9���h      B  , ,���������������f������f���������������      B  , ,���������������f������f���������������      B  , ,���������������f���o���f���o������������      B  , ,�������������j�������j���������������      B  , ,���������������j������j���������������      B  , ,���������������j������j���������������      B  , ,���������������j���o���j���o������������      B  , ,�������������j���S���j���S�����������      B  , ,���������������j���7���j���7������������      B  , ,���q�������q���j������j����������q����      B  , ,���U�������U���j�������j�����������U����      B  , ,���9�������9���j�������j�����������9����      B  , ,�������������[�������[���������������      B  , ,���E������E����������������������E���      B  , ,���)������)����������������������)���      B  , ,����������������������������������      B  , ,�������������������������������������      B  , ,�����������������������������������      B  , ,������������������c�������c����������      B  , ,������������������G�������G����������      B  , ,������������������+�������+����������      B  , ,���e������e��������������������e���      B  , ,���I������I����������������������I���      B  , ,���-������-����������������������-���      B  , ,����������������������������������      B  , ,�������������������������������������      B  , ,�������������������������������������      B  , ,������������������g�������g����������      B  , ,������������������K�������K����������      B  , ,������������������/�������/����������      B  , ,���i������i��������������������i���      B  , ,���M������M����������������������M���      B  , ,���-���d���-�����������������d���-���d      B  , ,������d��������������������d������d      B  , ,�������d���������������������d�������d      B  , ,�������d���������������������d�������d      B  , ,�������d����������g������g���d�������d      B  , ,�������d����������K������K���d�������d      B  , ,�������d����������/������/���d�������d      B  , ,���i���d���i���������������d���i���d      B  , ,���M���d���M�����������������d���M���d      B  , ,���I�������I���b�������b�����������I����      B  , ,���-�������-���b�������b�����������-����      B  , ,�������������b�������b���������������      B  , ,���������������b�������b����������������      B  , ,���������������b�������b����������������      B  , ,���������������b���g���b���g������������      B  , ,���������������b���K���b���K������������      B  , ,���������������b���/���b���/������������      B  , ,���i�������i���b������b����������i����      B  , ,���I���d���I�����������������d���I���d      B  , ,���M�������M���b�������b�����������M����      B  , ,���������������G���e���G���e������������      B  , ,���������������G���I���G���I������������      B  , ,���������������G���-���G���-������������      B  , ,���g�������g���G������G����������g����      B  , ,���K�������K���G�������G�����������K����      B  , ,���/�������/���G�������G�����������/����      B  , ,�������������G�������G���������������      B  , ,���������������G��á���G��á������������      B  , ,���������������G��ƅ���G��ƅ������������      B  , ,�������������b�������b���������������      B  , ,���������������b�������b����������������      B  , ,���������������b������b���������������      B  , ,���������������b���c���b���c������������      B  , ,���������������b���G���b���G������������      B  , ,���������������b���+���b���+������������      B  , ,���e�������e���b������b����������e����      B  , ,�������d����������G������G���d�������d      B  , ,�������d����������+������+���d�������d      B  , ,���e���d���e���������������d���e���d      B  , ,�������������G���)���G���)�����������      B  , ,����������������������������������      B  , ,�������������W�������W���������������      B  , ,����������������������������������      B  , ,���c�������c���G������G����������c����      B  , ,���G�������G���G�������G�����������G����      B  , ,���+�������+���G�������G�����������+����      B  , ,�������������G�������G���������������      B  , ,���������������G�������G����������������      B  , ,���������������G�������G����������������      B  , ,���E���d���E�����������������d���E���d      B  , ,���)���d���)�����������������d���)���d      B  , ,������d��������������������d������d      B  , ,�������d���������������������d�������d      B  , ,�������d�������������������d�������d      B  , ,�������d����������c������c���d�������d      B  , ,������Y��������������������Y������Y      B  , ,���E�������E���b�������b�����������E����      B  , ,���)�������)���b�������b�����������)����      B  , ,���������������G���E���G���E������������      B  , ,���������������G���a���G���a������������      B  , ,���������������f���+���f���+������������      B  , ,������	����������������������	������	      B  , ,���E���h���E�����������������h���E���h      B  , ,���)���h���)�����������������h���)���h      B  , ,������h��������������������h������h      B  , ,�������h���������������������h�������h      B  , ,�������h�������������������h�������h      B  , ,�������h����������c������c���h�������h      B  , ,�������h����������G������G���h�������h      B  , ,�������h����������+������+���h�������h      B  , ,���E�������E���j�������j�����������E����      B  , ,���)�������)���j�������j�����������)����      B  , ,�������������j�������j���������������      B  , ,���������������j�������j����������������      B  , ,���������������j������j���������������      B  , ,���������������j���c���j���c������������      B  , ,���������������j���G���j���G������������      B  , ,���������������j���+���j���+������������      B  , ,���e�������e���j������j����������e����      B  , ,�������������_�������_���������������      B  , ,���E������E����������������������E���      B  , ,���)������)����������������������)���      B  , ,����������������������������������      B  , ,�������������������������������������      B  , ,�����������������������������������      B  , ,������������������c�������c����������      B  , ,������������������G�������G����������      B  , ,������������������+�������+����������      B  , ,���e������e��������������������e���      B  , ,���e���h���e���������������h���e���h      B  , ,���e�������e���f������f����������e����      B  , ,������]��������������������]������]      B  , ,���E�������E���f�������f�����������E����      B  , ,���)�������)���f�������f�����������)����      B  , ,�������������f�������f���������������      B  , ,���������������f�������f����������������      B  , ,���������������f������f���������������      B  , ,���������������f���c���f���c������������      B  , ,���������������f���G���f���G������������      B  , ,���������������f���/���f���/������������      B  , ,���I������I����������������������I���      B  , ,���-������-����������������������-���      B  , ,����������������������������������      B  , ,�������������������������������������      B  , ,�������������������������������������      B  , ,������������������g�������g����������      B  , ,������������������K�������K����������      B  , ,������������������/�������/����������      B  , ,���i������i��������������������i���      B  , ,���I�������I���j�������j�����������I����      B  , ,���-�������-���j�������j�����������-����      B  , ,�������������j�������j���������������      B  , ,���������������j�������j����������������      B  , ,���������������j�������j����������������      B  , ,���������������j���g���j���g������������      B  , ,���������������j���K���j���K������������      B  , ,���������������j���/���j���/������������      B  , ,���i�������i���j������j����������i����      B  , ,���M�������M���j�������j�����������M����      B  , ,���M������M����������������������M���      B  , ,���i�������i���f������f����������i����      B  , ,���I���h���I�����������������h���I���h      B  , ,���-���h���-�����������������h���-���h      B  , ,������h��������������������h������h      B  , ,�������h���������������������h�������h      B  , ,�������h���������������������h�������h      B  , ,�������h����������g������g���h�������h      B  , ,�������h����������K������K���h�������h      B  , ,�������h����������/������/���h�������h      B  , ,���i���h���i���������������h���i���h      B  , ,���M���h���M�����������������h���M���h      B  , ,���M�������M���f�������f�����������M����      B  , ,���I�������I���f�������f�����������I����      B  , ,���-�������-���f�������f�����������-����      B  , ,�������������f�������f���������������      B  , ,���������������f�������f����������������      B  , ,���������������f�������f����������������      B  , ,���������������f���g���f���g������������      B  , ,���������������f���K���f���K������������      B  , ,���E������E����������������������E���      B  , ,���)������)����������������������)���      B  , ,����������������������������������      B  , ,�������������������������������������      B  , ,�����������������������������������      B  , ,������������������c�������c����������      B  , ,������������������G�������G����������      B  , ,������������������+�������+����������      B  , ,���e������e��������������������e���      B  , ,���I������I����������������������I���      B  , ,���-������-����������������������-���      B  , ,����������������������������������      B  , ,�������������������������������������      B  , ,�������������������������������������      B  , ,������������������g�������g����������      B  , ,������������������K�������K����������      B  , ,������������������/�������/����������      B  , ,���i������i��������������������i���      B  , ,���M������M����������������������M���      B  , ,������������������S������S������������      B  , ,���I�������I���n�������n�����������I����      B  , ,���-�������-���n�������n�����������-����      B  , ,�������������n�������n���������������      B  , ,���������������n�������n����������������      B  , ,���������������n�������n����������������      B  , ,���������������n���g���n���g������������      B  , ,���������������n���K���n���K������������      B  , ,���������������n���/���n���/������������      B  , ,���i�������i���n������n����������i����      B  , ,���M�������M���n�������n�����������M����      B  , ,���I���p���I�����������������p���I���p      B  , ,���-���p���-�����������������p���-���p      B  , ,������p��������������������p������p      B  , ,�������p���������������������p�������p      B  , ,�������p���������������������p�������p      B  , ,�������p����������g������g���p�������p      B  , ,�������p����������K������K���p�������p      B  , ,�������p����������/������/���p�������p      B  , ,���i���p���i���������������p���i���p      B  , ,���M���p���M�����������������p���M���p      B  , ,���I���l���I�����������������l���I���l      B  , ,���-���l���-�����������������l���-���l      B  , ,������l��������������������l������l      B  , ,�������l���������������������l�������l      B  , ,�������l���������������������l�������l      B  , ,�������l����������g������g���l�������l      B  , ,�������l����������K������K���l�������l      B  , ,�������l����������/������/���l�������l      B  , ,���i���l���i���������������l���i���l      B  , ,���M���l���M�����������������l���M���l      B  , ,���I������I����������������������I���      B  , ,���-������-����������������������-���      B  , ,����������������������������������      B  , ,�������������������������������������      B  , ,�������������������������������������      B  , ,������������������g�������g����������      B  , ,������������������K�������K����������      B  , ,������������������/�������/����������      B  , ,���i������i��������������������i���      B  , ,���M������M����������������������M���      B  , ,���E���p���E�����������������p���E���p      B  , ,���)���p���)�����������������p���)���p      B  , ,������p��������������������p������p      B  , ,�������p���������������������p�������p      B  , ,�������p�������������������p�������p      B  , ,�������p����������c������c���p�������p      B  , ,�������p����������G������G���p�������p      B  , ,�������p����������+������+���p�������p      B  , ,���e���p���e���������������p���e���p      B  , ,������l��������������������l������l      B  , ,�������l���������������������l�������l      B  , ,�������l�������������������l�������l      B  , ,�������l����������c������c���l�������l      B  , ,�������l����������G������G���l�������l      B  , ,�������l����������+������+���l�������l      B  , ,���e���l���e���������������l���e���l      B  , ,���E���l���E�����������������l���E���l      B  , ,������������c�������c�������������      B  , ,������e��������������������e������e      B  , ,���E�������E���n�������n�����������E����      B  , ,���)�������)���n�������n�����������)����      B  , ,�������������n�������n���������������      B  , ,���������������n�������n����������������      B  , ,���������������n������n���������������      B  , ,���������������n���c���n���c������������      B  , ,���������������n���G���n���G������������      B  , ,���������������n���+���n���+������������      B  , ,���e�������e���n������n����������e����      B  , ,���E������E����������������������E���      B  , ,���)������)����������������������)���      B  , ,����������������������������������      B  , ,�������������������������������������      B  , ,�����������������������������������      B  , ,������������������c�������c����������      B  , ,������������������G�������G����������      B  , ,������������������+�������+����������      B  , ,���e������e��������������������e���      B  , ,���)���l���)�����������������l���)���l      B  , ,��������������������������������      B  , ,��������������������������������      B  , ,���E�������E���r�������r�����������E����      B  , ,���)�������)���r�������r�����������)����      B  , ,�������������r�������r���������������      B  , ,���������������r�������r����������������      B  , ,���������������r������r���������������      B  , ,���������������r���c���r���c������������      B  , ,���������������r���G���r���G������������      B  , ,���������������r���+���r���+������������      B  , ,���e�������e���r������r����������e����      B  , ,��������������������������������      B  , ,������������������a������a������������      B  , ,������������������E������E������������      B  , ,����������������)������)�����������      B  , ,���c�������c�������������������c����      B  , ,���G�������G���������������������G����      B  , ,���+�������+���������������������+����      B  , ,�����������������������������������      B  , ,��������������������������������������      B  , ,��������������������������������������      B  , ,������������g�������g�������������      B  , ,���m�������m�������������������m����      B  , ,������������������k������k������������      B  , ,�����������������������������������      B  , ,���i�������i�������������������i����      B  , ,������������������g������g������������      B  , ,�����������������������������������      B  , ,���e�������e�������������������e����      B  , ,������������������c������c������������      B  , ,�����������������������������������      B  , ,���a�������a�������������������a����      B  , ,������������������_������_������������      B  , ,���	�������	���������������������	����      B  , ,���]�������]�������������������]����      B  , ,������������������[������[������������      B  , ,�����������������������������������      B  , ,���Y�������Y�������������������Y����      B  , ,������������������W������W������������      B  , ,�����������������������������������      B  , ,���U�������U���������������������U����      B  , ,������i��������������������i������i      B  , ,�������������r�������r���������������      B  , ,���������������r�������r����������������      B  , ,���������������r�������r����������������      B  , ,���������������r���g���r���g������������      B  , ,���������������r���K���r���K������������      B  , ,���������������r���/���r���/������������      B  , ,���i�������i���r������r����������i����      B  , ,���M�������M���r�������r�����������M����      B  , ,������������������e������e������������      B  , ,������������������I������I������������      B  , ,������������������-������-������������      B  , ,���g�������g�������������������g����      B  , ,���K�������K���������������������K����      B  , ,���/�������/���������������������/����      B  , ,�����������������������������������      B  , ,�����������������á�����á������������      B  , ,�����������������ƅ�����ƅ������������      B  , ,���I�������I���r�������r�����������I����      B  , ,���-�������-���r�������r�����������-����      B  , ,��������������������������������������      B  , ,���Q�������Q���������������������Q����      B  , ,������������������O������O������������      B  , ,��������������������������������������      B  , ,���M�������M���������������������M����      B  , ,������������������K������K������������      B  , ,��������������������������������������      B  , ,���I�������I���������������������I����      B  , ,������������������G������G������������      B  , ,��������������������������������������      B  , ,���E�������E���������������������E����      B  , ,������������������C������C������������      B  , ,��������������������������������������      B  , ,���A�������A���������������������A����      B  , ,������������������?������?������������      B  , ,����������������������������������      B  , ,���=�������=���������������������=����      B  , ,��đ������đ������;������;������đ����      B  , ,�����������������Ə�����Ə������������      B  , ,���9�������9���������������������9����      B  , ,������������������k�������k����������      B  , ,��إ�����إ�������O�������O�����إ���      B  , ,��ۉ�����ۉ�������3�������3�����ۉ���      B  , ,���m������m��������������������m���      B  , ,���Q������Q����������������������Q���      B  , ,���5������5����������������������5���      B  , ,����������������������������������      B  , ,�����������������������������������      B  , ,�����������������������������������      B  , ,������������������o�������o����������      B  , ,����������������S�������S���������      B  , ,������������������7�������7����������      B  , ,���q������q��������������������q���      B  , ,���U������U����������������������U���      B  , ,���9������9����������������������9���      B  , ,���5�������5���n�������n�����������5����      B  , ,���5�������5���r�������r�����������5����      B  , ,���5������5����������������������5���      B  , ,���5���p���5�����������������p���5���p      B  , ,���5���l���5�����������������l���5���l      B  , ,���1������1����������������������1���      B  , ,���������������Ϳ������Ϳ���������      B  , ,�����������������У������У����������      B  , ,�����������������Ӈ������Ӈ����������      B  , ,���9�������9���n�������n�����������9����      B  , ,�������������n�������n���������������      B  , ,���������������n������n���������������      B  , ,����������������������������������      B  , ,�����������������������������������      B  , ,�����������������������������������      B  , ,������������������o�������o����������      B  , ,����������������S�������S���������      B  , ,������������������7�������7����������      B  , ,���q������q��������������������q���      B  , ,���U������U����������������������U���      B  , ,���9������9����������������������9���      B  , ,���������������n������n���������������      B  , ,������p��������������������p������p      B  , ,�������p�������������������p�������p      B  , ,�������p�������������������p�������p      B  , ,�������p����������o������o���p�������p      B  , ,������p���������S������S���p������p      B  , ,�������p����������7������7���p�������p      B  , ,���q���p���q���������������p���q���p      B  , ,���U���p���U�����������������p���U���p      B  , ,���9���p���9�����������������p���9���p      B  , ,���������������n���o���n���o������������      B  , ,������l��������������������l������l      B  , ,�������l�������������������l�������l      B  , ,�������l�������������������l�������l      B  , ,�������l����������o������o���l�������l      B  , ,������l���������S������S���l������l      B  , ,�������l����������7������7���l�������l      B  , ,���q���l���q���������������l���q���l      B  , ,���U���l���U�����������������l���U���l      B  , ,���9���l���9�����������������l���9���l      B  , ,�������������n���S���n���S�����������      B  , ,���������������n���7���n���7������������      B  , ,���q�������q���n������n����������q����      B  , ,���U�������U���n�������n�����������U����      B  , ,���m���p���m���������������p���m���p      B  , ,���Q���p���Q�����������������p���Q���p      B  , ,������������������k�������k����������      B  , ,��إ�����إ�������O�������O�����إ���      B  , ,��ۉ�����ۉ�������3�������3�����ۉ���      B  , ,���m������m��������������������m���      B  , ,���Q������Q����������������������Q���      B  , ,��ۉ������ۉ���n���3���n���3������ۉ����      B  , ,���m�������m���n������n����������m����      B  , ,���Q�������Q���n�������n�����������Q����      B  , ,���������������n��У���n��У������������      B  , ,���������������n��Ӈ���n��Ӈ������������      B  , ,�������l���������Ӈ�����Ӈ���l�������l      B  , ,�������l����������k������k���l�������l      B  , ,��إ���l��إ������O������O���l��إ���l      B  , ,��ۉ���l��ۉ������3������3���l��ۉ���l      B  , ,���m���l���m���������������l���m���l      B  , ,���Q���l���Q�����������������l���Q���l      B  , ,���������������n���k���n���k������������      B  , ,���������������Ϳ������Ϳ���������      B  , ,�����������������У������У����������      B  , ,�����������������Ӈ������Ӈ����������      B  , ,��إ������إ���n���O���n���O������إ����      B  , ,������l��������Ϳ�����Ϳ���l������l      B  , ,�������l���������У�����У���l�������l      B  , ,���1���p���1�����������������p���1���p      B  , ,������p��������Ϳ�����Ϳ���p������p      B  , ,�������p���������У�����У���p�������p      B  , ,���1���l���1�����������������l���1���l      B  , ,���1������1����������������������1���      B  , ,���1�������1���n�������n�����������1����      B  , ,�������������n��Ϳ���n��Ϳ�����������      B  , ,�������p���������Ӈ�����Ӈ���p�������p      B  , ,�������p����������k������k���p�������p      B  , ,��إ���p��إ������O������O���p��إ���p      B  , ,��ۉ���p��ۉ������3������3���p��ۉ���p      B  , ,��إ������إ���r���O���r���O������إ����      B  , ,��ۉ������ۉ���r���3���r���3������ۉ����      B  , ,���m�������m���r������r����������m����      B  , ,���Q�������Q���r�������r�����������Q����      B  , ,���1�������1���r�������r�����������1����      B  , ,�������������r��Ϳ���r��Ϳ�����������      B  , ,��ȿ������ȿ������i������i������ȿ����      B  , ,��ˣ������ˣ������M������M������ˣ����      B  , ,��·������·������1������1������·����      B  , ,���k�������k�������������������k����      B  , ,���O�������O���������������������O����      B  , ,���3�������3���������������������3����      B  , ,�����������������������������������      B  , ,�����������������ݥ�����ݥ������������      B  , ,��������������������������������������      B  , ,������������������m������m������������      B  , ,���������������r��У���r��У������������      B  , ,���������������r��Ӈ���r��Ӈ������������      B  , ,���������������r���k���r���k������������      B  , ,��ȍ������ȍ������7������7������ȍ����      B  , ,�����������������ʋ�����ʋ������������      B  , ,���5�������5���������������������5����      B  , ,��̉������̉������3������3������̉����      B  , ,�����������������·�����·������������      B  , ,���1�������1���������������������1����      B  , ,��Ѕ������Ѕ������/������/������Ѕ����      B  , ,�����������������҃�����҃������������      B  , ,���-�������-���������������������-����      B  , ,��ԁ������ԁ������+������+������ԁ����      B  , ,������������������������������������      B  , ,���)�������)���������������������)����      B  , ,���}�������}������'������'�������}����      B  , ,������������������{������{������������      B  , ,���%�������%���������������������%����      B  , ,���y�������y������#������#�������y����      B  , ,������������������w������w������������      B  , ,���!�������!���������������������!����      B  , ,���u�������u�������������������u����      B  , ,������������������s������s������������      B  , ,�����������������������������������      B  , ,���������������r������r���������������      B  , ,����������������Q������Q�����������      B  , ,����������������5������5�����������      B  , ,���o�������o�������������������o����      B  , ,���S�������S���������������������S����      B  , ,���7�������7���������������������7����      B  , ,�����������������������������������      B  , ,��������������������������������������      B  , ,��������������������������������������      B  , ,������������������q������q������������      B  , ,���������������r������r���������������      B  , ,���������������r���o���r���o������������      B  , ,�������������r���S���r���S�����������      B  , ,���������������r���7���r���7������������      B  , ,���q�������q���r������r����������q����      B  , ,���U�������U���r�������r�����������U����      B  , ,���9�������9���r�������r�����������9����      B  , ,�������������r�������r���������������      B  , ,���q�������q�������������������q����      B  , ,������������������o������o������������      B  , ,�����������������������������������      B  , ,���m�������m�������������������m����      B  , ,������������������k������k������������      B  , ,���������������������������������      B  , ,���i�������i�������������������i����      B  , ,����������������g������g�����������      B  , ,���������������������������������      B  , ,���e�������e�������������������e����      B  , ,����������������c������c�����������      B  , ,���������������������������������      B  , ,���a�������a�������������������a����      B  , ,������������������_������_������������      B  , ,���	�������	���������������������	����      B  , ,���]�������]�������������������]����      B  , ,������������������[������[������������      B  , ,�����������������������������������      B  , ,���Y�������Y�������������������Y����      B  , ,������������������W������W������������      B  , ,�����������������������������������      B  , ,  nK���a  nK���  n����  n����a  nK���a      B  , ,  8	���  8	����  8�����  8����  8	���      B  , ,  :����  :�����  ;�����  ;����  :����      B  , ,  =����  =�����  >{����  >{���  =����      B  , ,  @����  @�����  A_����  A_���  @����      B  , ,  C����  C�����  DC����  DC���  C����      B  , ,  F}���  F}����  G'����  G'���  F}���      B  , ,  Ia���  Ia����  J����  J���  Ia���      B  , ,  LE���  LE����  L�����  L����  LE���      B  , ,  O)���  O)����  O�����  O����  O)���      B  , ,  R���  R����  R�����  R����  R���      B  , ,  T����  T�����  U�����  U����  T����      B  , ,  W����  W�����  X����  X���  W����      B  , ,  Z����  Z�����  [c����  [c���  Z����      B  , ,  ]����  ]�����  ^G����  ^G���  ]����      B  , ,  `����  `�����  a+����  a+���  `����      B  , ,  ce���  ce����  d����  d���  ce���      B  , ,  fI���  fI����  f�����  f����  fI���      B  , ,  i-���  i-����  i�����  i����  i-���      B  , ,  l���  l����  l�����  l����  l���      B  , ,  nK����  nK���[  n����[  n�����  nK����      B  , ,  T����d  T����  U����  U����d  T����d      B  , ,  W����d  W����  X���  X���d  W����d      B  , ,  Z����d  Z����  [c���  [c���d  Z����d      B  , ,  ]����d  ]����  ^G���  ^G���d  ]����d      B  , ,  `����d  `����  a+���  a+���d  `����d      B  , ,  ce���d  ce���  d���  d���d  ce���d      B  , ,  fI���d  fI���  f����  f����d  fI���d      B  , ,  i-���d  i-���  i����  i����d  i-���d      B  , ,  l���d  l���  l����  l����d  l���d      B  , ,  nK���  nK����  n�����  n����  nK���      B  , ,  T�����  T����b  U����b  U�����  T�����      B  , ,  W�����  W����b  X���b  X����  W�����      B  , ,  Z�����  Z����b  [c���b  [c����  Z�����      B  , ,  ]�����  ]����b  ^G���b  ^G����  ]�����      B  , ,  `�����  `����b  a+���b  a+����  `�����      B  , ,  ce����  ce���b  d���b  d����  ce����      B  , ,  fI����  fI���b  f����b  f�����  fI����      B  , ,  i-����  i-���b  i����b  i�����  i-����      B  , ,  l����  l���b  l����b  l�����  l����      B  , ,  nK���Y  nK���  n����  n����Y  nK���Y      B  , ,  S����  S���G  T)���G  T)����  S����      B  , ,  Vc����  Vc���G  W���G  W����  Vc����      B  , ,  YG����  YG���G  Y����G  Y�����  YG����      B  , ,  \+����  \+���G  \����G  \�����  \+����      B  , ,  _����  _���G  _����G  _�����  _����      B  , ,  a�����  a����G  b����G  b�����  a�����      B  , ,  d�����  d����G  e����G  e�����  d�����      B  , ,  g�����  g����G  he���G  he����  g�����      B  , ,  j�����  j����G  kI���G  kI����  j�����      B  , ,  nK���  nK����  n�����  n����  nK���      B  , ,  nK����  nK���W  n����W  n�����  nK����      B  , ,  :����d  :����  ;����  ;����d  :����d      B  , ,  =����d  =����  >{���  >{���d  =����d      B  , ,  @����d  @����  A_���  A_���d  @����d      B  , ,  C����d  C����  DC���  DC���d  C����d      B  , ,  F}���d  F}���  G'���  G'���d  F}���d      B  , ,  Ia���d  Ia���  J���  J���d  Ia���d      B  , ,  LE���d  LE���  L����  L����d  LE���d      B  , ,  O)���d  O)���  O����  O����d  O)���d      B  , ,  R���d  R���  R����  R����d  R���d      B  , ,  9{����  9{���G  :%���G  :%����  9{����      B  , ,  <_����  <_���G  =	���G  =	����  <_����      B  , ,  ?C����  ?C���G  ?����G  ?�����  ?C����      B  , ,  B'����  B'���G  B����G  B�����  B'����      B  , ,  E����  E���G  E����G  E�����  E����      B  , ,  G�����  G����G  H����G  H�����  G�����      B  , ,  J�����  J����G  K}���G  K}����  J�����      B  , ,  M�����  M����G  Na���G  Na����  M�����      B  , ,  P�����  P����G  QE���G  QE����  P�����      B  , ,  8	����  8	���b  8����b  8�����  8	����      B  , ,  :�����  :����b  ;����b  ;�����  :�����      B  , ,  =�����  =����b  >{���b  >{����  =�����      B  , ,  @�����  @����b  A_���b  A_����  @�����      B  , ,  C�����  C����b  DC���b  DC����  C�����      B  , ,  F}����  F}���b  G'���b  G'����  F}����      B  , ,  Ia����  Ia���b  J���b  J����  Ia����      B  , ,  LE����  LE���b  L����b  L�����  LE����      B  , ,  O)����  O)���b  O����b  O�����  O)����      B  , ,  R����  R���b  R����b  R�����  R����      B  , ,  8	���d  8	���  8����  8����d  8	���d      B  , ,  @����h  @����  A_���  A_���h  @����h      B  , ,  C����h  C����  DC���  DC���h  C����h      B  , ,  F}���h  F}���  G'���  G'���h  F}���h      B  , ,  Ia���h  Ia���  J���  J���h  Ia���h      B  , ,  LE���h  LE���  L����  L����h  LE���h      B  , ,  O)���h  O)���  O����  O����h  O)���h      B  , ,  R���h  R���  R����  R����h  R���h      B  , ,  @�����  @����f  A_���f  A_����  @�����      B  , ,  8	���  8	����  8�����  8����  8	���      B  , ,  8	����  8	���j  8����j  8�����  8	����      B  , ,  :�����  :����j  ;����j  ;�����  :�����      B  , ,  =�����  =����j  >{���j  >{����  =�����      B  , ,  @�����  @����j  A_���j  A_����  @�����      B  , ,  C�����  C����j  DC���j  DC����  C�����      B  , ,  F}����  F}���j  G'���j  G'����  F}����      B  , ,  Ia����  Ia���j  J���j  J����  Ia����      B  , ,  LE����  LE���j  L����j  L�����  LE����      B  , ,  O)����  O)���j  O����j  O�����  O)����      B  , ,  R����  R���j  R����j  R�����  R����      B  , ,  8	����  8	���f  8����f  8�����  8	����      B  , ,  :����  :�����  ;�����  ;����  :����      B  , ,  =����  =�����  >{����  >{���  =����      B  , ,  @����  @�����  A_����  A_���  @����      B  , ,  C����  C�����  DC����  DC���  C����      B  , ,  F}���  F}����  G'����  G'���  F}���      B  , ,  Ia���  Ia����  J����  J���  Ia���      B  , ,  LE���  LE����  L�����  L����  LE���      B  , ,  O)���  O)����  O�����  O����  O)���      B  , ,  R���  R����  R�����  R����  R���      B  , ,  C�����  C����f  DC���f  DC����  C�����      B  , ,  F}����  F}���f  G'���f  G'����  F}����      B  , ,  Ia����  Ia���f  J���f  J����  Ia����      B  , ,  LE����  LE���f  L����f  L�����  LE����      B  , ,  O)����  O)���f  O����f  O�����  O)����      B  , ,  R����  R���f  R����f  R�����  R����      B  , ,  :�����  :����f  ;����f  ;�����  :�����      B  , ,  =�����  =����f  >{���f  >{����  =�����      B  , ,  8	���h  8	���  8����  8����h  8	���h      B  , ,  :����h  :����  ;����  ;����h  :����h      B  , ,  =����h  =����  >{���  >{���h  =����h      B  , ,  W����  W�����  X����  X���  W����      B  , ,  Z����  Z�����  [c����  [c���  Z����      B  , ,  ]����  ]�����  ^G����  ^G���  ]����      B  , ,  `����  `�����  a+����  a+���  `����      B  , ,  ce���  ce����  d����  d���  ce���      B  , ,  fI���  fI����  f�����  f����  fI���      B  , ,  i-���  i-����  i�����  i����  i-���      B  , ,  l���  l����  l�����  l����  l���      B  , ,  nK����  nK���_  n����_  n�����  nK����      B  , ,  T�����  T����j  U����j  U�����  T�����      B  , ,  W�����  W����j  X���j  X����  W�����      B  , ,  Z�����  Z����j  [c���j  [c����  Z�����      B  , ,  ]�����  ]����j  ^G���j  ^G����  ]�����      B  , ,  `�����  `����j  a+���j  a+����  `�����      B  , ,  ce����  ce���j  d���j  d����  ce����      B  , ,  fI����  fI���j  f����j  f�����  fI����      B  , ,  i-����  i-���j  i����j  i�����  i-����      B  , ,  l����  l���j  l����j  l�����  l����      B  , ,  T����h  T����  U����  U����h  T����h      B  , ,  W����h  W����  X���  X���h  W����h      B  , ,  Z����h  Z����  [c���  [c���h  Z����h      B  , ,  ]����h  ]����  ^G���  ^G���h  ]����h      B  , ,  `����h  `����  a+���  a+���h  `����h      B  , ,  ce���h  ce���  d���  d���h  ce���h      B  , ,  fI���h  fI���  f����  f����h  fI���h      B  , ,  i-���h  i-���  i����  i����h  i-���h      B  , ,  l���h  l���  l����  l����h  l���h      B  , ,  nK���	  nK����  n�����  n����	  nK���	      B  , ,  T�����  T����f  U����f  U�����  T�����      B  , ,  W�����  W����f  X���f  X����  W�����      B  , ,  Z�����  Z����f  [c���f  [c����  Z�����      B  , ,  ]�����  ]����f  ^G���f  ^G����  ]�����      B  , ,  `�����  `����f  a+���f  a+����  `�����      B  , ,  ce����  ce���f  d���f  d����  ce����      B  , ,  fI����  fI���f  f����f  f�����  fI����      B  , ,  i-����  i-���f  i����f  i�����  i-����      B  , ,  l����  l���f  l����f  l�����  l����      B  , ,  nK���]  nK���  n����  n����]  nK���]      B  , ,  T����  T�����  U�����  U����  T����      B  , ,  !���  !����  �����  ����  !���      B  , ,  !���h  !���  ����  ����h  !���h      B  , ,  ���  ����  �����  ����  ���      B  , ,  ���  ����  �����  ����  ���      B  , ,  ����  �����  �����  ����  ����      B  , ,  	����  	�����  
s����  
s���  	����      B  , ,  ����  �����  W����  W���  ����      B  , ,  ����  �����  ;����  ;���  ����      B  , ,  u���  u����  ����  ���  u���      B  , ,  Y���  Y����  ����  ���  Y���      B  , ,  =���  =����  �����  ����  =���      B  , ,  !���  !����  �����  ����  !���      B  , ,  ���  ����  �����  ����  ���      B  , ,   ����   �����  !�����  !����   ����      B  , ,  #����  #�����  $w����  $w���  #����      B  , ,  &����  &�����  '[����  '[���  &����      B  , ,  )����  )�����  *?����  *?���  )����      B  , ,  ,y���  ,y����  -#����  -#���  ,y���      B  , ,  /]���  /]����  0����  0���  /]���      B  , ,  2A���  2A����  2�����  2����  2A���      B  , ,  5%���  5%����  5�����  5����  5%���      B  , ,  !���d  !���  ����  ����d  !���d      B  , ,  !����  !���j  ����j  �����  !����      B  , ,  !����  !���b  ����b  �����  !����      B  , ,  !����  !���f  ����f  �����  !����      B  , ,  &����d  &����  '[���  '[���d  &����d      B  , ,  )����d  )����  *?���  *?���d  )����d      B  , ,  ,y���d  ,y���  -#���  -#���d  ,y���d      B  , ,  /]���d  /]���  0���  0���d  /]���d      B  , ,  2A���d  2A���  2����  2����d  2A���d      B  , ,  5%���d  5%���  5����  5����d  5%���d      B  , ,  ���d  ���  ����  ����d  ���d      B  , ,   ����d   ����  !����  !����d   ����d      B  , ,  ����  ���b  ����b  �����  ����      B  , ,   �����   ����b  !����b  !�����   �����      B  , ,  #�����  #����b  $w���b  $w����  #�����      B  , ,  &�����  &����b  '[���b  '[����  &�����      B  , ,  )�����  )����b  *?���b  *?����  )�����      B  , ,  ,y����  ,y���b  -#���b  -#����  ,y����      B  , ,  /]����  /]���b  0���b  0����  /]����      B  , ,  2A����  2A���b  2����b  2�����  2A����      B  , ,  5%����  5%���b  5����b  5�����  5%����      B  , ,  �����  ����G  =���G  =����  �����      B  , ,  w����  w���G   !���G   !����  w����      B  , ,  "[����  "[���G  #���G  #����  "[����      B  , ,  %?����  %?���G  %����G  %�����  %?����      B  , ,  (#����  (#���G  (����G  (�����  (#����      B  , ,  +����  +���G  +����G  +�����  +����      B  , ,  -�����  -����G  .����G  .�����  -�����      B  , ,  0�����  0����G  1y���G  1y����  0�����      B  , ,  3�����  3����G  4]���G  4]����  3�����      B  , ,  6�����  6����G  7A���G  7A����  6�����      B  , ,  #����d  #����  $w���  $w���d  #����d      B  , ,  =���d  =���  ����  ����d  =���d      B  , ,  ����d  ����  ����  ����d  ����d      B  , ,  	����d  	����  
s���  
s���d  	����d      B  , ,  ����  ���b  ����b  �����  ����      B  , ,  ����  ���b  ����b  �����  ����      B  , ,  �����  ����b  ����b  �����  �����      B  , ,  s����  s���G  ���G  ����  s����      B  , ,  W����  W���G  	���G  	����  W����      B  , ,  ;����  ;���G  ����G  �����  ;����      B  , ,  ����  ���G  ����G  �����  ����      B  , ,  ����  ���G  ����G  �����  ����      B  , ,  �����  ����G  ����G  �����  �����      B  , ,  �����  ����G  u���G  u����  �����      B  , ,  �����  ����G  Y���G  Y����  �����      B  , ,  ���d  ���  ����  ����d  ���d      B  , ,  	�����  	����b  
s���b  
s����  	�����      B  , ,  �����  ����b  W���b  W����  �����      B  , ,  �����  ����b  ;���b  ;����  �����      B  , ,  u����  u���b  ���b  ����  u����      B  , ,  Y����  Y���b  ���b  ����  Y����      B  , ,  =����  =���b  ����b  �����  =����      B  , ,  ����d  ����  W���  W���d  ����d      B  , ,  ����d  ����  ;���  ;���d  ����d      B  , ,  u���d  u���  ���  ���d  u���d      B  , ,  Y���d  Y���  ���  ���d  Y���d      B  , ,  ���d  ���  ����  ����d  ���d      B  , ,  �����  ����G  9���G  9����  �����      B  , ,  ����  ���j  ����j  �����  ����      B  , ,  �����  ����j  ����j  �����  �����      B  , ,  	�����  	����f  
s���f  
s����  	�����      B  , ,  �����  ����f  W���f  W����  �����      B  , ,  �����  ����f  ;���f  ;����  �����      B  , ,  u����  u���f  ���f  ����  u����      B  , ,  	�����  	����j  
s���j  
s����  	�����      B  , ,  �����  ����j  W���j  W����  �����      B  , ,  �����  ����j  ;���j  ;����  �����      B  , ,  u����  u���j  ���j  ����  u����      B  , ,  Y����  Y���j  ���j  ����  Y����      B  , ,  =����  =���j  ����j  �����  =����      B  , ,  ����h  ����  ����  ����h  ����h      B  , ,  	����h  	����  
s���  
s���h  	����h      B  , ,  ����h  ����  W���  W���h  ����h      B  , ,  ����h  ����  ;���  ;���h  ����h      B  , ,  u���h  u���  ���  ���h  u���h      B  , ,  Y���h  Y���  ���  ���h  Y���h      B  , ,  =���h  =���  ����  ����h  =���h      B  , ,  ����  �����  ;����  ;���  ����      B  , ,  u���  u����  ����  ���  u���      B  , ,  ����  ���f  ����f  �����  ����      B  , ,  �����  ����f  ����f  �����  �����      B  , ,  Y���  Y����  ����  ���  Y���      B  , ,  Y����  Y���f  ���f  ����  Y����      B  , ,  =����  =���f  ����f  �����  =����      B  , ,  =���  =����  �����  ����  =���      B  , ,  ����  ���f  ����f  �����  ����      B  , ,  ����  �����  W����  W���  ����      B  , ,  ���h  ���  ����  ����h  ���h      B  , ,  ���h  ���  ����  ����h  ���h      B  , ,  ���  ����  �����  ����  ���      B  , ,  ���  ����  �����  ����  ���      B  , ,  ����  �����  �����  ����  ����      B  , ,  ����  ���j  ����j  �����  ����      B  , ,  	����  	�����  
s����  
s���  	����      B  , ,  ,y����  ,y���j  -#���j  -#����  ,y����      B  , ,  /]����  /]���j  0���j  0����  /]����      B  , ,  2A����  2A���j  2����j  2�����  2A����      B  , ,  5%����  5%���j  5����j  5�����  5%����      B  , ,  2A���h  2A���  2����  2����h  2A���h      B  , ,  5%���h  5%���  5����  5����h  5%���h      B  , ,  5%���  5%����  5�����  5����  5%���      B  , ,  ���  ����  �����  ����  ���      B  , ,   ����   �����  !�����  !����   ����      B  , ,  #����  #�����  $w����  $w���  #����      B  , ,  &����  &�����  '[����  '[���  &����      B  , ,  )����  )�����  *?����  *?���  )����      B  , ,  ,y���  ,y����  -#����  -#���  ,y���      B  , ,  /]���  /]����  0����  0���  /]���      B  , ,  2A���  2A����  2�����  2����  2A���      B  , ,  ���h  ���  ����  ����h  ���h      B  , ,   ����h   ����  !����  !����h   ����h      B  , ,  #����h  #����  $w���  $w���h  #����h      B  , ,  ����  ���f  ����f  �����  ����      B  , ,   �����   ����f  !����f  !�����   �����      B  , ,  #�����  #����f  $w���f  $w����  #�����      B  , ,  &�����  &����f  '[���f  '[����  &�����      B  , ,  )�����  )����f  *?���f  *?����  )�����      B  , ,  ,y����  ,y���f  -#���f  -#����  ,y����      B  , ,  /]����  /]���f  0���f  0����  /]����      B  , ,  2A����  2A���f  2����f  2�����  2A����      B  , ,  5%����  5%���f  5����f  5�����  5%����      B  , ,  &����h  &����  '[���  '[���h  &����h      B  , ,  )����h  )����  *?���  *?���h  )����h      B  , ,  ,y���h  ,y���  -#���  -#���h  ,y���h      B  , ,  /]���h  /]���  0���  0���h  /]���h      B  , ,  ����  ���j  ����j  �����  ����      B  , ,   �����   ����j  !����j  !�����   �����      B  , ,  #�����  #����j  $w���j  $w����  #�����      B  , ,  &�����  &����j  '[���j  '[����  &�����      B  , ,  )�����  )����j  *?���j  *?����  )�����      B  , ,  !���l  !���  ����  ����l  !���l      B  , ,  !���  !����  �����  ����  !���      B  , ,  ���  ����  �����  ����  ���      B  , ,  ���  ����  �����  ����  ���      B  , ,  ����  �����  �����  ����  ����      B  , ,  	����  	�����  
s����  
s���  	����      B  , ,  ����  �����  W����  W���  ����      B  , ,  ����  �����  ;����  ;���  ����      B  , ,  u���  u����  ����  ���  u���      B  , ,  Y���  Y����  ����  ���  Y���      B  , ,  =���  =����  �����  ����  =���      B  , ,  !���  !����  �����  ����  !���      B  , ,  ���  ����  �����  ����  ���      B  , ,   ����   �����  !�����  !����   ����      B  , ,  #����  #�����  $w����  $w���  #����      B  , ,  &����  &�����  '[����  '[���  &����      B  , ,  )����  )�����  *?����  *?���  )����      B  , ,  ,y���  ,y����  -#����  -#���  ,y���      B  , ,  /]���  /]����  0����  0���  /]���      B  , ,  2A���  2A����  2�����  2����  2A���      B  , ,  5%���  5%����  5�����  5����  5%���      B  , ,  !���p  !���  ����  ����p  !���p      B  , ,  !����  !���n  ����n  �����  !����      B  , ,  !����  !���r  ����r  �����  !����      B  , ,   ����l   ����  !����  !����l   ����l      B  , ,  #����l  #����  $w���  $w���l  #����l      B  , ,  5%���l  5%���  5����  5����l  5%���l      B  , ,  ���  ����  �����  ����  ���      B  , ,   ����   �����  !�����  !����   ����      B  , ,  #����  #�����  $w����  $w���  #����      B  , ,  &����  &�����  '[����  '[���  &����      B  , ,  ,y���  ,y����  -#����  -#���  ,y���      B  , ,  /]���  /]����  0����  0���  /]���      B  , ,  2A���  2A����  2�����  2����  2A���      B  , ,  5%���  5%����  5�����  5����  5%���      B  , ,  &����l  &����  '[���  '[���l  &����l      B  , ,  )����l  )����  *?���  *?���l  )����l      B  , ,  ,y���l  ,y���  -#���  -#���l  ,y���l      B  , ,  /]���l  /]���  0���  0���l  /]���l      B  , ,  2A���l  2A���  2����  2����l  2A���l      B  , ,  )����  )�����  *?����  *?���  )����      B  , ,  ���p  ���  ����  ����p  ���p      B  , ,   ����p   ����  !����  !����p   ����p      B  , ,  #����p  #����  $w���  $w���p  #����p      B  , ,  &����p  &����  '[���  '[���p  &����p      B  , ,  )����p  )����  *?���  *?���p  )����p      B  , ,  ,y���p  ,y���  -#���  -#���p  ,y���p      B  , ,  /]���p  /]���  0���  0���p  /]���p      B  , ,  2A���p  2A���  2����  2����p  2A���p      B  , ,  5%���p  5%���  5����  5����p  5%���p      B  , ,  5%����  5%���n  5����n  5�����  5%����      B  , ,  ����  ���n  ����n  �����  ����      B  , ,  ���l  ���  ����  ����l  ���l      B  , ,   �����   ����n  !����n  !�����   �����      B  , ,  #�����  #����n  $w���n  $w����  #�����      B  , ,  &�����  &����n  '[���n  '[����  &�����      B  , ,  )�����  )����n  *?���n  *?����  )�����      B  , ,  ,y����  ,y���n  -#���n  -#����  ,y����      B  , ,  /]����  /]���n  0���n  0����  /]����      B  , ,  2A����  2A���n  2����n  2�����  2A����      B  , ,  ���p  ���  ����  ����p  ���p      B  , ,  ����p  ����  ����  ����p  ����p      B  , ,  	����p  	����  
s���  
s���p  	����p      B  , ,  ����p  ����  W���  W���p  ����p      B  , ,  ����p  ����  ;���  ;���p  ����p      B  , ,  u���p  u���  ���  ���p  u���p      B  , ,  Y���p  Y���  ���  ���p  Y���p      B  , ,  =���p  =���  ����  ����p  =���p      B  , ,  ���  ����  �����  ����  ���      B  , ,  ����  �����  �����  ����  ����      B  , ,  	����  	�����  
s����  
s���  	����      B  , ,  ����  �����  W����  W���  ����      B  , ,  ����  �����  ;����  ;���  ����      B  , ,  u���  u����  ����  ���  u���      B  , ,  Y���  Y����  ����  ���  Y���      B  , ,  =���  =����  �����  ����  =���      B  , ,  =���l  =���  ����  ����l  =���l      B  , ,  ����l  ����  W���  W���l  ����l      B  , ,  �����  ����n  ;���n  ;����  �����      B  , ,  u����  u���n  ���n  ����  u����      B  , ,  Y����  Y���n  ���n  ����  Y����      B  , ,  =����  =���n  ����n  �����  =����      B  , ,  ����l  ����  ;���  ;���l  ����l      B  , ,  u���l  u���  ���  ���l  u���l      B  , ,  Y���l  Y���  ���  ���l  Y���l      B  , ,  ���  ����  �����  ����  ���      B  , ,  ����  ���n  ����n  �����  ����      B  , ,  ����  ���n  ����n  �����  ����      B  , ,  �����  ����n  ����n  �����  �����      B  , ,  	�����  	����n  
s���n  
s����  	�����      B  , ,  �����  ����n  W���n  W����  �����      B  , ,  ���p  ���  ����  ����p  ���p      B  , ,  ���l  ���  ����  ����l  ���l      B  , ,  ���l  ���  ����  ����l  ���l      B  , ,  ����l  ����  ����  ����l  ����l      B  , ,  	����l  	����  
s���  
s���l  	����l      B  , ,  	�����  	����r  
s���r  
s����  	�����      B  , ,  �����  ����r  W���r  W����  �����      B  , ,  �����  ����r  ;���r  ;����  �����      B  , ,  u����  u���r  ���r  ����  u����      B  , ,  Y����  Y���r  ���r  ����  Y����      B  , ,  =����  =���r  ����r  �����  =����      B  , ,  �����  ����  u���  u����  �����      B  , ,  �����  ����  Y���  Y����  �����      B  , ,  �����  ����  9���  9����  �����      B  , ,  s����  s���  ���  ����  s����      B  , ,  W����  W���  	���  	����  W����      B  , ,  ;����  ;���  ����  �����  ;����      B  , ,  ����  ���  ����  �����  ����      B  , ,  ����  ���  ����  �����  ����      B  , ,  �����  ����  ����  �����  �����      B  , ,  ����  ���r  ����r  �����  ����      B  , ,  ����  ���r  ����r  �����  ����      B  , ,  �����  ����r  ����r  �����  �����      B  , ,   U����   U���   ����   �����   U����      B  , ,  �����  ����  S���  S����  �����      B  , ,  �����  ����  ����  �����  �����      B  , ,  Q����  Q���  ����  �����  Q����      B  , ,  �����  ����  O���  O����  �����      B  , ,  �����  ����  ����  �����  �����      B  , ,  M����  M���  ����  �����  M����      B  , ,  	�����  	����  
K���  
K����  	�����      B  , ,  
�����  
����  ����  �����  
�����      B  , ,  I����  I���  ����  �����  I����      B  , ,  �����  ����  G���  G����  �����      B  , ,  �����  ����  ����  �����  �����      B  , ,  E����  E���  ����  �����  E����      B  , ,  �����  ����  C���  C����  �����      B  , ,  �����  ����  ����  �����  �����      B  , ,  A����  A���  ����  �����  A����      B  , ,  �����  ����  ?���  ?����  �����      B  , ,  �����  ����  ����  �����  �����      B  , ,  =����  =���  ����  �����  =����      B  , ,  �����  ����  ;���  ;����  �����      B  , ,  �����  ����  ����  �����  �����      B  , ,  &�����  &����r  '[���r  '[����  &�����      B  , ,  )�����  )����r  *?���r  *?����  )�����      B  , ,  ,y����  ,y���r  -#���r  -#����  ,y����      B  , ,  /]����  /]���r  0���r  0����  /]����      B  , ,  2A����  2A���r  2����r  2�����  2A����      B  , ,  5%����  5%���r  5����r  5�����  5%����      B  , ,  "[����  "[���  #���  #����  "[����      B  , ,  %?����  %?���  %����  %�����  %?����      B  , ,  (#����  (#���  (����  (�����  (#����      B  , ,  +����  +���  +����  +�����  +����      B  , ,  -�����  -����  .����  .�����  -�����      B  , ,  0�����  0����  1y���  1y����  0�����      B  , ,  3�����  3����  4]���  4]����  3�����      B  , ,  6�����  6����  7A���  7A����  6�����      B  , ,  �����  ����  =���  =����  �����      B  , ,  w����  w���   !���   !����  w����      B  , ,  ����  ���r  ����r  �����  ����      B  , ,   �����   ����r  !����r  !�����   �����      B  , ,  #�����  #����r  $w���r  $w����  #�����      B  , ,  9����  9���  ����  �����  9����      B  , ,  �����  ����  7���  7����  �����      B  , ,  �����  ����  ����  �����  �����      B  , ,   5����   5���   ����   �����   5����      B  , ,  !�����  !����  "3���  "3����  !�����      B  , ,  "�����  "����  #����  #�����  "�����      B  , ,  $1����  $1���  $����  $�����  $1����      B  , ,  %�����  %����  &/���  &/����  %�����      B  , ,  &�����  &����  '����  '�����  &�����      B  , ,  (-����  (-���  (����  (�����  (-����      B  , ,  )�����  )����  *+���  *+����  )�����      B  , ,  *�����  *����  +���  +����  *�����      B  , ,  ,)����  ,)���  ,����  ,�����  ,)����      B  , ,  -}����  -}���  .'���  .'����  -}����      B  , ,  .�����  .����  /{���  /{����  .�����      B  , ,  0%����  0%���  0����  0�����  0%����      B  , ,  1y����  1y���  2#���  2#����  1y����      B  , ,  2�����  2����  3w���  3w����  2�����      B  , ,  4!����  4!���  4����  4�����  4!����      B  , ,  5u����  5u���  6���  6����  5u����      B  , ,  6�����  6����  7s���  7s����  6�����      B  , ,  8	���  8	����  8�����  8����  8	���      B  , ,  :����  :�����  ;�����  ;����  :����      B  , ,  =����  =�����  >{����  >{���  =����      B  , ,  @����  @�����  A_����  A_���  @����      B  , ,  C����  C�����  DC����  DC���  C����      B  , ,  F}���  F}����  G'����  G'���  F}���      B  , ,  Ia���  Ia����  J����  J���  Ia���      B  , ,  LE���  LE����  L�����  L����  LE���      B  , ,  O)���  O)����  O�����  O����  O)���      B  , ,  R���  R����  R�����  R����  R���      B  , ,  T����  T�����  U�����  U����  T����      B  , ,  W����  W�����  X����  X���  W����      B  , ,  Z����  Z�����  [c����  [c���  Z����      B  , ,  ]����  ]�����  ^G����  ^G���  ]����      B  , ,  `����  `�����  a+����  a+���  `����      B  , ,  ce���  ce����  d����  d���  ce���      B  , ,  fI���  fI����  f�����  f����  fI���      B  , ,  i-���  i-����  i�����  i����  i-���      B  , ,  l���  l����  l�����  l����  l���      B  , ,  R�����  R����  SW���  SW����  R�����      B  , ,  l���l  l���  l����  l����l  l���l      B  , ,  nK���  nK���  n����  n����  nK���      B  , ,  T����l  T����  U����  U����l  T����l      B  , ,  W����l  W����  X���  X���l  W����l      B  , ,  Z����l  Z����  [c���  [c���l  Z����l      B  , ,  ]����l  ]����  ^G���  ^G���l  ]����l      B  , ,  `����l  `����  a+���  a+���l  `����l      B  , ,  ce���l  ce���  d���  d���l  ce���l      B  , ,  T�����  T����n  U����n  U�����  T�����      B  , ,  W�����  W����n  X���n  X����  W�����      B  , ,  Z�����  Z����n  [c���n  [c����  Z�����      B  , ,  ]�����  ]����n  ^G���n  ^G����  ]�����      B  , ,  `�����  `����n  a+���n  a+����  `�����      B  , ,  ce����  ce���n  d���n  d����  ce����      B  , ,  `����p  `����  a+���  a+���p  `����p      B  , ,  ce���p  ce���  d���  d���p  ce���p      B  , ,  fI���p  fI���  f����  f����p  fI���p      B  , ,  i-���p  i-���  i����  i����p  i-���p      B  , ,  l���p  l���  l����  l����p  l���p      B  , ,  nK���  nK���  n����  n����  nK���      B  , ,  l����  l���n  l����n  l�����  l����      B  , ,  nK���e  nK���  n����  n����e  nK���e      B  , ,  fI���l  fI���  f����  f����l  fI���l      B  , ,  i-���l  i-���  i����  i����l  i-���l      B  , ,  T����  T�����  U�����  U����  T����      B  , ,  W����  W�����  X����  X���  W����      B  , ,  Z����  Z�����  [c����  [c���  Z����      B  , ,  ]����  ]�����  ^G����  ^G���  ]����      B  , ,  `����  `�����  a+����  a+���  `����      B  , ,  ce���  ce����  d����  d���  ce���      B  , ,  fI���  fI����  f�����  f����  fI���      B  , ,  i-���  i-����  i�����  i����  i-���      B  , ,  l���  l����  l�����  l����  l���      B  , ,  fI����  fI���n  f����n  f�����  fI����      B  , ,  i-����  i-���n  i����n  i�����  i-����      B  , ,  T����p  T����  U����  U����p  T����p      B  , ,  W����p  W����  X���  X���p  W����p      B  , ,  Z����p  Z����  [c���  [c���p  Z����p      B  , ,  ]����p  ]����  ^G���  ^G���p  ]����p      B  , ,  nK���  nK���c  n����c  n����  nK���      B  , ,  8	���  8	����  8�����  8����  8	���      B  , ,  :����  :�����  ;�����  ;����  :����      B  , ,  8	���l  8	���  8����  8����l  8	���l      B  , ,  :����l  :����  ;����  ;����l  :����l      B  , ,  =����l  =����  >{���  >{���l  =����l      B  , ,  @����l  @����  A_���  A_���l  @����l      B  , ,  C����l  C����  DC���  DC���l  C����l      B  , ,  F}���l  F}���  G'���  G'���l  F}���l      B  , ,  Ia���l  Ia���  J���  J���l  Ia���l      B  , ,  LE���l  LE���  L����  L����l  LE���l      B  , ,  O)���l  O)���  O����  O����l  O)���l      B  , ,  R���l  R���  R����  R����l  R���l      B  , ,  =����  =�����  >{����  >{���  =����      B  , ,  @����  @�����  A_����  A_���  @����      B  , ,  C����  C�����  DC����  DC���  C����      B  , ,  F}���  F}����  G'����  G'���  F}���      B  , ,  Ia���  Ia����  J����  J���  Ia���      B  , ,  LE���  LE����  L�����  L����  LE���      B  , ,  8	����  8	���n  8����n  8�����  8	����      B  , ,  :�����  :����n  ;����n  ;�����  :�����      B  , ,  =�����  =����n  >{���n  >{����  =�����      B  , ,  @�����  @����n  A_���n  A_����  @�����      B  , ,  C�����  C����n  DC���n  DC����  C�����      B  , ,  F}����  F}���n  G'���n  G'����  F}����      B  , ,  Ia����  Ia���n  J���n  J����  Ia����      B  , ,  8	���p  8	���  8����  8����p  8	���p      B  , ,  :����p  :����  ;����  ;����p  :����p      B  , ,  =����p  =����  >{���  >{���p  =����p      B  , ,  @����p  @����  A_���  A_���p  @����p      B  , ,  C����p  C����  DC���  DC���p  C����p      B  , ,  F}���p  F}���  G'���  G'���p  F}���p      B  , ,  Ia���p  Ia���  J���  J���p  Ia���p      B  , ,  LE���p  LE���  L����  L����p  LE���p      B  , ,  O)���p  O)���  O����  O����p  O)���p      B  , ,  R���p  R���  R����  R����p  R���p      B  , ,  LE����  LE���n  L����n  L�����  LE����      B  , ,  O)����  O)���n  O����n  O�����  O)����      B  , ,  R����  R���n  R����n  R�����  R����      B  , ,  O)���  O)����  O�����  O����  O)���      B  , ,  R���  R����  R�����  R����  R���      B  , ,  O)����  O)���r  O����r  O�����  O)����      B  , ,  R����  R���r  R����r  R�����  R����      B  , ,  J�����  J����  K}���  K}����  J�����      B  , ,  M�����  M����  Na���  Na����  M�����      B  , ,  P�����  P����  QE���  QE����  P�����      B  , ,  E����  E���  E����  E�����  E����      B  , ,  G�����  G����  H����  H�����  G�����      B  , ,  8	����  8	���r  8����r  8�����  8	����      B  , ,  :�����  :����r  ;����r  ;�����  :�����      B  , ,  =�����  =����r  >{���r  >{����  =�����      B  , ,  @�����  @����r  A_���r  A_����  @�����      B  , ,  C�����  C����r  DC���r  DC����  C�����      B  , ,  F}����  F}���r  G'���r  G'����  F}����      B  , ,  Ia����  Ia���r  J���r  J����  Ia����      B  , ,  9{����  9{���  :%���  :%����  9{����      B  , ,  <_����  <_���  =	���  =	����  <_����      B  , ,  ?C����  ?C���  ?����  ?�����  ?C����      B  , ,  B'����  B'���  B����  B�����  B'����      B  , ,  8����  8���  8����  8�����  8����      B  , ,  9q����  9q���  :���  :����  9q����      B  , ,  :�����  :����  ;o���  ;o����  :�����      B  , ,  <����  <���  <����  <�����  <����      B  , ,  =m����  =m���  >���  >����  =m����      B  , ,  >�����  >����  ?k���  ?k����  >�����      B  , ,  @����  @���  @����  @�����  @����      B  , ,  Ai����  Ai���  B���  B����  Ai����      B  , ,  B�����  B����  Cg���  Cg����  B�����      B  , ,  D����  D���  D����  D�����  D����      B  , ,  Ee����  Ee���  F���  F����  Ee����      B  , ,  F�����  F����  Gc���  Gc����  F�����      B  , ,  H����  H���  H����  H�����  H����      B  , ,  Ia����  Ia���  J���  J����  Ia����      B  , ,  J�����  J����  K_���  K_����  J�����      B  , ,  L	����  L	���  L����  L�����  L	����      B  , ,  M]����  M]���  N���  N����  M]����      B  , ,  N�����  N����  O[���  O[����  N�����      B  , ,  P����  P���  P����  P�����  P����      B  , ,  QY����  QY���  R���  R����  QY����      B  , ,  LE����  LE���r  L����r  L�����  LE����      B  , ,  nK���  nK���g  n����g  n����  nK���      B  , ,  \+����  \+���  \����  \�����  \+����      B  , ,  _����  _���  _����  _�����  _����      B  , ,  a�����  a����  b����  b�����  a�����      B  , ,  d�����  d����  e����  e�����  d�����      B  , ,  g�����  g����  he���  he����  g�����      B  , ,  j�����  j����  kI���  kI����  j�����      B  , ,  nK���  nK���  n����  n����  nK���      B  , ,  S����  S���  T)���  T)����  S����      B  , ,  Vc����  Vc���  W���  W����  Vc����      B  , ,  T�����  T����r  U����r  U�����  T�����      B  , ,  W�����  W����r  X���r  X����  W�����      B  , ,  Z�����  Z����r  [c���r  [c����  Z�����      B  , ,  ]�����  ]����r  ^G���r  ^G����  ]�����      B  , ,  `�����  `����r  a+���r  a+����  `�����      B  , ,  ce����  ce���r  d���r  d����  ce����      B  , ,  fI����  fI���r  f����r  f�����  fI����      B  , ,  i-����  i-���r  i����r  i�����  i-����      B  , ,  l����  l���r  l����r  l�����  l����      B  , ,  nK���i  nK���  n����  n����i  nK���i      B  , ,  YG����  YG���  Y����  Y�����  YG����      B  , ,  T����  T���  T����  T�����  T����      B  , ,  UU����  UU���  U����  U�����  UU����      B  , ,  V�����  V����  WS���  WS����  V�����      B  , ,  W�����  W����  X����  X�����  W�����      B  , ,  YQ����  YQ���  Y����  Y�����  YQ����      B  , ,  Z�����  Z����  [O���  [O����  Z�����      B  , ,  [�����  [����  \����  \�����  [�����      B  , ,  ]M����  ]M���  ]����  ]�����  ]M����      B  , ,  ^�����  ^����  _K���  _K����  ^�����      B  , ,  _�����  _����  `����  `�����  _�����      B  , ,  aI����  aI���  a����  a�����  aI����      B  , ,  b�����  b����  cG���  cG����  b�����      B  , ,  c�����  c����  d����  d�����  c�����      B  , ,  eE����  eE���  e����  e�����  eE����      B  , ,  f�����  f����  gC���  gC����  f�����      B  , ,  g�����  g����  h����  h�����  g�����      B  , ,  iA����  iA���  i����  i�����  iA����      B  , ,  j�����  j����  k?���  k?����  j�����      B  , ,  k�����  k����  l����  l�����  k�����      _   ,���G  ���G  �   �  �   �  ���G        _   ,���S���9���S  �����  ��������9���S���9      _   ,���7���9���7  �����  ��������9���7���9      _   ,������9���  �����  ��������9������9      _   ,�������9����  ����q  ����q���9�������9      _   ,�������9����  ����U  ����U���9�������9      _   ,�������9����  ����9  ����9���9�������9      _   ,�������9����  ����  �������9�������9      _   ,�������9����  ����  �������9�������9      _   ,���s���9���s  �����  ��������9���s���9      _   ,���W���9���W  �����  ��������9���W���9      _   ,���;���9���;  �����  ��������9���;���9      _   ,������9���  �����  ��������9������9      _   ,������9���  ����u  ����u���9������9      _   ,�������9����  ����Y  ����Y���9�������9      _   ,�������9����  ����=  ����=���9�������9      _   ,�������9����  ����!  ����!���9�������9      _   ,�����9��  ����  �������9�����9      _   ,���w���9���w  �����  ��������9���w���9      _   ,���[���9���[  �����  ��������9���[���9      _   ,���?���9���?  ���̱  ���̱���9���?���9      _   ,���#���9���#  ���ϕ  ���ϕ���9���#���9      _   ,������9���  ����y  ����y���9������9      _   ,�������9����  ����]  ����]���9�������9      _   ,�������9����  ����A  ����A���9�������9      _   ,��ٳ���9��ٳ  ����%  ����%���9��ٳ���9      _   ,��ܗ���9��ܗ  ����	  ����	���9��ܗ���9      _   ,���{���9���{  �����  ��������9���{���9      _   ,���_���9���_  �����  ��������9���_���9      _   ,���C���9���C  ����  �������9���C���9      _   ,���'���9���'  ����  �������9���'���9      _   ,������9���  ����}  ����}���9������9      _   ,�������9����  ����a  ����a���9�������9      _   ,�������9����  ����E  ����E���9�������9      _   ,������9���  ����)  ����)���9������9      _   ,�������9����  ����  �������9�������9      _   ,������9���  �����  ��������9������9      _   ,���c���9���c  �����  ��������9���c���9      _   ,���G���9���G  �   �  �   ����9���G���9      _   ,  +���9  +  �  �  �  ����9  +���9      _   ,  ���9    �  �  �  ����9  ���9      _   ,  ����9  �  �  	e  �  	e���9  ����9      _   ,  
����9  
�  �  I  �  I���9  
����9      _   ,  ����9  �  �  -  �  -���9  ����9      _   ,  ����9  �  �    �  ���9  ����9      _   ,  ����9  �  �  �  �  ����9  ����9      _   ,  g���9  g  �  �  �  ����9  g���9      _   ,  K���9  K  �  �  �  ����9  K���9      _   ,  /���9  /  �  �  �  ����9  /���9      _   ,  ���9    �   �  �   ����9  ���9      _   ,  !����9  !�  �  #i  �  #i���9  !����9      _   ,  $����9  $�  �  &M  �  &M���9  $����9      _   ,  '����9  '�  �  )1  �  )1���9  '����9      _   ,  *����9  *�  �  ,  �  ,���9  *����9      _   ,  -����9  -�  �  .�  �  .����9  -����9      _   ,  0k���9  0k  �  1�  �  1����9  0k���9      _   ,  3O���9  3O  �  4�  �  4����9  3O���9      _   ,  63���9  63  �  7�  �  7����9  63���9      _   ,  9���9  9  �  :�  �  :����9  9���9      _   ,  ;����9  ;�  �  =m  �  =m���9  ;����9      _   ,  >����9  >�  �  @Q  �  @Q���9  >����9      _   ,  A����9  A�  �  C5  �  C5���9  A����9      _   ,  D����9  D�  �  F  �  F���9  D����9      _   ,  G����9  G�  �  H�  �  H����9  G����9      _   ,  Jo���9  Jo  �  K�  �  K����9  Jo���9      _   ,  MS���9  MS  �  N�  �  N����9  MS���9      _   ,  P7���9  P7  �  Q�  �  Q����9  P7���9      _   ,  S���9  S  �  T�  �  T����9  S���9      _   ,  U����9  U�  �  Wq  �  Wq���9  U����9      _   ,  X����9  X�  �  ZU  �  ZU���9  X����9      _   ,  [����9  [�  �  ]9  �  ]9���9  [����9      _   ,  ^����9  ^�  �  `  �  `���9  ^����9      _   ,  a����9  a�  �  c  �  c���9  a����9      _   ,  ds���9  ds  �  e�  �  e����9  ds���9      _   ,  gW���9  gW  �  h�  �  h����9  gW���9      _   ,  j;���9  j;  �  k�  �  k����9  j;���9      _   ,���G������G����   �����   �������G���      _   ,  �    �  �  	e  �  	e    �        _   ,  
�    
�  �  I  �  I    
�        _   ,  �    �  �  -  �  -    �        _   ,  �    �  �    �      �        _   ,  �    �  �  �  �  �    �        _   ,  g    g  �  �  �  �    g        _   ,  K    K  �  �  �  �    K        _   ,  /    /  �  �  �  �    /        _   ,        �   �  �   �            _   ,  !�    !�  �  #i  �  #i    !�        _   ,  $�    $�  �  &M  �  &M    $�        _   ,  '�    '�  �  )1  �  )1    '�        _   ,  *�    *�  �  ,  �  ,    *�        _   ,  -�    -�  �  .�  �  .�    -�        _   ,  0k    0k  �  1�  �  1�    0k        _   ,  3O    3O  �  4�  �  4�    3O        _   ,  63    63  �  7�  �  7�    63        _   ,  9    9  �  :�  �  :�    9        _   ,  ;�    ;�  �  =m  �  =m    ;�        _   ,  >�    >�  �  @Q  �  @Q    >�        _   ,  A�    A�  �  C5  �  C5    A�        _   ,  D�    D�  �  F  �  F    D�        _   ,  G�    G�  �  H�  �  H�    G�        _   ,  Jo    Jo  �  K�  �  K�    Jo        _   ,  MS    MS  �  N�  �  N�    MS        _   ,  P7    P7  �  Q�  �  Q�    P7        _   ,  S    S  �  T�  �  T�    S        _   ,  U�    U�  �  Wq  �  Wq    U�        _   ,  X�    X�  �  ZU  �  ZU    X�        _   ,  [�    [�  �  ]9  �  ]9    [�        _   ,  ^�    ^�  �  `  �  `    ^�        _   ,  a�    a�  �  c  �  c    a�        _   ,  ds    ds  �  e�  �  e�    ds        _   ,  gW    gW  �  h�  �  h�    gW        _   ,  j;    j;  �  k�  �  k�    j;        _   ,  +    +  �  �  �  �    +        _   ,        �  �  �  �            _   ,����  ����  ����q  ����q  ����        _   ,����  ����  ����U  ����U  ����        _   ,����  ����  ����9  ����9  ����        _   ,����  ����  ����  ����  ����        _   ,����  ����  ����  ����  ����        _   ,���s  ���s  �����  �����  ���s        _   ,���W  ���W  �����  �����  ���W        _   ,���;  ���;  �����  �����  ���;        _   ,���  ���  �����  �����  ���        _   ,���  ���  ����u  ����u  ���        _   ,����  ����  ����Y  ����Y  ����        _   ,����  ����  ����=  ����=  ����        _   ,����  ����  ����!  ����!  ����        _   ,��  ��  ����  ����  ��        _   ,���w  ���w  �����  �����  ���w        _   ,���[  ���[  �����  �����  ���[        _   ,���?  ���?  ���̱  ���̱  ���?        _   ,���#  ���#  ���ϕ  ���ϕ  ���#        _   ,���  ���  ����y  ����y  ���        _   ,����  ����  ����]  ����]  ����        _   ,����  ����  ����A  ����A  ����        _   ,��ٳ  ��ٳ  ����%  ����%  ��ٳ        _   ,��ܗ  ��ܗ  ����	  ����	  ��ܗ        _   ,���{  ���{  �����  �����  ���{        _   ,���_  ���_  �����  �����  ���_        _   ,���C  ���C  ����  ����  ���C        _   ,���'  ���'  ����  ����  ���'        _   ,���  ���  ����}  ����}  ���        _   ,����  ����  ����a  ����a  ����        _   ,����  ����  ����E  ����E  ����        _   ,���  ���  ����)  ����)  ���        _   ,����  ����  ����  ����  ����        _   ,���  ���  �����  �����  ���        _   ,���c  ���c  �����  �����  ���c        _   ,���S  ���S  �����  �����  ���S        _   ,���7  ���7  �����  �����  ���7        _   ,���  ���  �����  �����  ���        _   ,���7������7����������������������7���      _   ,����������������������������������      _   ,������������������q�������q����������      _   ,������������������U�������U����������      _   ,������������������9�������9����������      _   ,�����������������������������������      _   ,�����������������������������������      _   ,���s������s����������������������s���      _   ,���W������W����������������������W���      _   ,���;������;����������������������;���      _   ,����������������������������������      _   ,����������������u�������u���������      _   ,������������������Y�������Y����������      _   ,������������������=�������=����������      _   ,������������������!�������!����������      _   ,�����������������������������      _   ,���w������w����������������������w���      _   ,���[������[����������������������[���      _   ,���?������?������̱������̱������?���      _   ,���#������#������ϕ������ϕ������#���      _   ,����������������y�������y���������      _   ,������������������]�������]����������      _   ,������������������A�������A����������      _   ,��ٳ�����ٳ�������%�������%�����ٳ���      _   ,��ܗ�����ܗ�������	�������	�����ܗ���      _   ,���{������{����������������������{���      _   ,���_������_����������������������_���      _   ,���C������C��������������������C���      _   ,���'������'��������������������'���      _   ,����������������}�������}���������      _   ,������������������a�������a����������      _   ,������������������E�������E����������      _   ,����������������)�������)���������      _   ,�����������������������������������      _   ,����������������������������������      _   ,���c������c����������������������c���      _   ,���S������S����������������������S���      _   ,  +���  +����  �����  ����  +���      _   ,  ���  ����  �����  ����  ���      _   ,  ����  �����  	e����  	e���  ����      _   ,  
����  
�����  I����  I���  
����      _   ,  ����  �����  -����  -���  ����      _   ,  ����  �����  ����  ���  ����      _   ,  ����  �����  �����  ����  ����      _   ,  g���  g����  �����  ����  g���      _   ,  K���  K����  �����  ����  K���      _   ,  /���  /����  �����  ����  /���      _   ,  ���  ����   �����   ����  ���      _   ,  !����  !�����  #i����  #i���  !����      _   ,  $����  $�����  &M����  &M���  $����      _   ,  '����  '�����  )1����  )1���  '����      _   ,  *����  *�����  ,����  ,���  *����      _   ,  -����  -�����  .�����  .����  -����      _   ,  0k���  0k����  1�����  1����  0k���      _   ,  3O���  3O����  4�����  4����  3O���      _   ,  63���  63����  7�����  7����  63���      _   ,  9���  9����  :�����  :����  9���      _   ,  ;����  ;�����  =m����  =m���  ;����      _   ,  >����  >�����  @Q����  @Q���  >����      _   ,  A����  A�����  C5����  C5���  A����      _   ,  D����  D�����  F����  F���  D����      _   ,  G����  G�����  H�����  H����  G����      _   ,  Jo���  Jo����  K�����  K����  Jo���      _   ,  MS���  MS����  N�����  N����  MS���      _   ,  P7���  P7����  Q�����  Q����  P7���      _   ,  S���  S����  T�����  T����  S���      _   ,  U����  U�����  Wq����  Wq���  U����      _   ,  X����  X�����  ZU����  ZU���  X����      _   ,  [����  [�����  ]9����  ]9���  [����      _   ,  ^����  ^�����  `����  `���  ^����      _   ,  a����  a�����  c����  c���  a����      _   ,  ds���  ds����  e�����  e����  ds���      _   ,  gW���  gW����  h�����  h����  gW���      _   ,  j;���  j;����  k�����  k����  j;���      C   ,���  q���    n�    n�  q���  q      C   ,���������  q����  q�������������      C   ,���  s���     �     �  s���  s      C   ,���   ����  c   �  c   �   ����   �      C   ,�������������G   ����G   ������������      C   ,�������������   ����   ������������      C   ,  nK���  nK  q  n�  q  n����  nK���      C   ,�������������  n����  n������������      C   ,  6  s  6    7�    7�  s  6  s      C   ,        �  �  �  �            C   ,        �  �  �  �            C   ,  �    �  �  �  �  �    �        C   ,  	�    	�  �  
s  �  
s    	�        C   ,  �    �  �  W  �  W    �        C   ,  �    �  �  ;  �  ;    �        C   ,  u    u  �    �      u        C   ,  Y    Y  �    �      Y        C   ,  =    =  �  �  �  �    =        C   ,  !    !  �  �  �  �    !        C   ,        �  �  �  �            C   ,   �     �  �  !�  �  !�     �        C   ,  #�    #�  �  $w  �  $w    #�        C   ,  &�    &�  �  '[  �  '[    &�        C   ,  )�    )�  �  *?  �  *?    )�        C   ,  ,y    ,y  �  -#  �  -#    ,y        C   ,  /]    /]  �  0  �  0    /]        C   ,  2A    2A  �  2�  �  2�    2A        C   ,  5%    5%  �  5�  �  5�    5%        C   ,  8	    8	  �  8�  �  8�    8	        C   ,  :�    :�  �  ;�  �  ;�    :�        C   ,  =�    =�  �  >{  �  >{    =�        C   ,  @�    @�  �  A_  �  A_    @�        C   ,  C�    C�  �  DC  �  DC    C�        C   ,  F}    F}  �  G'  �  G'    F}        C   ,  Ia    Ia  �  J  �  J    Ia        C   ,  LE    LE  �  L�  �  L�    LE        C   ,  O)    O)  �  O�  �  O�    O)        C   ,  R    R  �  R�  �  R�    R        C   ,  T�    T�  �  U�  �  U�    T�        C   ,  W�    W�  �  X  �  X    W�        C   ,  Z�    Z�  �  [c  �  [c    Z�        C   ,  ]�    ]�  �  ^G  �  ^G    ]�        C   ,  `�    `�  �  a+  �  a+    `�        C   ,  ce    ce  �  d  �  d    ce        C   ,  fI    fI  �  f�  �  f�    fI        C   ,  i-    i-  �  i�  �  i�    i-        C   ,  l    l  �  l�  �  l�    l        C   ,  6   �  6  c  7�  c  7�   �  6   �      C   ,  A�  s  A�    C]    C]  s  A�  s      C   ,  D  s  D    FA    FA  s  D  s      C   ,  Gc  s  Gc    I%    I%  s  Gc  s      C   ,  JG  s  JG    L	    L	  s  JG  s      C   ,  M+  s  M+    N�    N�  s  M+  s      C   ,  P  s  P    Q�    Q�  s  P  s      C   ,  R�  s  R�    T�    T�  s  R�  s      C   ,  U�  s  U�    W�    W�  s  U�  s      C   ,  X�  s  X�    Z}    Z}  s  X�  s      C   ,  [�  s  [�    ]a    ]a  s  [�  s      C   ,  ^�  s  ^�    `E    `E  s  ^�  s      C   ,  ag  s  ag    c)    c)  s  ag  s      C   ,  dK  s  dK    f    f  s  dK  s      C   ,  g/  s  g/    h�    h�  s  g/  s      C   ,  j  s  j    k�    k�  s  j  s      C   ,  8�  s  8�    :�    :�  s  8�  s      C   ,  ;�  s  ;�    =�    =�  s  ;�  s      C   ,  >�  s  >�    @y    @y  s  >�  s      C   ,  !�  s  !�    #�    #�  s  !�  s      C   ,  $�  s  $�    &u    &u  s  $�  s      C   ,  '�  s  '�    )Y    )Y  s  '�  s      C   ,  *{  s  *{    ,=    ,=  s  *{  s      C   ,  -_  s  -_    /!    /!  s  -_  s      C   ,  0C  s  0C    2    2  s  0C  s      C   ,  3'  s  3'    4�    4�  s  3'  s      C   ,  w  s  w    9    9  s  w  s      C   ,  [  s  [          s  [  s      C   ,  ?  s  ?          s  ?  s      C   ,  #  s  #    �    �  s  #  s      C   ,    s      �    �  s    s      C   ,    s      �    �  s    s      C   ,  �  s  �     �     �  s  �  s      C   ,  �  s  �    �    �  s  �  s      C   ,  �  s  �    	�    	�  s  �  s      C   ,  
�  s  
�    q    q  s  
�  s      C   ,  �  s  �    U    U  s  �  s      C   ,  w   �  w  c  9  c  9   �  w   �      C   ,  [   �  [  c    c     �  [   �      C   ,  ?   �  ?  c    c     �  ?   �      C   ,  #   �  #  c  �  c  �   �  #   �      C   ,     �    c  �  c  �   �     �      C   ,  �   �  �  c   �  c   �   �  �   �      C   ,  !�   �  !�  c  #�  c  #�   �  !�   �      C   ,  $�   �  $�  c  &u  c  &u   �  $�   �      C   ,  '�   �  '�  c  )Y  c  )Y   �  '�   �      C   ,  *{   �  *{  c  ,=  c  ,=   �  *{   �      C   ,  -_   �  -_  c  /!  c  /!   �  -_   �      C   ,  0C   �  0C  c  2  c  2   �  0C   �      C   ,  3'   �  3'  c  4�  c  4�   �  3'   �      C   ,     �    c  �  c  �   �     �      C   ,  �   �  �  c  �  c  �   �  �   �      C   ,  �   �  �  c  	�  c  	�   �  �   �      C   ,  
�   �  
�  c  q  c  q   �  
�   �      C   ,  �   �  �  c  U  c  U   �  �   �      C   ,  D   �  D  c  FA  c  FA   �  D   �      C   ,  Gc   �  Gc  c  I%  c  I%   �  Gc   �      C   ,  JG   �  JG  c  L	  c  L	   �  JG   �      C   ,  M+   �  M+  c  N�  c  N�   �  M+   �      C   ,  P   �  P  c  Q�  c  Q�   �  P   �      C   ,  R�   �  R�  c  T�  c  T�   �  R�   �      C   ,  U�   �  U�  c  W�  c  W�   �  U�   �      C   ,  X�   �  X�  c  Z}  c  Z}   �  X�   �      C   ,  [�   �  [�  c  ]a  c  ]a   �  [�   �      C   ,  ^�   �  ^�  c  `E  c  `E   �  ^�   �      C   ,  ag   �  ag  c  c)  c  c)   �  ag   �      C   ,  dK   �  dK  c  f  c  f   �  dK   �      C   ,  g/   �  g/  c  h�  c  h�   �  g/   �      C   ,  j   �  j  c  k�  c  k�   �  j   �      C   ,  8�   �  8�  c  :�  c  :�   �  8�   �      C   ,  ;�   �  ;�  c  =�  c  =�   �  ;�   �      C   ,  >�   �  >�  c  @y  c  @y   �  >�   �      C   ,  A�   �  A�  c  C]  c  C]   �  A�   �      C   ,���3  s���3  ����  ����  s���3  s      C   ,���E  ���E  �����  �����  ���E        C   ,���3   ����3  c����  c����   ����3   �      C   ,���)  ���)  �����  �����  ���)        C   ,���  ���  �����  �����  ���        C   ,����  ����  �����  �����  ����        C   ,����  ����  ����  ����  ����        C   ,����  ����  ����c  ����c  ����        C   ,����  ����  ����G  ����G  ����        C   ,����  ����  ����+  ����+  ����        C   ,���e  ���e  ����  ����  ���e        C   ,���I  ���I  �����  �����  ���I        C   ,���-  ���-  �����  �����  ���-        C   ,���  ���  �����  �����  ���        C   ,����  ����  �����  �����  ����        C   ,����  ����  �����  �����  ����        C   ,����  ����  ����g  ����g  ����        C   ,����  ����  ����K  ����K  ����        C   ,����  ����  ����/  ����/  ����        C   ,���i  ���i  ����  ����  ���i        C   ,���M  ���M  �����  �����  ���M        C   ,���1  ���1  �����  �����  ���1        C   ,���  ���  ���Ϳ  ���Ϳ  ���        C   ,����  ����  ���У  ���У  ����        C   ,����  ����  ���Ӈ  ���Ӈ  ����        C   ,����  ����  ����k  ����k  ����        C   ,��إ  ��إ  ����O  ����O  ��إ        C   ,��ۉ  ��ۉ  ����3  ����3  ��ۉ        C   ,���m  ���m  ����  ����  ���m        C   ,���Q  ���Q  �����  �����  ���Q        C   ,���5  ���5  �����  �����  ���5        C   ,���  ���  �����  �����  ���        C   ,����  ����  ����  ����  ����        C   ,����  ����  ����  ����  ����        C   ,����  ����  ����o  ����o  ����        C   ,���  ���  ����S  ����S  ���        C   ,����  ����  ����7  ����7  ����        C   ,���q  ���q  ����  ����  ���q        C   ,���U  ���U  �����  �����  ���U        C   ,���9  ���9  �����  �����  ���9        C   ,����  s����  ��Յ  ��Յ  s����  s      C   ,��֧  s��֧  ���i  ���i  s��֧  s      C   ,��ً  s��ً  ���M  ���M  s��ً  s      C   ,���o  s���o  ���1  ���1  s���o  s      C   ,���S  s���S  ���  ���  s���S  s      C   ,���7  s���7  ����  ����  s���7  s      C   ,���  s���  ����  ����  s���  s      C   ,����  s����  ����  ����  s����  s      C   ,����  s����  ���  ���  s����  s      C   ,����  s����  ���  ���  s����  s      C   ,���  s���  ���m  ���m  s���  s      C   ,���  s���  ���Q  ���Q  s���  s      C   ,���s  s���s  ���5  ���5  s���s  s      C   ,���W  s���W  ���  ���  s���W  s      C   ,���;  s���;  ����  ����  s���;  s      C   ,���  s���  ����  ����  s���  s      C   ,����  s����  ��Ͻ  ��Ͻ  s����  s      C   ,����  s����  ��ҡ  ��ҡ  s����  s      C   ,����  s����  ����  ����  s����  s      C   ,����  s����  ���e  ���e  s����  s      C   ,����  s����  ���I  ���I  s����  s      C   ,���k  s���k  ���-  ���-  s���k  s      C   ,���O  s���O  ���  ���  s���O  s      C   ,����  s����  ���E  ���E  s����  s      C   ,���g  s���g  ���)  ���)  s���g  s      C   ,���K  s���K  ���  ���  s���K  s      C   ,���/  s���/  ����  ����  s���/  s      C   ,���  s���  ����  ����  s���  s      C   ,����  s����  ����  ����  s����  s      C   ,����  s����  ����  ����  s����  s      C   ,���+  s���+  ����  ����  s���+  s      C   ,���  s���  ����  ����  s���  s      C   ,����  s����  ����  ����  s����  s      C   ,����  s����  ����  ����  s����  s      C   ,����  s����  ���}  ���}  s����  s      C   ,����  s����  ���a  ���a  s����  s      C   ,���g   ����g  c���)  c���)   ����g   �      C   ,���K   ����K  c���  c���   ����K   �      C   ,���/   ����/  c����  c����   ����/   �      C   ,���   ����  c����  c����   ����   �      C   ,����   �����  c����  c����   �����   �      C   ,����   �����  c����  c����   �����   �      C   ,����   �����  c����  c����   �����   �      C   ,����   �����  c���e  c���e   �����   �      C   ,����   �����  c���I  c���I   �����   �      C   ,���k   ����k  c���-  c���-   ����k   �      C   ,���O   ����O  c���  c���   ����O   �      C   ,���+   ����+  c����  c����   ����+   �      C   ,���   ����  c����  c����   ����   �      C   ,����   �����  c����  c����   �����   �      C   ,����   �����  c����  c����   �����   �      C   ,����   �����  c���}  c���}   �����   �      C   ,����   �����  c���a  c���a   �����   �      C   ,����   �����  c���E  c���E   �����   �      C   ,���o   ����o  c���1  c���1   ����o   �      C   ,���S   ����S  c���  c���   ����S   �      C   ,���7   ����7  c����  c����   ����7   �      C   ,���   ����  c����  c����   ����   �      C   ,����   �����  c����  c����   �����   �      C   ,����   �����  c���  c���   �����   �      C   ,����   �����  c���  c���   �����   �      C   ,���   ����  c���m  c���m   ����   �      C   ,���   ����  c���Q  c���Q   ����   �      C   ,���s   ����s  c���5  c���5   ����s   �      C   ,���W   ����W  c���  c���   ����W   �      C   ,���;   ����;  c����  c����   ����;   �      C   ,���   ����  c����  c����   ����   �      C   ,����   �����  c��Ͻ  c��Ͻ   �����   �      C   ,����   �����  c��ҡ  c��ҡ   �����   �      C   ,����   �����  c��Յ  c��Յ   �����   �      C   ,��֧   ���֧  c���i  c���i   ���֧   �      C   ,��ً   ���ً  c���M  c���M   ���ً   �      C   ,���3�������3���G�������G�����������3����      C   ,���E���7���E�������������������7���E���7      C   ,���)���7���)�������������������7���)���7      C   ,������7����������������������7������7      C   ,�������7�����������������������7�������7      C   ,�������7���������������������7�������7      C   ,�������7�����������c�������c���7�������7      C   ,�������7�����������G�������G���7�������7      C   ,�������7�����������+�������+���7�������7      C   ,���e���7���e�����������������7���e���7      C   ,���I���7���I�������������������7���I���7      C   ,���-���7���-�������������������7���-���7      C   ,������7����������������������7������7      C   ,�������7�����������������������7�������7      C   ,�������7�����������������������7�������7      C   ,�������7�����������g�������g���7�������7      C   ,�������7�����������K�������K���7�������7      C   ,�������7�����������/�������/���7�������7      C   ,���i���7���i�����������������7���i���7      C   ,���M���7���M�������������������7���M���7      C   ,���1���7���1�������������������7���1���7      C   ,������7���������Ϳ������Ϳ���7������7      C   ,�������7����������У������У���7�������7      C   ,�������7����������Ӈ������Ӈ���7�������7      C   ,�������7�����������k�������k���7�������7      C   ,��إ���7��إ�������O�������O���7��إ���7      C   ,��ۉ���7��ۉ�������3�������3���7��ۉ���7      C   ,���m���7���m�����������������7���m���7      C   ,���Q���7���Q�������������������7���Q���7      C   ,���5���7���5�������������������7���5���7      C   ,������7����������������������7������7      C   ,�������7���������������������7�������7      C   ,�������7���������������������7�������7      C   ,�������7�����������o�������o���7�������7      C   ,������7����������S�������S���7������7      C   ,�������7�����������7�������7���7�������7      C   ,���q���7���q�����������������7���q���7      C   ,���U���7���U�������������������7���U���7      C   ,���9���7���9�������������������7���9���7      C   ,���3�������3���������������������3����      C   ,���������������G��Յ���G��Յ������������      C   ,��֧������֧���G���i���G���i������֧����      C   ,��ً������ً���G���M���G���M������ً����      C   ,���o�������o���G���1���G���1�������o����      C   ,���S�������S���G������G����������S����      C   ,���7�������7���G�������G�����������7����      C   ,�������������G�������G���������������      C   ,���������������G�������G����������������      C   ,���������������G������G���������������      C   ,���������������G������G���������������      C   ,�������������G���m���G���m�����������      C   ,�������������G���Q���G���Q�����������      C   ,���s�������s���G���5���G���5�������s����      C   ,���W�������W���G������G����������W����      C   ,���;�������;���G�������G�����������;����      C   ,�������������G�������G���������������      C   ,���������������G��Ͻ���G��Ͻ������������      C   ,���������������G��ҡ���G��ҡ������������      C   ,���������������G���}���G���}������������      C   ,���������������G���a���G���a������������      C   ,���������������G���E���G���E������������      C   ,���g�������g���G���)���G���)�������g����      C   ,���K�������K���G������G����������K����      C   ,���+�������+���G�������G�����������+����      C   ,���/�������/���G�������G�����������/����      C   ,�������������G�������G���������������      C   ,���������������G�������G����������������      C   ,���������������G�������G����������������      C   ,���������������G�������G����������������      C   ,���������������G���e���G���e������������      C   ,���������������G���I���G���I������������      C   ,���k�������k���G���-���G���-�������k����      C   ,���O�������O���G������G����������O����      C   ,�������������G�������G���������������      C   ,���������������G�������G����������������      C   ,���������������G�������G����������������      C   ,������������������}������}������������      C   ,������������������a������a������������      C   ,������������������E������E������������      C   ,���g�������g������)������)�������g����      C   ,���K�������K�������������������K����      C   ,���/�������/���������������������/����      C   ,�����������������������������������      C   ,��������������������������������������      C   ,��������������������������������������      C   ,��������������������������������������      C   ,������������������e������e������������      C   ,������������������I������I������������      C   ,���k�������k������-������-�������k����      C   ,���O�������O�������������������O����      C   ,���+�������+���������������������+����      C   ,�����������������������������������      C   ,��������������������������������������      C   ,��������������������������������������      C   ,�����������������Յ�����Յ������������      C   ,��֧������֧������i������i������֧����      C   ,��ً������ً������M������M������ً����      C   ,���o�������o������1������1�������o����      C   ,���S�������S�������������������S����      C   ,���7�������7���������������������7����      C   ,�����������������������������������      C   ,��������������������������������������      C   ,������������������������������������      C   ,������������������������������������      C   ,����������������m������m�����������      C   ,����������������Q������Q�����������      C   ,���s�������s������5������5�������s����      C   ,���W�������W�������������������W����      C   ,���;�������;���������������������;����      C   ,�����������������������������������      C   ,�����������������Ͻ�����Ͻ������������      C   ,�����������������ҡ�����ҡ������������      C   ,  	����7  	�����  
s����  
s���7  	����7      C   ,  ����7  �����  W����  W���7  ����7      C   ,  ����7  �����  ;����  ;���7  ����7      C   ,  u���7  u����  ����  ���7  u���7      C   ,  Y���7  Y����  ����  ���7  Y���7      C   ,  =���7  =����  �����  ����7  =���7      C   ,  !���7  !����  �����  ����7  !���7      C   ,  ���7  ����  �����  ����7  ���7      C   ,   ����7   �����  !�����  !����7   ����7      C   ,  #����7  #�����  $w����  $w���7  #����7      C   ,  &����7  &�����  '[����  '[���7  &����7      C   ,  )����7  )�����  *?����  *?���7  )����7      C   ,  ,y���7  ,y����  -#����  -#���7  ,y���7      C   ,  /]���7  /]����  0����  0���7  /]���7      C   ,  2A���7  2A����  2�����  2����7  2A���7      C   ,  5%���7  5%����  5�����  5����7  5%���7      C   ,  8	���7  8	����  8�����  8����7  8	���7      C   ,  :����7  :�����  ;�����  ;����7  :����7      C   ,  =����7  =�����  >{����  >{���7  =����7      C   ,  @����7  @�����  A_����  A_���7  @����7      C   ,  C����7  C�����  DC����  DC���7  C����7      C   ,  F}���7  F}����  G'����  G'���7  F}���7      C   ,  Ia���7  Ia����  J����  J���7  Ia���7      C   ,  LE���7  LE����  L�����  L����7  LE���7      C   ,  O)���7  O)����  O�����  O����7  O)���7      C   ,  R���7  R����  R�����  R����7  R���7      C   ,  T����7  T�����  U�����  U����7  T����7      C   ,  W����7  W�����  X����  X���7  W����7      C   ,  Z����7  Z�����  [c����  [c���7  Z����7      C   ,  ]����7  ]�����  ^G����  ^G���7  ]����7      C   ,  `����7  `�����  a+����  a+���7  `����7      C   ,  ce���7  ce����  d����  d���7  ce���7      C   ,  fI���7  fI����  f�����  f����7  fI���7      C   ,  i-���7  i-����  i�����  i����7  i-���7      C   ,  l���7  l����  l�����  l����7  l���7      C   ,  6����  6���G  7����G  7�����  6����      C   ,  ���7  ����  �����  ����7  ���7      C   ,  6����  6���  7����  7�����  6����      C   ,  ���7  ����  �����  ����7  ���7      C   ,  ����7  �����  �����  ����7  ����7      C   ,  D����  D���G  FA���G  FA����  D����      C   ,  Gc����  Gc���G  I%���G  I%����  Gc����      C   ,  JG����  JG���G  L	���G  L	����  JG����      C   ,  M+����  M+���G  N����G  N�����  M+����      C   ,  P����  P���G  Q����G  Q�����  P����      C   ,  R�����  R����G  T����G  T�����  R�����      C   ,  U�����  U����G  W����G  W�����  U�����      C   ,  X�����  X����G  Z}���G  Z}����  X�����      C   ,  [�����  [����G  ]a���G  ]a����  [�����      C   ,  ^�����  ^����G  `E���G  `E����  ^�����      C   ,  ag����  ag���G  c)���G  c)����  ag����      C   ,  dK����  dK���G  f���G  f����  dK����      C   ,  g/����  g/���G  h����G  h�����  g/����      C   ,  j����  j���G  k����G  k�����  j����      C   ,  8�����  8����G  :����G  :�����  8�����      C   ,  ;�����  ;����G  =����G  =�����  ;�����      C   ,  >�����  >����G  @y���G  @y����  >�����      C   ,  A�����  A����G  C]���G  C]����  A�����      C   ,  ?����  ?���G  ���G  ����  ?����      C   ,  #����  #���G  ����G  �����  #����      C   ,  ����  ���G  ����G  �����  ����      C   ,  �����  ����G   ����G   �����  �����      C   ,  !�����  !����G  #����G  #�����  !�����      C   ,  $�����  $����G  &u���G  &u����  $�����      C   ,  '�����  '����G  )Y���G  )Y����  '�����      C   ,  *{����  *{���G  ,=���G  ,=����  *{����      C   ,  -_����  -_���G  /!���G  /!����  -_����      C   ,  0C����  0C���G  2���G  2����  0C����      C   ,  3'����  3'���G  4����G  4�����  3'����      C   ,  �����  ����G  ����G  �����  �����      C   ,  �����  ����G  	����G  	�����  �����      C   ,  ����  ���G  ����G  �����  ����      C   ,  
�����  
����G  q���G  q����  
�����      C   ,  �����  ����G  U���G  U����  �����      C   ,  w����  w���G  9���G  9����  w����      C   ,  [����  [���G  ���G  ����  [����      C   ,  
�����  
����  q���  q����  
�����      C   ,  �����  ����  U���  U����  �����      C   ,  w����  w���  9���  9����  w����      C   ,  [����  [���  ���  ����  [����      C   ,  ?����  ?���  ���  ����  ?����      C   ,  #����  #���  ����  �����  #����      C   ,  ����  ���  ����  �����  ����      C   ,  �����  ����   ����   �����  �����      C   ,  !�����  !����  #����  #�����  !�����      C   ,  $�����  $����  &u���  &u����  $�����      C   ,  '�����  '����  )Y���  )Y����  '�����      C   ,  *{����  *{���  ,=���  ,=����  *{����      C   ,  -_����  -_���  /!���  /!����  -_����      C   ,  0C����  0C���  2���  2����  0C����      C   ,  3'����  3'���  4����  4�����  3'����      C   ,  ����  ���  ����  �����  ����      C   ,  �����  ����  ����  �����  �����      C   ,  �����  ����  	����  	�����  �����      C   ,  >�����  >����  @y���  @y����  >�����      C   ,  A�����  A����  C]���  C]����  A�����      C   ,  D����  D���  FA���  FA����  D����      C   ,  Gc����  Gc���  I%���  I%����  Gc����      C   ,  JG����  JG���  L	���  L	����  JG����      C   ,  M+����  M+���  N����  N�����  M+����      C   ,  P����  P���  Q����  Q�����  P����      C   ,  R�����  R����  T����  T�����  R�����      C   ,  U�����  U����  W����  W�����  U�����      C   ,  X�����  X����  Z}���  Z}����  X�����      C   ,  [�����  [����  ]a���  ]a����  [�����      C   ,  ^�����  ^����  `E���  `E����  ^�����      C   ,  ag����  ag���  c)���  c)����  ag����      C   ,  dK����  dK���  f���  f����  dK����      C   ,  g/����  g/���  h����  h�����  g/����      C   ,  j����  j���  k����  k�����  j����      C   ,  8�����  8����  :����  :�����  8�����      C   ,  ;�����  ;����  =����  =�����  ;�����      C  , ,����  s����     U     U  s����  s      C  , ,����   �����  c   U  c   U   �����   �      C  , ,���������������G   U���G   U������������      C  , ,���������������   U���   U������������      C  , ,  8	  �  8	  ,  8�  ,  8�  �  8	  �      C  , ,  :�  �  :�  ,  ;�  ,  ;�  �  :�  �      C  , ,  =�  �  =�  ,  >{  ,  >{  �  =�  �      C  , ,  @�  �  @�  ,  A_  ,  A_  �  @�  �      C  , ,  C�  �  C�  ,  DC  ,  DC  �  C�  �      C  , ,  F}  �  F}  ,  G'  ,  G'  �  F}  �      C  , ,  Ia  �  Ia  ,  J  ,  J  �  Ia  �      C  , ,  LE  �  LE  ,  L�  ,  L�  �  LE  �      C  , ,  O)  �  O)  ,  O�  ,  O�  �  O)  �      C  , ,  R  �  R  ,  R�  ,  R�  �  R  �      C  , ,  T�  �  T�  ,  U�  ,  U�  �  T�  �      C  , ,  W�  �  W�  ,  X  ,  X  �  W�  �      C  , ,  Z�  �  Z�  ,  [c  ,  [c  �  Z�  �      C  , ,  ]�  �  ]�  ,  ^G  ,  ^G  �  ]�  �      C  , ,  `�  �  `�  ,  a+  ,  a+  �  `�  �      C  , ,  ce  �  ce  ,  d  ,  d  �  ce  �      C  , ,  fI  �  fI  ,  f�  ,  f�  �  fI  �      C  , ,  i-  �  i-  ,  i�  ,  i�  �  i-  �      C  , ,  l  �  l  ,  l�  ,  l�  �  l  �      C  , ,  R  �  R  �  R�  �  R�  �  R  �      C  , ,  T�  �  T�  �  U�  �  U�  �  T�  �      C  , ,  W�  �  W�  �  X  �  X  �  W�  �      C  , ,  Z�  �  Z�  �  [c  �  [c  �  Z�  �      C  , ,  ]�  �  ]�  �  ^G  �  ^G  �  ]�  �      C  , ,  `�  �  `�  �  a+  �  a+  �  `�  �      C  , ,  ce  �  ce  �  d  �  d  �  ce  �      C  , ,  fI  �  fI  �  f�  �  f�  �  fI  �      C  , ,  i-  �  i-  �  i�  �  i�  �  i-  �      C  , ,  l  �  l  �  l�  �  l�  �  l  �      C  , ,  S  s  S    T)    T)  s  S  s      C  , ,  Vc  s  Vc    W    W  s  Vc  s      C  , ,  YG  s  YG    Y�    Y�  s  YG  s      C  , ,  \+  s  \+    \�    \�  s  \+  s      C  , ,  _  s  _    _�    _�  s  _  s      C  , ,  a�  s  a�    b�    b�  s  a�  s      C  , ,  d�  s  d�    e�    e�  s  d�  s      C  , ,  g�  s  g�    he    he  s  g�  s      C  , ,  j�  s  j�    kI    kI  s  j�  s      C  , ,  R  R  R  �  R�  �  R�  R  R  R      C  , ,  T�  R  T�  �  U�  �  U�  R  T�  R      C  , ,  W�  R  W�  �  X  �  X  R  W�  R      C  , ,  Z�  R  Z�  �  [c  �  [c  R  Z�  R      C  , ,  ]�  R  ]�  �  ^G  �  ^G  R  ]�  R      C  , ,  `�  R  `�  �  a+  �  a+  R  `�  R      C  , ,  ce  R  ce  �  d  �  d  R  ce  R      C  , ,  fI  R  fI  �  f�  �  f�  R  fI  R      C  , ,  i-  R  i-  �  i�  �  i�  R  i-  R      C  , ,  l  R  l  �  l�  �  l�  R  l  R      C  , ,  :�  R  :�  �  ;�  �  ;�  R  :�  R      C  , ,  =�  R  =�  �  >{  �  >{  R  =�  R      C  , ,  @�  R  @�  �  A_  �  A_  R  @�  R      C  , ,  C�  R  C�  �  DC  �  DC  R  C�  R      C  , ,  F}  R  F}  �  G'  �  G'  R  F}  R      C  , ,  Ia  R  Ia  �  J  �  J  R  Ia  R      C  , ,  LE  R  LE  �  L�  �  L�  R  LE  R      C  , ,  O)  R  O)  �  O�  �  O�  R  O)  R      C  , ,  P�  s  P�    QE    QE  s  P�  s      C  , ,  6�  s  6�    7A    7A  s  6�  s      C  , ,  9{  s  9{    :%    :%  s  9{  s      C  , ,  <_  s  <_    =	    =	  s  <_  s      C  , ,  ?C  s  ?C    ?�    ?�  s  ?C  s      C  , ,  B'  s  B'    B�    B�  s  B'  s      C  , ,  E  s  E    E�    E�  s  E  s      C  , ,  G�  s  G�    H�    H�  s  G�  s      C  , ,  J�  s  J�    K}    K}  s  J�  s      C  , ,  M�  s  M�    Na    Na  s  M�  s      C  , ,  8	  �  8	  �  8�  �  8�  �  8	  �      C  , ,  :�  �  :�  �  ;�  �  ;�  �  :�  �      C  , ,  =�  �  =�  �  >{  �  >{  �  =�  �      C  , ,  @�  �  @�  �  A_  �  A_  �  @�  �      C  , ,  C�  �  C�  �  DC  �  DC  �  C�  �      C  , ,  F}  �  F}  �  G'  �  G'  �  F}  �      C  , ,  Ia  �  Ia  �  J  �  J  �  Ia  �      C  , ,  LE  �  LE  �  L�  �  L�  �  LE  �      C  , ,  O)  �  O)  �  O�  �  O�  �  O)  �      C  , ,  8	  R  8	  �  8�  �  8�  R  8	  R      C  , ,  8	    8	  �  8�  �  8�    8	        C  , ,  :�    :�  �  ;�  �  ;�    :�        C  , ,  =�    =�  �  >{  �  >{    =�        C  , ,  @�    @�  �  A_  �  A_    @�        C  , ,  C�    C�  �  DC  �  DC    C�        C  , ,  F}    F}  �  G'  �  G'    F}        C  , ,  Ia    Ia  �  J  �  J    Ia        C  , ,  LE    LE  �  L�  �  L�    LE        C  , ,  O)    O)  �  O�  �  O�    O)        C  , ,  8	  �  8	  \  8�  \  8�  �  8	  �      C  , ,  :�  �  :�  \  ;�  \  ;�  �  :�  �      C  , ,  =�  �  =�  \  >{  \  >{  �  =�  �      C  , ,  @�  �  @�  \  A_  \  A_  �  @�  �      C  , ,  C�  �  C�  \  DC  \  DC  �  C�  �      C  , ,  F}  �  F}  \  G'  \  G'  �  F}  �      C  , ,  Ia  �  Ia  \  J  \  J  �  Ia  �      C  , ,  LE  �  LE  \  L�  \  L�  �  LE  �      C  , ,  O)  �  O)  \  O�  \  O�  �  O)  �      C  , ,  8	  J  8	  �  8�  �  8�  J  8	  J      C  , ,  :�  J  :�  �  ;�  �  ;�  J  :�  J      C  , ,  =�  J  =�  �  >{  �  >{  J  =�  J      C  , ,  @�  J  @�  �  A_  �  A_  J  @�  J      C  , ,  C�  J  C�  �  DC  �  DC  J  C�  J      C  , ,  F}  J  F}  �  G'  �  G'  J  F}  J      C  , ,  Ia  J  Ia  �  J  �  J  J  Ia  J      C  , ,  LE  J  LE  �  L�  �  L�  J  LE  J      C  , ,  O)  J  O)  �  O�  �  O�  J  O)  J      C  , ,  i-    i-  �  i�  �  i�    i-        C  , ,  R  �  R  \  R�  \  R�  �  R  �      C  , ,  T�  �  T�  \  U�  \  U�  �  T�  �      C  , ,  W�  �  W�  \  X  \  X  �  W�  �      C  , ,  Z�  �  Z�  \  [c  \  [c  �  Z�  �      C  , ,  ]�  �  ]�  \  ^G  \  ^G  �  ]�  �      C  , ,  `�  �  `�  \  a+  \  a+  �  `�  �      C  , ,  ce  �  ce  \  d  \  d  �  ce  �      C  , ,  fI  �  fI  \  f�  \  f�  �  fI  �      C  , ,  i-  �  i-  \  i�  \  i�  �  i-  �      C  , ,  l  �  l  \  l�  \  l�  �  l  �      C  , ,  l    l  �  l�  �  l�    l        C  , ,  R    R  �  R�  �  R�    R        C  , ,  T�    T�  �  U�  �  U�    T�        C  , ,  W�    W�  �  X  �  X    W�        C  , ,  Z�    Z�  �  [c  �  [c    Z�        C  , ,  ]�    ]�  �  ^G  �  ^G    ]�        C  , ,  `�    `�  �  a+  �  a+    `�        C  , ,  ce    ce  �  d  �  d    ce        C  , ,  fI    fI  �  f�  �  f�    fI        C  , ,  R  J  R  �  R�  �  R�  J  R  J      C  , ,  T�  J  T�  �  U�  �  U�  J  T�  J      C  , ,  W�  J  W�  �  X  �  X  J  W�  J      C  , ,  Z�  J  Z�  �  [c  �  [c  J  Z�  J      C  , ,  ]�  J  ]�  �  ^G  �  ^G  J  ]�  J      C  , ,  `�  J  `�  �  a+  �  a+  J  `�  J      C  , ,  ce  J  ce  �  d  �  d  J  ce  J      C  , ,  fI  J  fI  �  f�  �  f�  J  fI  J      C  , ,  i-  J  i-  �  i�  �  i�  J  i-  J      C  , ,  l  J  l  �  l�  �  l�  J  l  J      C  , ,  !    !  �  �  �  �    !        C  , ,  !  �  !  �  �  �  �  �  !  �      C  , ,  !  �  !  \  �  \  �  �  !  �      C  , ,  !  R  !  �  �  �  �  R  !  R      C  , ,    �    ,  �  ,  �  �    �      C  , ,    �    ,  �  ,  �  �    �      C  , ,  �  �  �  ,  �  ,  �  �  �  �      C  , ,  	�  �  	�  ,  
s  ,  
s  �  	�  �      C  , ,  !  J  !  �  �  �  �  J  !  J      C  , ,  �  �  �  ,  W  ,  W  �  �  �      C  , ,  �  �  �  ,  ;  ,  ;  �  �  �      C  , ,  u  �  u  ,    ,    �  u  �      C  , ,  Y  �  Y  ,    ,    �  Y  �      C  , ,  =  �  =  ,  �  ,  �  �  =  �      C  , ,  !  �  !  ,  �  ,  �  �  !  �      C  , ,    �    ,  �  ,  �  �    �      C  , ,   �  �   �  ,  !�  ,  !�  �   �  �      C  , ,  #�  �  #�  ,  $w  ,  $w  �  #�  �      C  , ,  &�  �  &�  ,  '[  ,  '[  �  &�  �      C  , ,  )�  �  )�  ,  *?  ,  *?  �  )�  �      C  , ,  ,y  �  ,y  ,  -#  ,  -#  �  ,y  �      C  , ,  /]  �  /]  ,  0  ,  0  �  /]  �      C  , ,  2A  �  2A  ,  2�  ,  2�  �  2A  �      C  , ,  5%  �  5%  ,  5�  ,  5�  �  5%  �      C  , ,  5%  R  5%  �  5�  �  5�  R  5%  R      C  , ,  �  s  �    =    =  s  �  s      C  , ,  w  s  w     !     !  s  w  s      C  , ,  0�  s  0�    1y    1y  s  0�  s      C  , ,    �    �  �  �  �  �    �      C  , ,   �  �   �  �  !�  �  !�  �   �  �      C  , ,  #�  �  #�  �  $w  �  $w  �  #�  �      C  , ,  &�  �  &�  �  '[  �  '[  �  &�  �      C  , ,  )�  �  )�  �  *?  �  *?  �  )�  �      C  , ,  ,y  �  ,y  �  -#  �  -#  �  ,y  �      C  , ,  /]  �  /]  �  0  �  0  �  /]  �      C  , ,  2A  �  2A  �  2�  �  2�  �  2A  �      C  , ,  5%  �  5%  �  5�  �  5�  �  5%  �      C  , ,  3�  s  3�    4]    4]  s  3�  s      C  , ,  -�  s  -�    .�    .�  s  -�  s      C  , ,    R    �  �  �  �  R    R      C  , ,   �  R   �  �  !�  �  !�  R   �  R      C  , ,  #�  R  #�  �  $w  �  $w  R  #�  R      C  , ,  &�  R  &�  �  '[  �  '[  R  &�  R      C  , ,  )�  R  )�  �  *?  �  *?  R  )�  R      C  , ,  ,y  R  ,y  �  -#  �  -#  R  ,y  R      C  , ,  /]  R  /]  �  0  �  0  R  /]  R      C  , ,  2A  R  2A  �  2�  �  2�  R  2A  R      C  , ,  "[  s  "[    #    #  s  "[  s      C  , ,  %?  s  %?    %�    %�  s  %?  s      C  , ,  (#  s  (#    (�    (�  s  (#  s      C  , ,  +  s  +    +�    +�  s  +  s      C  , ,  	�  R  	�  �  
s  �  
s  R  	�  R      C  , ,    �    �  �  �  �  �    �      C  , ,    �    �  �  �  �  �    �      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,  �  R  �  �  W  �  W  R  �  R      C  , ,  �  R  �  �  ;  �  ;  R  �  R      C  , ,  u  R  u  �    �    R  u  R      C  , ,  Y  R  Y  �    �    R  Y  R      C  , ,  	�  �  	�  �  
s  �  
s  �  	�  �      C  , ,  =  R  =  �  �  �  �  R  =  R      C  , ,  ;  s  ;    �    �  s  ;  s      C  , ,  �  �  �  �  W  �  W  �  �  �      C  , ,  �  �  �  �  ;  �  ;  �  �  �      C  , ,  u  �  u  �    �    �  u  �      C  , ,  Y  �  Y  �    �    �  Y  �      C  , ,  =  �  =  �  �  �  �  �  =  �      C  , ,    s      �    �  s    s      C  , ,    s      �    �  s    s      C  , ,  �  s  �    �    �  s  �  s      C  , ,    R    �  �  �  �  R    R      C  , ,  �  s  �    u    u  s  �  s      C  , ,  �  s  �    Y    Y  s  �  s      C  , ,    R    �  �  �  �  R    R      C  , ,  �  R  �  �  �  �  �  R  �  R      C  , ,  �  s  �    9    9  s  �  s      C  , ,  s  s  s          s  s  s      C  , ,  W  s  W    	    	  s  W  s      C  , ,  �  J  �  �  ;  �  ;  J  �  J      C  , ,  u  J  u  �    �    J  u  J      C  , ,  Y  J  Y  �    �    J  Y  J      C  , ,  =  J  =  �  �  �  �  J  =  J      C  , ,  �    �  �  W  �  W    �        C  , ,  �    �  �  ;  �  ;    �        C  , ,  u    u  �    �      u        C  , ,  Y    Y  �    �      Y        C  , ,  =    =  �  �  �  �    =        C  , ,        �  �  �  �            C  , ,        �  �  �  �            C  , ,    �    \  �  \  �  �    �      C  , ,    �    \  �  \  �  �    �      C  , ,  �  �  �  \  �  \  �  �  �  �      C  , ,  	�  �  	�  \  
s  \  
s  �  	�  �      C  , ,  �  �  �  \  W  \  W  �  �  �      C  , ,  �  �  �  \  ;  \  ;  �  �  �      C  , ,  u  �  u  \    \    �  u  �      C  , ,  Y  �  Y  \    \    �  Y  �      C  , ,  =  �  =  \  �  \  �  �  =  �      C  , ,  �    �  �  �  �  �    �        C  , ,  	�    	�  �  
s  �  
s    	�        C  , ,    J    �  �  �  �  J    J      C  , ,    J    �  �  �  �  J    J      C  , ,  �  J  �  �  �  �  �  J  �  J      C  , ,  	�  J  	�  �  
s  �  
s  J  	�  J      C  , ,  �  J  �  �  W  �  W  J  �  J      C  , ,  )�  J  )�  �  *?  �  *?  J  )�  J      C  , ,  ,y  J  ,y  �  -#  �  -#  J  ,y  J      C  , ,  /]  J  /]  �  0  �  0  J  /]  J      C  , ,  2A  J  2A  �  2�  �  2�  J  2A  J      C  , ,  5%  J  5%  �  5�  �  5�  J  5%  J      C  , ,  #�  �  #�  \  $w  \  $w  �  #�  �      C  , ,  &�  �  &�  \  '[  \  '[  �  &�  �      C  , ,  )�  �  )�  \  *?  \  *?  �  )�  �      C  , ,  ,y  �  ,y  \  -#  \  -#  �  ,y  �      C  , ,  /]  �  /]  \  0  \  0  �  /]  �      C  , ,  2A  �  2A  \  2�  \  2�  �  2A  �      C  , ,  5%  �  5%  \  5�  \  5�  �  5%  �      C  , ,  #�    #�  �  $w  �  $w    #�        C  , ,  &�    &�  �  '[  �  '[    &�        C  , ,  )�    )�  �  *?  �  *?    )�        C  , ,  ,y    ,y  �  -#  �  -#    ,y        C  , ,  /]    /]  �  0  �  0    /]        C  , ,  2A    2A  �  2�  �  2�    2A        C  , ,  5%    5%  �  5�  �  5�    5%        C  , ,        �  �  �  �            C  , ,   �     �  �  !�  �  !�     �        C  , ,    �    \  �  \  �  �    �      C  , ,   �  �   �  \  !�  \  !�  �   �  �      C  , ,    J    �  �  �  �  J    J      C  , ,   �  J   �  �  !�  �  !�  J   �  J      C  , ,  #�  J  #�  �  $w  �  $w  J  #�  J      C  , ,  &�  J  &�  �  '[  �  '[  J  &�  J      C  , ,  !  	�  !  
�  �  
�  �  	�  !  	�      C  , ,  !  z  !  	$  �  	$  �  z  !  z      C  , ,  !    !  �  �  �  �    !        C  , ,  !  �  !  T  �  T  �  �  !  �      C  , ,  !  B  !  �  �  �  �  B  !  B      C  , ,  !  �  !  �  �  �  �  �  !  �      C  , ,  ,y  	�  ,y  
�  -#  
�  -#  	�  ,y  	�      C  , ,  /]  	�  /]  
�  0  
�  0  	�  /]  	�      C  , ,  2A  	�  2A  
�  2�  
�  2�  	�  2A  	�      C  , ,  5%  	�  5%  
�  5�  
�  5�  	�  5%  	�      C  , ,    	�    
�  �  
�  �  	�    	�      C  , ,    z    	$  �  	$  �  z    z      C  , ,   �  z   �  	$  !�  	$  !�  z   �  z      C  , ,  #�  z  #�  	$  $w  	$  $w  z  #�  z      C  , ,  &�  z  &�  	$  '[  	$  '[  z  &�  z      C  , ,  )�  z  )�  	$  *?  	$  *?  z  )�  z      C  , ,  ,y  z  ,y  	$  -#  	$  -#  z  ,y  z      C  , ,  /]  z  /]  	$  0  	$  0  z  /]  z      C  , ,  2A  z  2A  	$  2�  	$  2�  z  2A  z      C  , ,  5%  z  5%  	$  5�  	$  5�  z  5%  z      C  , ,   �  	�   �  
�  !�  
�  !�  	�   �  	�      C  , ,        �  �  �  �            C  , ,   �     �  �  !�  �  !�     �        C  , ,  #�    #�  �  $w  �  $w    #�        C  , ,  &�    &�  �  '[  �  '[    &�        C  , ,  )�    )�  �  *?  �  *?    )�        C  , ,  ,y    ,y  �  -#  �  -#    ,y        C  , ,  /]    /]  �  0  �  0    /]        C  , ,  2A    2A  �  2�  �  2�    2A        C  , ,  5%    5%  �  5�  �  5�    5%        C  , ,  #�  	�  #�  
�  $w  
�  $w  	�  #�  	�      C  , ,    �    T  �  T  �  �    �      C  , ,   �  �   �  T  !�  T  !�  �   �  �      C  , ,  #�  �  #�  T  $w  T  $w  �  #�  �      C  , ,  &�  �  &�  T  '[  T  '[  �  &�  �      C  , ,  )�  �  )�  T  *?  T  *?  �  )�  �      C  , ,  ,y  �  ,y  T  -#  T  -#  �  ,y  �      C  , ,  /]  �  /]  T  0  T  0  �  /]  �      C  , ,  2A  �  2A  T  2�  T  2�  �  2A  �      C  , ,  5%  �  5%  T  5�  T  5�  �  5%  �      C  , ,  &�  	�  &�  
�  '[  
�  '[  	�  &�  	�      C  , ,  )�  	�  )�  
�  *?  
�  *?  	�  )�  	�      C  , ,  Y    Y  �    �      Y        C  , ,  =    =  �  �  �  �    =        C  , ,  �  z  �  	$  W  	$  W  z  �  z      C  , ,  �  z  �  	$  ;  	$  ;  z  �  z      C  , ,  u  z  u  	$    	$    z  u  z      C  , ,  Y  z  Y  	$    	$    z  Y  z      C  , ,  =  z  =  	$  �  	$  �  z  =  z      C  , ,  Y  	�  Y  
�    
�    	�  Y  	�      C  , ,  =  	�  =  
�  �  
�  �  	�  =  	�      C  , ,  	�  	�  	�  
�  
s  
�  
s  	�  	�  	�      C  , ,  �  	�  �  
�  W  
�  W  	�  �  	�      C  , ,  �  	�  �  
�  ;  
�  ;  	�  �  	�      C  , ,    �    T  �  T  �  �    �      C  , ,    �    T  �  T  �  �    �      C  , ,  �  �  �  T  �  T  �  �  �  �      C  , ,  	�  �  	�  T  
s  T  
s  �  	�  �      C  , ,  �  �  �  T  W  T  W  �  �  �      C  , ,  �  �  �  T  ;  T  ;  �  �  �      C  , ,  u  �  u  T    T    �  u  �      C  , ,  Y  �  Y  T    T    �  Y  �      C  , ,  =  �  =  T  �  T  �  �  =  �      C  , ,  u  	�  u  
�    
�    	�  u  	�      C  , ,    z    	$  �  	$  �  z    z      C  , ,    z    	$  �  	$  �  z    z      C  , ,  �  z  �  	$  �  	$  �  z  �  z      C  , ,  	�  z  	�  	$  
s  	$  
s  z  	�  z      C  , ,        �  �  �  �            C  , ,        �  �  �  �            C  , ,  �    �  �  �  �  �    �        C  , ,  	�    	�  �  
s  �  
s    	�        C  , ,  �    �  �  W  �  W    �        C  , ,  �    �  �  ;  �  ;    �        C  , ,  u    u  �    �      u        C  , ,    	�    
�  �  
�  �  	�    	�      C  , ,    	�    
�  �  
�  �  	�    	�      C  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      C  , ,  �  B  �  �  ;  �  ;  B  �  B      C  , ,  u  B  u  �    �    B  u  B      C  , ,  Y  B  Y  �    �    B  Y  B      C  , ,  =  B  =  �  �  �  �  B  =  B      C  , ,    B    �  �  �  �  B    B      C  , ,    �    �  �  �  �  �    �      C  , ,    �    �  �  �  �  �    �      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,  	�  �  	�  �  
s  �  
s  �  	�  �      C  , ,  �  �  �  �  W  �  W  �  �  �      C  , ,  �  �  �  �  ;  �  ;  �  �  �      C  , ,  u  �  u  �    �    �  u  �      C  , ,  Y  �  Y  �    �    �  Y  �      C  , ,  =  �  =  �  �  �  �  �  =  �      C  , ,    B    �  �  �  �  B    B      C  , ,  �  B  �  �  �  �  �  B  �  B      C  , ,  �   �  �  c  9  c  9   �  �   �      C  , ,  s   �  s  c    c     �  s   �      C  , ,  W   �  W  c  	  c  	   �  W   �      C  , ,  ;   �  ;  c  �  c  �   �  ;   �      C  , ,     �    c  �  c  �   �     �      C  , ,     �    c  �  c  �   �     �      C  , ,  �   �  �  c  �  c  �   �  �   �      C  , ,  �   �  �  c  u  c  u   �  �   �      C  , ,  �   �  �  c  Y  c  Y   �  �   �      C  , ,  	�  B  	�  �  
s  �  
s  B  	�  B      C  , ,  �  B  �  �  W  �  W  B  �  B      C  , ,  &�  �  &�  �  '[  �  '[  �  &�  �      C  , ,  )�  �  )�  �  *?  �  *?  �  )�  �      C  , ,  ,y  �  ,y  �  -#  �  -#  �  ,y  �      C  , ,  /]  �  /]  �  0  �  0  �  /]  �      C  , ,  2A  �  2A  �  2�  �  2�  �  2A  �      C  , ,  5%  �  5%  �  5�  �  5�  �  5%  �      C  , ,   �  B   �  �  !�  �  !�  B   �  B      C  , ,  #�  B  #�  �  $w  �  $w  B  #�  B      C  , ,  &�  B  &�  �  '[  �  '[  B  &�  B      C  , ,  )�  B  )�  �  *?  �  *?  B  )�  B      C  , ,  ,y  B  ,y  �  -#  �  -#  B  ,y  B      C  , ,  /]  B  /]  �  0  �  0  B  /]  B      C  , ,  2A  B  2A  �  2�  �  2�  B  2A  B      C  , ,  5%  B  5%  �  5�  �  5�  B  5%  B      C  , ,    B    �  �  �  �  B    B      C  , ,    �    �  �  �  �  �    �      C  , ,  �   �  �  c  =  c  =   �  �   �      C  , ,  w   �  w  c   !  c   !   �  w   �      C  , ,  "[   �  "[  c  #  c  #   �  "[   �      C  , ,  %?   �  %?  c  %�  c  %�   �  %?   �      C  , ,  (#   �  (#  c  (�  c  (�   �  (#   �      C  , ,  +   �  +  c  +�  c  +�   �  +   �      C  , ,  -�   �  -�  c  .�  c  .�   �  -�   �      C  , ,  0�   �  0�  c  1y  c  1y   �  0�   �      C  , ,  3�   �  3�  c  4]  c  4]   �  3�   �      C  , ,   �  �   �  �  !�  �  !�  �   �  �      C  , ,  #�  �  #�  �  $w  �  $w  �  #�  �      C  , ,  R  �  R  T  R�  T  R�  �  R  �      C  , ,  T�  �  T�  T  U�  T  U�  �  T�  �      C  , ,  W�  �  W�  T  X  T  X  �  W�  �      C  , ,  Z�  �  Z�  T  [c  T  [c  �  Z�  �      C  , ,  ]�  �  ]�  T  ^G  T  ^G  �  ]�  �      C  , ,  `�  �  `�  T  a+  T  a+  �  `�  �      C  , ,  ce  �  ce  T  d  T  d  �  ce  �      C  , ,  fI  �  fI  T  f�  T  f�  �  fI  �      C  , ,  i-  �  i-  T  i�  T  i�  �  i-  �      C  , ,  l  �  l  T  l�  T  l�  �  l  �      C  , ,  R  	�  R  
�  R�  
�  R�  	�  R  	�      C  , ,  T�  	�  T�  
�  U�  
�  U�  	�  T�  	�      C  , ,  W�  	�  W�  
�  X  
�  X  	�  W�  	�      C  , ,  Z�  	�  Z�  
�  [c  
�  [c  	�  Z�  	�      C  , ,  ]�  	�  ]�  
�  ^G  
�  ^G  	�  ]�  	�      C  , ,  `�  	�  `�  
�  a+  
�  a+  	�  `�  	�      C  , ,  ce  	�  ce  
�  d  
�  d  	�  ce  	�      C  , ,  fI  	�  fI  
�  f�  
�  f�  	�  fI  	�      C  , ,  i-  	�  i-  
�  i�  
�  i�  	�  i-  	�      C  , ,  l  	�  l  
�  l�  
�  l�  	�  l  	�      C  , ,  R    R  �  R�  �  R�    R        C  , ,  T�    T�  �  U�  �  U�    T�        C  , ,  W�    W�  �  X  �  X    W�        C  , ,  Z�    Z�  �  [c  �  [c    Z�        C  , ,  ]�    ]�  �  ^G  �  ^G    ]�        C  , ,  `�    `�  �  a+  �  a+    `�        C  , ,  ce    ce  �  d  �  d    ce        C  , ,  fI    fI  �  f�  �  f�    fI        C  , ,  i-    i-  �  i�  �  i�    i-        C  , ,  l    l  �  l�  �  l�    l        C  , ,  R  z  R  	$  R�  	$  R�  z  R  z      C  , ,  T�  z  T�  	$  U�  	$  U�  z  T�  z      C  , ,  W�  z  W�  	$  X  	$  X  z  W�  z      C  , ,  Z�  z  Z�  	$  [c  	$  [c  z  Z�  z      C  , ,  ]�  z  ]�  	$  ^G  	$  ^G  z  ]�  z      C  , ,  `�  z  `�  	$  a+  	$  a+  z  `�  z      C  , ,  ce  z  ce  	$  d  	$  d  z  ce  z      C  , ,  fI  z  fI  	$  f�  	$  f�  z  fI  z      C  , ,  i-  z  i-  	$  i�  	$  i�  z  i-  z      C  , ,  l  z  l  	$  l�  	$  l�  z  l  z      C  , ,  C�    C�  �  DC  �  DC    C�        C  , ,  F}    F}  �  G'  �  G'    F}        C  , ,  Ia    Ia  �  J  �  J    Ia        C  , ,  LE    LE  �  L�  �  L�    LE        C  , ,  O)    O)  �  O�  �  O�    O)        C  , ,  @�  	�  @�  
�  A_  
�  A_  	�  @�  	�      C  , ,  C�  	�  C�  
�  DC  
�  DC  	�  C�  	�      C  , ,  F}  	�  F}  
�  G'  
�  G'  	�  F}  	�      C  , ,  Ia  	�  Ia  
�  J  
�  J  	�  Ia  	�      C  , ,  LE  	�  LE  
�  L�  
�  L�  	�  LE  	�      C  , ,  O)  	�  O)  
�  O�  
�  O�  	�  O)  	�      C  , ,  F}  �  F}  T  G'  T  G'  �  F}  �      C  , ,  Ia  �  Ia  T  J  T  J  �  Ia  �      C  , ,  LE  �  LE  T  L�  T  L�  �  LE  �      C  , ,  O)  �  O)  T  O�  T  O�  �  O)  �      C  , ,  8	  z  8	  	$  8�  	$  8�  z  8	  z      C  , ,  :�  z  :�  	$  ;�  	$  ;�  z  :�  z      C  , ,  =�  z  =�  	$  >{  	$  >{  z  =�  z      C  , ,  @�  z  @�  	$  A_  	$  A_  z  @�  z      C  , ,  C�  z  C�  	$  DC  	$  DC  z  C�  z      C  , ,  F}  z  F}  	$  G'  	$  G'  z  F}  z      C  , ,  Ia  z  Ia  	$  J  	$  J  z  Ia  z      C  , ,  LE  z  LE  	$  L�  	$  L�  z  LE  z      C  , ,  O)  z  O)  	$  O�  	$  O�  z  O)  z      C  , ,  =�  �  =�  T  >{  T  >{  �  =�  �      C  , ,  @�  �  @�  T  A_  T  A_  �  @�  �      C  , ,  C�  �  C�  T  DC  T  DC  �  C�  �      C  , ,  8	  	�  8	  
�  8�  
�  8�  	�  8	  	�      C  , ,  :�  	�  :�  
�  ;�  
�  ;�  	�  :�  	�      C  , ,  =�  	�  =�  
�  >{  
�  >{  	�  =�  	�      C  , ,  8	    8	  �  8�  �  8�    8	        C  , ,  :�    :�  �  ;�  �  ;�    :�        C  , ,  =�    =�  �  >{  �  >{    =�        C  , ,  @�    @�  �  A_  �  A_    @�        C  , ,  8	  �  8	  T  8�  T  8�  �  8	  �      C  , ,  :�  �  :�  T  ;�  T  ;�  �  :�  �      C  , ,  C�  B  C�  �  DC  �  DC  B  C�  B      C  , ,  F}  B  F}  �  G'  �  G'  B  F}  B      C  , ,  Ia  B  Ia  �  J  �  J  B  Ia  B      C  , ,  LE  B  LE  �  L�  �  L�  B  LE  B      C  , ,  O)  B  O)  �  O�  �  O�  B  O)  B      C  , ,  8	  B  8	  �  8�  �  8�  B  8	  B      C  , ,  8	  �  8	  �  8�  �  8�  �  8	  �      C  , ,  :�  �  :�  �  ;�  �  ;�  �  :�  �      C  , ,  =�  �  =�  �  >{  �  >{  �  =�  �      C  , ,  @�  �  @�  �  A_  �  A_  �  @�  �      C  , ,  C�  �  C�  �  DC  �  DC  �  C�  �      C  , ,  F}  �  F}  �  G'  �  G'  �  F}  �      C  , ,  Ia  �  Ia  �  J  �  J  �  Ia  �      C  , ,  LE  �  LE  �  L�  �  L�  �  LE  �      C  , ,  O)  �  O)  �  O�  �  O�  �  O)  �      C  , ,  :�  B  :�  �  ;�  �  ;�  B  :�  B      C  , ,  6�   �  6�  c  7A  c  7A   �  6�   �      C  , ,  9{   �  9{  c  :%  c  :%   �  9{   �      C  , ,  <_   �  <_  c  =	  c  =	   �  <_   �      C  , ,  ?C   �  ?C  c  ?�  c  ?�   �  ?C   �      C  , ,  B'   �  B'  c  B�  c  B�   �  B'   �      C  , ,  E   �  E  c  E�  c  E�   �  E   �      C  , ,  G�   �  G�  c  H�  c  H�   �  G�   �      C  , ,  J�   �  J�  c  K}  c  K}   �  J�   �      C  , ,  M�   �  M�  c  Na  c  Na   �  M�   �      C  , ,  P�   �  P�  c  QE  c  QE   �  P�   �      C  , ,  =�  B  =�  �  >{  �  >{  B  =�  B      C  , ,  @�  B  @�  �  A_  �  A_  B  @�  B      C  , ,  T�  �  T�  �  U�  �  U�  �  T�  �      C  , ,  W�  �  W�  �  X  �  X  �  W�  �      C  , ,  Z�  �  Z�  �  [c  �  [c  �  Z�  �      C  , ,  ]�  �  ]�  �  ^G  �  ^G  �  ]�  �      C  , ,  `�  �  `�  �  a+  �  a+  �  `�  �      C  , ,  ce  �  ce  �  d  �  d  �  ce  �      C  , ,  fI  �  fI  �  f�  �  f�  �  fI  �      C  , ,  i-  �  i-  �  i�  �  i�  �  i-  �      C  , ,  l  �  l  �  l�  �  l�  �  l  �      C  , ,  i-  B  i-  �  i�  �  i�  B  i-  B      C  , ,  l  B  l  �  l�  �  l�  B  l  B      C  , ,  R  B  R  �  R�  �  R�  B  R  B      C  , ,  T�  B  T�  �  U�  �  U�  B  T�  B      C  , ,  W�  B  W�  �  X  �  X  B  W�  B      C  , ,  Z�  B  Z�  �  [c  �  [c  B  Z�  B      C  , ,  ]�  B  ]�  �  ^G  �  ^G  B  ]�  B      C  , ,  `�  B  `�  �  a+  �  a+  B  `�  B      C  , ,  ce  B  ce  �  d  �  d  B  ce  B      C  , ,  S   �  S  c  T)  c  T)   �  S   �      C  , ,  Vc   �  Vc  c  W  c  W   �  Vc   �      C  , ,  YG   �  YG  c  Y�  c  Y�   �  YG   �      C  , ,  \+   �  \+  c  \�  c  \�   �  \+   �      C  , ,  _   �  _  c  _�  c  _�   �  _   �      C  , ,  a�   �  a�  c  b�  c  b�   �  a�   �      C  , ,  d�   �  d�  c  e�  c  e�   �  d�   �      C  , ,  g�   �  g�  c  he  c  he   �  g�   �      C  , ,  j�   �  j�  c  kI  c  kI   �  j�   �      C  , ,  fI  B  fI  �  f�  �  f�  B  fI  B      C  , ,  R  �  R  �  R�  �  R�  �  R  �      C  , ,���5  ���5  �����  �����  ���5        C  , ,���5  ����5  �����  �����  ����5  �      C  , ,���5  ����5  \����  \����  ����5  �      C  , ,���5  R���5  �����  �����  R���5  R      C  , ,���5  J���5  �����  �����  J���5  J      C  , ,���1  ����1  ,����  ,����  ����1  �      C  , ,���  ����  ,��Ϳ  ,��Ϳ  ����  �      C  , ,����  �����  ,��У  ,��У  �����  �      C  , ,����  �����  ,��Ӈ  ,��Ӈ  �����  �      C  , ,����  �����  ,���k  ,���k  �����  �      C  , ,��إ  ���إ  ,���O  ,���O  ���إ  �      C  , ,��ۉ  ���ۉ  ,���3  ,���3  ���ۉ  �      C  , ,���m  ����m  ,���  ,���  ����m  �      C  , ,���Q  ����Q  ,����  ,����  ����Q  �      C  , ,���5  ����5  ,����  ,����  ����5  �      C  , ,���  ����  ,����  ,����  ����  �      C  , ,����  �����  ,���  ,���  �����  �      C  , ,����  �����  ,���  ,���  �����  �      C  , ,����  �����  ,���o  ,���o  �����  �      C  , ,���  ����  ,���S  ,���S  ����  �      C  , ,����  �����  ,���7  ,���7  �����  �      C  , ,���q  ����q  ,���  ,���  ����q  �      C  , ,���U  ����U  ,����  ,����  ����U  �      C  , ,���9  ����9  ,����  ,����  ����9  �      C  , ,����  R����  ����  ����  R����  R      C  , ,����  R����  ����o  ����o  R����  R      C  , ,���  R���  ����S  ����S  R���  R      C  , ,����  R����  ����7  ����7  R����  R      C  , ,���q  R���q  ����  ����  R���q  R      C  , ,���U  R���U  �����  �����  R���U  R      C  , ,���9  R���9  �����  �����  R���9  R      C  , ,���7  s���7  ����  ����  s���7  s      C  , ,���  s���  ����  ����  s���  s      C  , ,����  s����  ����  ����  s����  s      C  , ,����  s����  ����  ����  s����  s      C  , ,����  s����  ���q  ���q  s����  s      C  , ,���  s���  ���Q  ���Q  s���  s      C  , ,���  s���  ���5  ���5  s���  s      C  , ,���  ����  �����  �����  ����  �      C  , ,����  �����  ����  ����  �����  �      C  , ,����  �����  ����  ����  �����  �      C  , ,����  �����  ����o  ����o  �����  �      C  , ,���  ����  ����S  ����S  ����  �      C  , ,����  �����  ����7  ����7  �����  �      C  , ,���q  ����q  ����  ����  ����q  �      C  , ,���U  ����U  �����  �����  ����U  �      C  , ,���9  ����9  �����  �����  ����9  �      C  , ,���o  s���o  ���  ���  s���o  s      C  , ,���S  s���S  ����  ����  s���S  s      C  , ,���  R���  �����  �����  R���  R      C  , ,����  R����  ����  ����  R����  R      C  , ,��إ  ���إ  ����O  ����O  ���إ  �      C  , ,��ۉ  ���ۉ  ����3  ����3  ���ۉ  �      C  , ,���m  ����m  ����  ����  ����m  �      C  , ,���Q  ����Q  �����  �����  ����Q  �      C  , ,��·  s��·  ���1  ���1  s��·  s      C  , ,���k  s���k  ���  ���  s���k  s      C  , ,���O  s���O  ����  ����  s���O  s      C  , ,���3  s���3  ����  ����  s���3  s      C  , ,���  s���  ����  ����  s���  s      C  , ,����  s����  ��ݥ  ��ݥ  s����  s      C  , ,����  s����  ����  ����  s����  s      C  , ,����  s����  ���m  ���m  s����  s      C  , ,��ˣ  s��ˣ  ���M  ���M  s��ˣ  s      C  , ,���1  ����1  �����  �����  ����1  �      C  , ,���  ����  ���Ϳ  ���Ϳ  ����  �      C  , ,���1  R���1  �����  �����  R���1  R      C  , ,���  R���  ���Ϳ  ���Ϳ  R���  R      C  , ,����  R����  ���У  ���У  R����  R      C  , ,����  R����  ���Ӈ  ���Ӈ  R����  R      C  , ,����  R����  ����k  ����k  R����  R      C  , ,��إ  R��إ  ����O  ����O  R��إ  R      C  , ,��ۉ  R��ۉ  ����3  ����3  R��ۉ  R      C  , ,���m  R���m  ����  ����  R���m  R      C  , ,���Q  R���Q  �����  �����  R���Q  R      C  , ,����  �����  ���У  ���У  �����  �      C  , ,����  �����  ���Ӈ  ���Ӈ  �����  �      C  , ,����  �����  ����k  ����k  �����  �      C  , ,����  J����  ���У  ���У  J����  J      C  , ,����  J����  ���Ӈ  ���Ӈ  J����  J      C  , ,����  J����  ����k  ����k  J����  J      C  , ,��إ  J��إ  ����O  ����O  J��إ  J      C  , ,��ۉ  J��ۉ  ����3  ����3  J��ۉ  J      C  , ,���m  J���m  ����  ����  J���m  J      C  , ,���Q  J���Q  �����  �����  J���Q  J      C  , ,����  ����  ����k  ����k  ����        C  , ,��إ  ��إ  ����O  ����O  ��إ        C  , ,��ۉ  ��ۉ  ����3  ����3  ��ۉ        C  , ,���m  ���m  ����  ����  ���m        C  , ,���Q  ���Q  �����  �����  ���Q        C  , ,���1  ���1  �����  �����  ���1        C  , ,���  ���  ���Ϳ  ���Ϳ  ���        C  , ,���1  ����1  \����  \����  ����1  �      C  , ,���  ����  \��Ϳ  \��Ϳ  ����  �      C  , ,����  �����  \��У  \��У  �����  �      C  , ,����  �����  \��Ӈ  \��Ӈ  �����  �      C  , ,����  �����  \���k  \���k  �����  �      C  , ,��إ  ���إ  \���O  \���O  ���إ  �      C  , ,��ۉ  ���ۉ  \���3  \���3  ���ۉ  �      C  , ,���m  ����m  \���  \���  ����m  �      C  , ,���Q  ����Q  \����  \����  ����Q  �      C  , ,����  ����  ���У  ���У  ����        C  , ,����  ����  ���Ӈ  ���Ӈ  ����        C  , ,���1  J���1  �����  �����  J���1  J      C  , ,���  J���  ���Ϳ  ���Ϳ  J���  J      C  , ,����  J����  ����  ����  J����  J      C  , ,����  J����  ����  ����  J����  J      C  , ,����  J����  ����o  ����o  J����  J      C  , ,���  J���  ����S  ����S  J���  J      C  , ,����  J����  ����7  ����7  J����  J      C  , ,���q  J���q  ����  ����  J���q  J      C  , ,���U  J���U  �����  �����  J���U  J      C  , ,���9  J���9  �����  �����  J���9  J      C  , ,����  �����  \���  \���  �����  �      C  , ,����  �����  \���o  \���o  �����  �      C  , ,���  ����  \���S  \���S  ����  �      C  , ,����  �����  \���7  \���7  �����  �      C  , ,���q  ����q  \���  \���  ����q  �      C  , ,���U  ����U  \����  \����  ����U  �      C  , ,���9  ����9  \����  \����  ����9  �      C  , ,����  ����  ����  ����  ����        C  , ,����  ����  ����o  ����o  ����        C  , ,���  ���  ����S  ����S  ���        C  , ,����  ����  ����7  ����7  ����        C  , ,���q  ���q  ����  ����  ���q        C  , ,���U  ���U  �����  �����  ���U        C  , ,���9  ���9  �����  �����  ���9        C  , ,���  ���  �����  �����  ���        C  , ,����  ����  ����  ����  ����        C  , ,���  ����  \����  \����  ����  �      C  , ,����  �����  \���  \���  �����  �      C  , ,���  J���  �����  �����  J���  J      C  , ,���E  ����E  ,����  ,����  ����E  �      C  , ,���)  ����)  ,����  ,����  ����)  �      C  , ,���  ����  ,����  ,����  ����  �      C  , ,����  �����  ,����  ,����  �����  �      C  , ,����  �����  ,���  ,���  �����  �      C  , ,����  �����  ,���c  ,���c  �����  �      C  , ,����  �����  ,���G  ,���G  �����  �      C  , ,����  �����  ,���+  ,���+  �����  �      C  , ,���e  ����e  ,���  ,���  ����e  �      C  , ,���I  ����I  ,����  ,����  ����I  �      C  , ,���-  ����-  ,����  ,����  ����-  �      C  , ,���  ����  ,����  ,����  ����  �      C  , ,����  �����  ,����  ,����  �����  �      C  , ,����  �����  ,����  ,����  �����  �      C  , ,����  �����  ,���g  ,���g  �����  �      C  , ,����  �����  ,���K  ,���K  �����  �      C  , ,����  �����  ,���/  ,���/  �����  �      C  , ,���i  ����i  ,���  ,���  ����i  �      C  , ,���M  ����M  ,����  ,����  ����M  �      C  , ,���-  ����-  �����  �����  ����-  �      C  , ,���  ����  �����  �����  ����  �      C  , ,����  �����  �����  �����  �����  �      C  , ,����  �����  �����  �����  �����  �      C  , ,����  �����  ����g  ����g  �����  �      C  , ,����  �����  ����K  ����K  �����  �      C  , ,����  �����  ����/  ����/  �����  �      C  , ,���i  ����i  ����  ����  ����i  �      C  , ,���M  ����M  �����  �����  ����M  �      C  , ,����  s����  ���e  ���e  s����  s      C  , ,����  s����  ���I  ���I  s����  s      C  , ,����  s����  ���-  ���-  s����  s      C  , ,���g  s���g  ���  ���  s���g  s      C  , ,���K  s���K  ����  ����  s���K  s      C  , ,���/  s���/  ����  ����  s���/  s      C  , ,���  s���  ����  ����  s���  s      C  , ,����  s����  ��á  ��á  s����  s      C  , ,����  s����  ��ƅ  ��ƅ  s����  s      C  , ,��ȿ  s��ȿ  ���i  ���i  s��ȿ  s      C  , ,���-  R���-  �����  �����  R���-  R      C  , ,���  R���  �����  �����  R���  R      C  , ,����  R����  �����  �����  R����  R      C  , ,����  R����  �����  �����  R����  R      C  , ,����  R����  ����g  ����g  R����  R      C  , ,����  R����  ����K  ����K  R����  R      C  , ,����  R����  ����/  ����/  R����  R      C  , ,���i  R���i  ����  ����  R���i  R      C  , ,���M  R���M  �����  �����  R���M  R      C  , ,����  R����  ����  ����  R����  R      C  , ,����  R����  ����c  ����c  R����  R      C  , ,����  R����  ����G  ����G  R����  R      C  , ,����  R����  ����+  ����+  R����  R      C  , ,���e  R���e  ����  ����  R���e  R      C  , ,���I  R���I  �����  �����  R���I  R      C  , ,����  s����  ����  ����  s����  s      C  , ,����  s����  ���E  ���E  s����  s      C  , ,����  s����  ����  ����  s����  s      C  , ,���)  R���)  �����  �����  R���)  R      C  , ,���+  s���+  ����  ����  s���+  s      C  , ,���  s���  ����  ����  s���  s      C  , ,���c  s���c  ���  ���  s���c  s      C  , ,���G  s���G  ����  ����  s���G  s      C  , ,����  s����  ���a  ���a  s����  s      C  , ,���E  R���E  �����  �����  R���E  R      C  , ,���E  ����E  �����  �����  ����E  �      C  , ,���)  ����)  �����  �����  ����)  �      C  , ,���  ����  �����  �����  ����  �      C  , ,����  �����  �����  �����  �����  �      C  , ,����  �����  ����  ����  �����  �      C  , ,����  �����  ����c  ����c  �����  �      C  , ,����  �����  ����G  ����G  �����  �      C  , ,����  �����  ����+  ����+  �����  �      C  , ,���e  ����e  ����  ����  ����e  �      C  , ,���I  ����I  �����  �����  ����I  �      C  , ,���  R���  �����  �����  R���  R      C  , ,����  R����  �����  �����  R����  R      C  , ,���  s���  ���)  ���)  s���  s      C  , ,���E  ���E  �����  �����  ���E        C  , ,���E  J���E  �����  �����  J���E  J      C  , ,���)  J���)  �����  �����  J���)  J      C  , ,���  J���  �����  �����  J���  J      C  , ,����  J����  �����  �����  J����  J      C  , ,����  J����  ����  ����  J����  J      C  , ,����  J����  ����c  ����c  J����  J      C  , ,����  J����  ����G  ����G  J����  J      C  , ,����  J����  ����+  ����+  J����  J      C  , ,���e  J���e  ����  ����  J���e  J      C  , ,���I  J���I  �����  �����  J���I  J      C  , ,���)  ���)  �����  �����  ���)        C  , ,���  ���  �����  �����  ���        C  , ,����  ����  �����  �����  ����        C  , ,����  ����  ����  ����  ����        C  , ,����  ����  ����c  ����c  ����        C  , ,����  ����  ����G  ����G  ����        C  , ,����  ����  ����+  ����+  ����        C  , ,���e  ���e  ����  ����  ���e        C  , ,���E  ����E  \����  \����  ����E  �      C  , ,���)  ����)  \����  \����  ����)  �      C  , ,���  ����  \����  \����  ����  �      C  , ,����  �����  \����  \����  �����  �      C  , ,����  �����  \���  \���  �����  �      C  , ,����  �����  \���c  \���c  �����  �      C  , ,����  �����  \���G  \���G  �����  �      C  , ,����  �����  \���+  \���+  �����  �      C  , ,���e  ����e  \���  \���  ����e  �      C  , ,���I  ����I  \����  \����  ����I  �      C  , ,���I  ���I  �����  �����  ���I        C  , ,����  ����  �����  �����  ����        C  , ,����  ����  ����g  ����g  ����        C  , ,����  ����  ����K  ����K  ����        C  , ,����  ����  ����/  ����/  ����        C  , ,���i  ���i  ����  ����  ���i        C  , ,���M  ���M  �����  �����  ���M        C  , ,���-  J���-  �����  �����  J���-  J      C  , ,���  J���  �����  �����  J���  J      C  , ,����  J����  �����  �����  J����  J      C  , ,����  J����  �����  �����  J����  J      C  , ,����  J����  ����g  ����g  J����  J      C  , ,����  J����  ����K  ����K  J����  J      C  , ,����  J����  ����/  ����/  J����  J      C  , ,���i  J���i  ����  ����  J���i  J      C  , ,���M  J���M  �����  �����  J���M  J      C  , ,���-  ���-  �����  �����  ���-        C  , ,���  ���  �����  �����  ���        C  , ,���-  ����-  \����  \����  ����-  �      C  , ,���  ����  \����  \����  ����  �      C  , ,����  �����  \����  \����  �����  �      C  , ,����  �����  \����  \����  �����  �      C  , ,����  �����  \���g  \���g  �����  �      C  , ,����  �����  \���K  \���K  �����  �      C  , ,����  �����  \���/  \���/  �����  �      C  , ,���i  ����i  \���  \���  ����i  �      C  , ,���M  ����M  \����  \����  ����M  �      C  , ,����  ����  �����  �����  ����        C  , ,���-  ����-  T����  T����  ����-  �      C  , ,���  ����  T����  T����  ����  �      C  , ,����  �����  T����  T����  �����  �      C  , ,����  �����  T����  T����  �����  �      C  , ,����  �����  T���g  T���g  �����  �      C  , ,����  �����  T���K  T���K  �����  �      C  , ,����  �����  T���/  T���/  �����  �      C  , ,���i  ����i  T���  T���  ����i  �      C  , ,���M  ����M  T����  T����  ����M  �      C  , ,���-  ���-  �����  �����  ���-        C  , ,���  ���  �����  �����  ���        C  , ,����  ����  �����  �����  ����        C  , ,����  ����  �����  �����  ����        C  , ,����  ����  ����g  ����g  ����        C  , ,����  ����  ����K  ����K  ����        C  , ,����  ����  ����/  ����/  ����        C  , ,���i  ���i  ����  ����  ���i        C  , ,���M  ���M  �����  �����  ���M        C  , ,����  	�����  
�����  
�����  	�����  	�      C  , ,����  	�����  
�����  
�����  	�����  	�      C  , ,����  	�����  
����g  
����g  	�����  	�      C  , ,����  	�����  
����K  
����K  	�����  	�      C  , ,����  	�����  
����/  
����/  	�����  	�      C  , ,���i  	����i  
����  
����  	����i  	�      C  , ,���M  	����M  
�����  
�����  	����M  	�      C  , ,���-  z���-  	$����  	$����  z���-  z      C  , ,���  z���  	$����  	$����  z���  z      C  , ,����  z����  	$����  	$����  z����  z      C  , ,����  z����  	$����  	$����  z����  z      C  , ,����  z����  	$���g  	$���g  z����  z      C  , ,����  z����  	$���K  	$���K  z����  z      C  , ,����  z����  	$���/  	$���/  z����  z      C  , ,���i  z���i  	$���  	$���  z���i  z      C  , ,���M  z���M  	$����  	$����  z���M  z      C  , ,���-  	����-  
�����  
�����  	����-  	�      C  , ,���  	����  
�����  
�����  	����  	�      C  , ,����  �����  T���+  T���+  �����  �      C  , ,����  	�����  
�����  
�����  	�����  	�      C  , ,����  	�����  
����  
����  	�����  	�      C  , ,����  	�����  
����c  
����c  	�����  	�      C  , ,����  	�����  
����G  
����G  	�����  	�      C  , ,����  	�����  
����+  
����+  	�����  	�      C  , ,���e  	����e  
����  
����  	����e  	�      C  , ,���E  z���E  	$����  	$����  z���E  z      C  , ,���)  z���)  	$����  	$����  z���)  z      C  , ,���  z���  	$����  	$����  z���  z      C  , ,����  z����  	$����  	$����  z����  z      C  , ,����  z����  	$���  	$���  z����  z      C  , ,����  z����  	$���c  	$���c  z����  z      C  , ,����  z����  	$���G  	$���G  z����  z      C  , ,����  z����  	$���+  	$���+  z����  z      C  , ,���e  z���e  	$���  	$���  z���e  z      C  , ,���I  z���I  	$����  	$����  z���I  z      C  , ,���e  ����e  T���  T���  ����e  �      C  , ,����  ����  �����  �����  ����        C  , ,����  ����  ����  ����  ����        C  , ,����  ����  ����c  ����c  ����        C  , ,����  ����  ����G  ����G  ����        C  , ,����  ����  ����+  ����+  ����        C  , ,���e  ���e  ����  ����  ���e        C  , ,���I  ���I  �����  �����  ���I        C  , ,���I  ����I  T����  T����  ����I  �      C  , ,���I  	����I  
�����  
�����  	����I  	�      C  , ,����  �����  T���c  T���c  �����  �      C  , ,����  �����  T���G  T���G  �����  �      C  , ,���E  ���E  �����  �����  ���E        C  , ,���)  ���)  �����  �����  ���)        C  , ,���  ���  �����  �����  ���        C  , ,���E  ����E  T����  T����  ����E  �      C  , ,���)  ����)  T����  T����  ����)  �      C  , ,���  ����  T����  T����  ����  �      C  , ,����  �����  T����  T����  �����  �      C  , ,����  �����  T���  T���  �����  �      C  , ,���E  	����E  
�����  
�����  	����E  	�      C  , ,���)  	����)  
�����  
�����  	����)  	�      C  , ,���  	����  
�����  
�����  	����  	�      C  , ,����  B����  ����c  ����c  B����  B      C  , ,����  B����  ����G  ����G  B����  B      C  , ,����  B����  ����+  ����+  B����  B      C  , ,���e  B���e  ����  ����  B���e  B      C  , ,���I  B���I  �����  �����  B���I  B      C  , ,����  �����  ����c  ����c  �����  �      C  , ,����  �����  ����G  ����G  �����  �      C  , ,����  �����  ����+  ����+  �����  �      C  , ,���e  ����e  ����  ����  ����e  �      C  , ,���I  ����I  �����  �����  ����I  �      C  , ,���E  ����E  �����  �����  ����E  �      C  , ,���)  ����)  �����  �����  ����)  �      C  , ,���  ����  �����  �����  ����  �      C  , ,����  �����  �����  �����  �����  �      C  , ,����  �����  ����  ����  �����  �      C  , ,���E  B���E  �����  �����  B���E  B      C  , ,���)  B���)  �����  �����  B���)  B      C  , ,���  B���  �����  �����  B���  B      C  , ,����   �����  c���a  c���a   �����   �      C  , ,����   �����  c���E  c���E   �����   �      C  , ,���   ����  c���)  c���)   ����   �      C  , ,���c   ����c  c���  c���   ����c   �      C  , ,���G   ����G  c����  c����   ����G   �      C  , ,���+   ����+  c����  c����   ����+   �      C  , ,���   ����  c����  c����   ����   �      C  , ,����   �����  c����  c����   �����   �      C  , ,����   �����  c����  c����   �����   �      C  , ,����  B����  �����  �����  B����  B      C  , ,����  B����  ����  ����  B����  B      C  , ,����  B����  ����K  ����K  B����  B      C  , ,����  B����  ����/  ����/  B����  B      C  , ,���i  B���i  ����  ����  B���i  B      C  , ,���M  B���M  �����  �����  B���M  B      C  , ,���-  ����-  �����  �����  ����-  �      C  , ,���  ����  �����  �����  ����  �      C  , ,����   �����  c���e  c���e   �����   �      C  , ,����   �����  c���I  c���I   �����   �      C  , ,����   �����  c���-  c���-   �����   �      C  , ,���g   ����g  c���  c���   ����g   �      C  , ,���K   ����K  c����  c����   ����K   �      C  , ,���/   ����/  c����  c����   ����/   �      C  , ,���   ����  c����  c����   ����   �      C  , ,����   �����  c��á  c��á   �����   �      C  , ,����   �����  c��ƅ  c��ƅ   �����   �      C  , ,��ȿ   ���ȿ  c���i  c���i   ���ȿ   �      C  , ,����  �����  �����  �����  �����  �      C  , ,����  �����  �����  �����  �����  �      C  , ,����  �����  ����g  ����g  �����  �      C  , ,����  �����  ����K  ����K  �����  �      C  , ,����  �����  ����/  ����/  �����  �      C  , ,���i  ����i  ����  ����  ����i  �      C  , ,���M  ����M  �����  �����  ����M  �      C  , ,���-  B���-  �����  �����  B���-  B      C  , ,���  B���  �����  �����  B���  B      C  , ,����  B����  �����  �����  B����  B      C  , ,����  B����  �����  �����  B����  B      C  , ,����  B����  ����g  ����g  B����  B      C  , ,���5  ����5  �����  �����  ����5  �      C  , ,���5  ���5  �����  �����  ���5        C  , ,���5  B���5  �����  �����  B���5  B      C  , ,���5  ����5  T����  T����  ����5  �      C  , ,���5  z���5  	$����  	$����  z���5  z      C  , ,���5  	����5  
�����  
�����  	����5  	�      C  , ,���  ���  ����S  ����S  ���        C  , ,����  ����  ����7  ����7  ����        C  , ,���q  ���q  ����  ����  ���q        C  , ,���U  ���U  �����  �����  ���U        C  , ,���9  ���9  �����  �����  ���9        C  , ,���  ���  �����  �����  ���        C  , ,����  ����  ����  ����  ����        C  , ,���  ����  T����  T����  ����  �      C  , ,����  �����  T���  T���  �����  �      C  , ,����  �����  T���  T���  �����  �      C  , ,����  �����  T���o  T���o  �����  �      C  , ,���  ����  T���S  T���S  ����  �      C  , ,����  �����  T���7  T���7  �����  �      C  , ,���q  ����q  T���  T���  ����q  �      C  , ,���U  ����U  T����  T����  ����U  �      C  , ,���9  ����9  T����  T����  ����9  �      C  , ,����  ����  ����  ����  ����        C  , ,���  z���  	$����  	$����  z���  z      C  , ,����  z����  	$���  	$���  z����  z      C  , ,����  z����  	$���  	$���  z����  z      C  , ,����  z����  	$���o  	$���o  z����  z      C  , ,���  z���  	$���S  	$���S  z���  z      C  , ,����  z����  	$���7  	$���7  z����  z      C  , ,���q  z���q  	$���  	$���  z���q  z      C  , ,���U  z���U  	$����  	$����  z���U  z      C  , ,���9  z���9  	$����  	$����  z���9  z      C  , ,����  ����  ����o  ����o  ����        C  , ,���  	����  
�����  
�����  	����  	�      C  , ,����  	�����  
����  
����  	�����  	�      C  , ,����  	�����  
����  
����  	�����  	�      C  , ,����  	�����  
����o  
����o  	�����  	�      C  , ,���  	����  
����S  
����S  	����  	�      C  , ,����  	�����  
����7  
����7  	�����  	�      C  , ,���q  	����q  
����  
����  	����q  	�      C  , ,���U  	����U  
�����  
�����  	����U  	�      C  , ,���9  	����9  
�����  
�����  	����9  	�      C  , ,����  z����  	$��У  	$��У  z����  z      C  , ,����  z����  	$��Ӈ  	$��Ӈ  z����  z      C  , ,����  z����  	$���k  	$���k  z����  z      C  , ,��إ  z��إ  	$���O  	$���O  z��إ  z      C  , ,��ۉ  z��ۉ  	$���3  	$���3  z��ۉ  z      C  , ,���m  z���m  	$���  	$���  z���m  z      C  , ,���Q  z���Q  	$����  	$����  z���Q  z      C  , ,���  ����  T��Ϳ  T��Ϳ  ����  �      C  , ,����  �����  T��У  T��У  �����  �      C  , ,����  �����  T��Ӈ  T��Ӈ  �����  �      C  , ,����  �����  T���k  T���k  �����  �      C  , ,��إ  ���إ  T���O  T���O  ���إ  �      C  , ,��ۉ  ���ۉ  T���3  T���3  ���ۉ  �      C  , ,���m  ����m  T���  T���  ����m  �      C  , ,���Q  ����Q  T����  T����  ����Q  �      C  , ,����  ����  ���У  ���У  ����        C  , ,����  ����  ���Ӈ  ���Ӈ  ����        C  , ,���1  	����1  
�����  
�����  	����1  	�      C  , ,���  	����  
���Ϳ  
���Ϳ  	����  	�      C  , ,����  	�����  
���У  
���У  	�����  	�      C  , ,����  	�����  
���Ӈ  
���Ӈ  	�����  	�      C  , ,����  	�����  
����k  
����k  	�����  	�      C  , ,��إ  	���إ  
����O  
����O  	���إ  	�      C  , ,��ۉ  	���ۉ  
����3  
����3  	���ۉ  	�      C  , ,���m  	����m  
����  
����  	����m  	�      C  , ,���Q  	����Q  
�����  
�����  	����Q  	�      C  , ,����  ����  ����k  ����k  ����        C  , ,��إ  ��إ  ����O  ����O  ��إ        C  , ,��ۉ  ��ۉ  ����3  ����3  ��ۉ        C  , ,���m  ���m  ����  ����  ���m        C  , ,���Q  ���Q  �����  �����  ���Q        C  , ,���1  ���1  �����  �����  ���1        C  , ,���  ���  ���Ϳ  ���Ϳ  ���        C  , ,���1  ����1  T����  T����  ����1  �      C  , ,���1  z���1  	$����  	$����  z���1  z      C  , ,���  z���  	$��Ϳ  	$��Ϳ  z���  z      C  , ,����  �����  ���У  ���У  �����  �      C  , ,����  �����  ���Ӈ  ���Ӈ  �����  �      C  , ,����  �����  ����k  ����k  �����  �      C  , ,��ˣ   ���ˣ  c���M  c���M   ���ˣ   �      C  , ,��·   ���·  c���1  c���1   ���·   �      C  , ,���k   ����k  c���  c���   ����k   �      C  , ,���O   ����O  c����  c����   ����O   �      C  , ,���3   ����3  c����  c����   ����3   �      C  , ,���   ����  c����  c����   ����   �      C  , ,����   �����  c��ݥ  c��ݥ   �����   �      C  , ,����   �����  c����  c����   �����   �      C  , ,����   �����  c���m  c���m   �����   �      C  , ,��إ  ���إ  ����O  ����O  ���إ  �      C  , ,��ۉ  ���ۉ  ����3  ����3  ���ۉ  �      C  , ,���m  ����m  ����  ����  ����m  �      C  , ,���1  B���1  �����  �����  B���1  B      C  , ,���  B���  ���Ϳ  ���Ϳ  B���  B      C  , ,����  B����  ���У  ���У  B����  B      C  , ,����  B����  ���Ӈ  ���Ӈ  B����  B      C  , ,����  B����  ����k  ����k  B����  B      C  , ,��إ  B��إ  ����O  ����O  B��إ  B      C  , ,��ۉ  B��ۉ  ����3  ����3  B��ۉ  B      C  , ,���m  B���m  ����  ����  B���m  B      C  , ,���Q  B���Q  �����  �����  B���Q  B      C  , ,���Q  ����Q  �����  �����  ����Q  �      C  , ,���1  ����1  �����  �����  ����1  �      C  , ,���  ����  ���Ϳ  ���Ϳ  ����  �      C  , ,���U  ����U  �����  �����  ����U  �      C  , ,���9  ����9  �����  �����  ����9  �      C  , ,���  ����  �����  �����  ����  �      C  , ,����  �����  ����  ����  �����  �      C  , ,���  B���  �����  �����  B���  B      C  , ,���   ����  c���Q  c���Q   ����   �      C  , ,���   ����  c���5  c���5   ����   �      C  , ,���o   ����o  c���  c���   ����o   �      C  , ,���S   ����S  c����  c����   ����S   �      C  , ,���7   ����7  c����  c����   ����7   �      C  , ,���   ����  c����  c����   ����   �      C  , ,����   �����  c����  c����   �����   �      C  , ,����   �����  c����  c����   �����   �      C  , ,����   �����  c���q  c���q   �����   �      C  , ,����  B����  ����  ����  B����  B      C  , ,����  B����  ����  ����  B����  B      C  , ,����  B����  ����o  ����o  B����  B      C  , ,���  B���  ����S  ����S  B���  B      C  , ,����  B����  ����7  ����7  B����  B      C  , ,���q  B���q  ����  ����  B���q  B      C  , ,���U  B���U  �����  �����  B���U  B      C  , ,���9  B���9  �����  �����  B���9  B      C  , ,����  �����  ����  ����  �����  �      C  , ,����  �����  ����o  ����o  �����  �      C  , ,���  ����  ����S  ����S  ����  �      C  , ,����  �����  ����7  ����7  �����  �      C  , ,���q  ����q  ����  ����  ����q  �      C  , ,���5���|���5���&�������&�������|���5���|      C  , ,���5������5����������������������5���      C  , ,���5�������5���V�������V�����������5����      C  , ,���5���D���5�������������������D���5���D      C  , ,���5�������5�����������������������5����      C  , ,���5���t���5�����������������t���5���t      C  , ,���������������G�������G����������������      C  , ,���������������G�������G����������������      C  , ,���������������G���q���G���q������������      C  , ,�������������G���Q���G���Q�����������      C  , ,������|������&�������&�������|������|      C  , ,�������|�������&������&������|�������|      C  , ,�������|�������&������&������|�������|      C  , ,�������|�������&���o���&���o���|�������|      C  , ,������|������&���S���&���S���|������|      C  , ,�������|�������&���7���&���7���|�������|      C  , ,���q���|���q���&������&������|���q���|      C  , ,���U���|���U���&�������&�������|���U���|      C  , ,���9���|���9���&�������&�������|���9���|      C  , ,�������������G���5���G���5�����������      C  , ,����������������������������������      C  , ,�����������������������������������      C  , ,�����������������������������������      C  , ,������������������o�������o����������      C  , ,����������������S�������S���������      C  , ,������������������7�������7����������      C  , ,���q������q��������������������q���      C  , ,���U������U����������������������U���      C  , ,���9������9����������������������9���      C  , ,���o�������o���G������G����������o����      C  , ,���S�������S���G�������G�����������S����      C  , ,���7�������7���G�������G�����������7����      C  , ,�������������G�������G���������������      C  , ,���������������G��ݥ���G��ݥ������������      C  , ,���������������G�������G����������������      C  , ,���������������G���m���G���m������������      C  , ,���1���|���1���&�������&�������|���1���|      C  , ,���1������1����������������������1���      C  , ,���������������Ϳ������Ϳ���������      C  , ,�����������������У������У����������      C  , ,�����������������Ӈ������Ӈ����������      C  , ,������������������k�������k����������      C  , ,��إ�����إ�������O�������O�����إ���      C  , ,��ۉ�����ۉ�������3�������3�����ۉ���      C  , ,���m������m��������������������m���      C  , ,���Q������Q����������������������Q���      C  , ,������|������&��Ϳ���&��Ϳ���|������|      C  , ,�������|�������&��У���&��У���|�������|      C  , ,�������|�������&��Ӈ���&��Ӈ���|�������|      C  , ,�������|�������&���k���&���k���|�������|      C  , ,��إ���|��إ���&���O���&���O���|��إ���|      C  , ,��ۉ���|��ۉ���&���3���&���3���|��ۉ���|      C  , ,���m���|���m���&������&������|���m���|      C  , ,���Q���|���Q���&�������&�������|���Q���|      C  , ,��ˣ������ˣ���G���M���G���M������ˣ����      C  , ,��·������·���G���1���G���1������·����      C  , ,���k�������k���G������G����������k����      C  , ,���O�������O���G�������G�����������O����      C  , ,���3�������3���G�������G�����������3����      C  , ,�������������G�������G���������������      C  , ,���������������V���k���V���k������������      C  , ,��إ������إ���V���O���V���O������إ����      C  , ,��ۉ������ۉ���V���3���V���3������ۉ����      C  , ,���m�������m���V������V����������m����      C  , ,���Q�������Q���V�������V�����������Q����      C  , ,���1�������1���V�������V�����������1����      C  , ,���1���D���1�������������������D���1���D      C  , ,������D���������Ϳ������Ϳ���D������D      C  , ,�������D����������У������У���D�������D      C  , ,�������D����������Ӈ������Ӈ���D�������D      C  , ,�������D�����������k�������k���D�������D      C  , ,��إ���D��إ�������O�������O���D��إ���D      C  , ,��ۉ���D��ۉ�������3�������3���D��ۉ���D      C  , ,���m���D���m�����������������D���m���D      C  , ,���Q���D���Q�������������������D���Q���D      C  , ,�������������V��Ϳ���V��Ϳ�����������      C  , ,���1�������1�����������������������1����      C  , ,����������������Ϳ������Ϳ�����������      C  , ,������������������У������У������������      C  , ,������������������Ӈ������Ӈ������������      C  , ,�������������������k�������k������������      C  , ,��إ������إ�������O�������O������إ����      C  , ,��ۉ������ۉ�������3�������3������ۉ����      C  , ,���m�������m���������������������m����      C  , ,���Q�������Q�����������������������Q����      C  , ,���������������V��У���V��У������������      C  , ,���1���t���1�����������������t���1���t      C  , ,������t��������Ϳ�����Ϳ���t������t      C  , ,�������t���������У�����У���t�������t      C  , ,�������t���������Ӈ�����Ӈ���t�������t      C  , ,�������t����������k������k���t�������t      C  , ,��إ���t��إ������O������O���t��إ���t      C  , ,��ۉ���t��ۉ������3������3���t��ۉ���t      C  , ,���m���t���m���������������t���m���t      C  , ,���Q���t���Q�����������������t���Q���t      C  , ,���������������V��Ӈ���V��Ӈ������������      C  , ,���������������V���o���V���o������������      C  , ,�������������V���S���V���S�����������      C  , ,���������������V���7���V���7������������      C  , ,���q�������q���V������V����������q����      C  , ,���U�������U���V�������V�����������U����      C  , ,���9�������9���V�������V�����������9����      C  , ,�������������V�������V���������������      C  , ,������D����������������������D������D      C  , ,�������������������������������������      C  , ,��������������������������������������      C  , ,��������������������������������������      C  , ,�������������������o�������o������������      C  , ,�����������������S�������S�����������      C  , ,�������������������7�������7������������      C  , ,���q�������q���������������������q����      C  , ,���U�������U�����������������������U����      C  , ,���9�������9�����������������������9����      C  , ,�������D���������������������D�������D      C  , ,�������D���������������������D�������D      C  , ,�������D�����������o�������o���D�������D      C  , ,������D����������S�������S���D������D      C  , ,�������D�����������7�������7���D�������D      C  , ,���q���D���q�����������������D���q���D      C  , ,���U���D���U�������������������D���U���D      C  , ,���9���D���9�������������������D���9���D      C  , ,���������������V������V���������������      C  , ,���������������V������V���������������      C  , ,������t��������������������t������t      C  , ,�������t�������������������t�������t      C  , ,�������t�������������������t�������t      C  , ,�������t����������o������o���t�������t      C  , ,������t���������S������S���t������t      C  , ,�������t����������7������7���t�������t      C  , ,���q���t���q���������������t���q���t      C  , ,���U���t���U�����������������t���U���t      C  , ,���9���t���9�����������������t���9���t      C  , ,���������������G���e���G���e������������      C  , ,���������������G���I���G���I������������      C  , ,���������������G���-���G���-������������      C  , ,���g�������g���G������G����������g����      C  , ,���K�������K���G�������G�����������K����      C  , ,���/�������/���G�������G�����������/����      C  , ,�������������G�������G���������������      C  , ,���������������G��á���G��á������������      C  , ,���������������G��ƅ���G��ƅ������������      C  , ,��ȿ������ȿ���G���i���G���i������ȿ����      C  , ,���-������-����������������������-���      C  , ,����������������������������������      C  , ,�������������������������������������      C  , ,�������������������������������������      C  , ,������������������g�������g����������      C  , ,������������������K�������K����������      C  , ,������������������/�������/����������      C  , ,���i������i��������������������i���      C  , ,���M������M����������������������M���      C  , ,���-���|���-���&�������&�������|���-���|      C  , ,������|������&�������&�������|������|      C  , ,�������|�������&�������&�������|�������|      C  , ,�������|�������&�������&�������|�������|      C  , ,�������|�������&���g���&���g���|�������|      C  , ,�������|�������&���K���&���K���|�������|      C  , ,�������|�������&���/���&���/���|�������|      C  , ,���i���|���i���&������&������|���i���|      C  , ,���M���|���M���&�������&�������|���M���|      C  , ,���������������G�������G����������������      C  , ,���+�������+���G�������G�����������+����      C  , ,�������������G�������G���������������      C  , ,�������������G���)���G���)�����������      C  , ,���������������G���a���G���a������������      C  , ,���E���|���E���&�������&�������|���E���|      C  , ,���E������E����������������������E���      C  , ,���)������)����������������������)���      C  , ,���)���|���)���&�������&�������|���)���|      C  , ,������|������&�������&�������|������|      C  , ,�������|�������&�������&�������|�������|      C  , ,�������|�������&������&������|�������|      C  , ,�������|�������&���c���&���c���|�������|      C  , ,�������|�������&���G���&���G���|�������|      C  , ,�������|�������&���+���&���+���|�������|      C  , ,���e���|���e���&������&������|���e���|      C  , ,���I���|���I���&�������&�������|���I���|      C  , ,����������������������������������      C  , ,�������������������������������������      C  , ,�����������������������������������      C  , ,������������������c�������c����������      C  , ,������������������G�������G����������      C  , ,������������������+�������+����������      C  , ,���e������e��������������������e���      C  , ,���I������I����������������������I���      C  , ,���������������G�������G����������������      C  , ,���c�������c���G������G����������c����      C  , ,���G�������G���G�������G�����������G����      C  , ,���������������G���E���G���E������������      C  , ,���I���D���I�������������������D���I���D      C  , ,���E���D���E�������������������D���E���D      C  , ,���)���D���)�������������������D���)���D      C  , ,������D����������������������D������D      C  , ,�������D�����������������������D�������D      C  , ,�������D���������������������D�������D      C  , ,�������D�����������c�������c���D�������D      C  , ,�������D�����������G�������G���D�������D      C  , ,�������D�����������+�������+���D�������D      C  , ,���e���D���e�����������������D���e���D      C  , ,���E�������E�����������������������E����      C  , ,���)�������)�����������������������)����      C  , ,�������������������������������������      C  , ,����������������������������������������      C  , ,��������������������������������������      C  , ,�������������������c�������c������������      C  , ,�������������������G�������G������������      C  , ,�������������������+�������+������������      C  , ,���E�������E���V�������V�����������E����      C  , ,���E���t���E�����������������t���E���t      C  , ,���)���t���)�����������������t���)���t      C  , ,������t��������������������t������t      C  , ,�������t���������������������t�������t      C  , ,�������t�������������������t�������t      C  , ,�������t����������c������c���t�������t      C  , ,�������t����������G������G���t�������t      C  , ,�������t����������+������+���t�������t      C  , ,���e���t���e���������������t���e���t      C  , ,���I���t���I�����������������t���I���t      C  , ,���)�������)���V�������V�����������)����      C  , ,�������������V�������V���������������      C  , ,���������������V�������V����������������      C  , ,���������������V������V���������������      C  , ,���������������V���c���V���c������������      C  , ,���������������V���G���V���G������������      C  , ,���������������V���+���V���+������������      C  , ,���e�������e���V������V����������e����      C  , ,���I�������I���V�������V�����������I����      C  , ,���e�������e���������������������e����      C  , ,���I�������I�����������������������I����      C  , ,�������D�����������/�������/���D�������D      C  , ,���i���D���i�����������������D���i���D      C  , ,���M���D���M�������������������D���M���D      C  , ,���-���D���-�������������������D���-���D      C  , ,������D����������������������D������D      C  , ,���-�������-�����������������������-����      C  , ,�������������������������������������      C  , ,���-���t���-�����������������t���-���t      C  , ,������t��������������������t������t      C  , ,�������t���������������������t�������t      C  , ,�������t���������������������t�������t      C  , ,�������t����������g������g���t�������t      C  , ,�������t����������K������K���t�������t      C  , ,�������t����������/������/���t�������t      C  , ,���i���t���i���������������t���i���t      C  , ,���M���t���M�����������������t���M���t      C  , ,����������������������������������������      C  , ,����������������������������������������      C  , ,�������������������g�������g������������      C  , ,�������������������K�������K������������      C  , ,�������������������/�������/������������      C  , ,���i�������i���������������������i����      C  , ,���M�������M�����������������������M����      C  , ,�������D�����������������������D�������D      C  , ,�������D�����������������������D�������D      C  , ,���-�������-���V�������V�����������-����      C  , ,�������������V�������V���������������      C  , ,���������������V�������V����������������      C  , ,���������������V�������V����������������      C  , ,���������������V���g���V���g������������      C  , ,���������������V���K���V���K������������      C  , ,���������������V���/���V���/������������      C  , ,���i�������i���V������V����������i����      C  , ,���M�������M���V�������V�����������M����      C  , ,�������D�����������g�������g���D�������D      C  , ,�������D�����������K�������K���D�������D      C  , ,���E�������E���~�������~�����������E����      C  , ,���)�������)���~�������~�����������)����      C  , ,�������������~�������~���������������      C  , ,���������������~�������~����������������      C  , ,���������������~������~���������������      C  , ,���������������~���c���~���c������������      C  , ,���������������~���G���~���G������������      C  , ,���������������~���+���~���+������������      C  , ,���e�������e���~������~����������e����      C  , ,���I�������I���~�������~�����������I����      C  , ,���-�������-���~�������~�����������-����      C  , ,�������������~�������~���������������      C  , ,���������������~�������~����������������      C  , ,���������������~�������~����������������      C  , ,���������������~���g���~���g������������      C  , ,���������������~���K���~���K������������      C  , ,���������������~���/���~���/������������      C  , ,���i�������i���~������~����������i����      C  , ,���M�������M���~�������~�����������M����      C  , ,������<����������������������<������<      C  , ,�������<�����������������������<�������<      C  , ,�������<�����������������������<�������<      C  , ,�������<�����������g�������g���<�������<      C  , ,�������<�����������K�������K���<�������<      C  , ,�������<�����������/�������/���<�������<      C  , ,���i���<���i�����������������<���i���<      C  , ,���M���<���M�������������������<���M���<      C  , ,���-������-����������������������-���      C  , ,����������������������������������      C  , ,�������������������������������������      C  , ,�������������������������������������      C  , ,������������������g�������g����������      C  , ,������������������K�������K����������      C  , ,������������������/�������/����������      C  , ,���i������i��������������������i���      C  , ,���M������M����������������������M���      C  , ,���-������-���N�������N����������-���      C  , ,������������N�������N�������������      C  , ,��������������N�������N��������������      C  , ,��������������N�������N��������������      C  , ,��������������N���g���N���g����������      C  , ,��������������N���K���N���K����������      C  , ,��������������N���/���N���/����������      C  , ,���i������i���N������N���������i���      C  , ,���M������M���N�������N����������M���      C  , ,���-���<���-�������������������<���-���<      C  , ,���I���<���I�������������������<���I���<      C  , ,���E������E���N�������N����������E���      C  , ,���)������)���N�������N����������)���      C  , ,������������N�������N�������������      C  , ,��������������N�������N��������������      C  , ,��������������N������N�������������      C  , ,��������������N���c���N���c����������      C  , ,��������������N���G���N���G����������      C  , ,��������������N���+���N���+����������      C  , ,���e������e���N������N���������e���      C  , ,���I������I���N�������N����������I���      C  , ,���)������)����������������������)���      C  , ,����������������������������������      C  , ,�������������������������������������      C  , ,�����������������������������������      C  , ,������������������c�������c����������      C  , ,������������������G�������G����������      C  , ,������������������+�������+����������      C  , ,���e������e��������������������e���      C  , ,���I������I����������������������I���      C  , ,���E���<���E�������������������<���E���<      C  , ,���)���<���)�������������������<���)���<      C  , ,������<����������������������<������<      C  , ,�������<�����������������������<�������<      C  , ,�������<���������������������<�������<      C  , ,�������<�����������c�������c���<�������<      C  , ,�������<�����������G�������G���<�������<      C  , ,�������<�����������+�������+���<�������<      C  , ,���e���<���e�����������������<���e���<      C  , ,���E������E����������������������E���      C  , ,���)���l���)�����������������l���)���l      C  , ,������l��������������������l������l      C  , ,�������l���������������������l�������l      C  , ,�������l�������������������l�������l      C  , ,�������l����������c������c���l�������l      C  , ,�������l����������G������G���l�������l      C  , ,�������l����������+������+���l�������l      C  , ,���e���l���e���������������l���e���l      C  , ,���I���l���I�����������������l���I���l      C  , ,���E������E��������������������E���      C  , ,���)������)��������������������)���      C  , ,��������������������������������      C  , ,�����������������������������������      C  , ,���������������������������������      C  , ,�����������������c������c����������      C  , ,�����������������G������G����������      C  , ,�����������������+������+����������      C  , ,���e������e������������������e���      C  , ,���I������I��������������������I���      C  , ,������������������a������a������������      C  , ,������������������E������E������������      C  , ,����������������)������)�����������      C  , ,���c�������c�������������������c����      C  , ,���G�������G���������������������G����      C  , ,���+�������+���������������������+����      C  , ,�����������������������������������      C  , ,��������������������������������������      C  , ,��������������������������������������      C  , ,���E���l���E�����������������l���E���l      C  , ,��������������������������������      C  , ,�����������������������������������      C  , ,�����������������������������������      C  , ,�����������������g������g����������      C  , ,�����������������K������K����������      C  , ,�����������������/������/����������      C  , ,���i������i������������������i���      C  , ,���M������M��������������������M���      C  , ,������l��������������������l������l      C  , ,�������l���������������������l�������l      C  , ,�������l���������������������l�������l      C  , ,�������l����������g������g���l�������l      C  , ,�������l����������K������K���l�������l      C  , ,�������l����������/������/���l�������l      C  , ,���i���l���i���������������l���i���l      C  , ,���M���l���M�����������������l���M���l      C  , ,���-���l���-�����������������l���-���l      C  , ,������������������e������e������������      C  , ,������������������I������I������������      C  , ,������������������-������-������������      C  , ,���g�������g�������������������g����      C  , ,���K�������K���������������������K����      C  , ,���/�������/���������������������/����      C  , ,�����������������������������������      C  , ,�����������������á�����á������������      C  , ,�����������������ƅ�����ƅ������������      C  , ,��ȿ������ȿ������i������i������ȿ����      C  , ,���-������-��������������������-���      C  , ,�������������~��Ϳ���~��Ϳ�����������      C  , ,���������������~��У���~��У������������      C  , ,���������������~��Ӈ���~��Ӈ������������      C  , ,���������������~���k���~���k������������      C  , ,��إ������إ���~���O���~���O������إ����      C  , ,��ۉ������ۉ���~���3���~���3������ۉ����      C  , ,���m�������m���~������~����������m����      C  , ,���Q�������Q���~�������~�����������Q����      C  , ,���5�������5���~�������~�����������5����      C  , ,�������������~�������~���������������      C  , ,���������������~������~���������������      C  , ,���������������~������~���������������      C  , ,���������������~���o���~���o������������      C  , ,�������������~���S���~���S�����������      C  , ,���������������~���7���~���7������������      C  , ,���q�������q���~������~����������q����      C  , ,���U�������U���~�������~�����������U����      C  , ,���9�������9���~�������~�����������9����      C  , ,���5������5����������������������5���      C  , ,���5���l���5�����������������l���5���l      C  , ,���5���<���5�������������������<���5���<      C  , ,���5������5��������������������5���      C  , ,���5������5���N�������N����������5���      C  , ,���1�������1���~�������~�����������1����      C  , ,������������������7�������7����������      C  , ,���q������q��������������������q���      C  , ,���U������U����������������������U���      C  , ,���9������9����������������������9���      C  , ,����������������������������������      C  , ,�����������������������������������      C  , ,������<����������������������<������<      C  , ,�������<���������������������<�������<      C  , ,�������<���������������������<�������<      C  , ,�������<�����������o�������o���<�������<      C  , ,������<����������S�������S���<������<      C  , ,�������<�����������7�������7���<�������<      C  , ,���q���<���q�����������������<���q���<      C  , ,���U���<���U�������������������<���U���<      C  , ,���9���<���9�������������������<���9���<      C  , ,�����������������������������������      C  , ,������������������o�������o����������      C  , ,������������N�������N�������������      C  , ,��������������N������N�������������      C  , ,��������������N������N�������������      C  , ,��������������N���o���N���o����������      C  , ,������������N���S���N���S���������      C  , ,��������������N���7���N���7����������      C  , ,���q������q���N������N���������q���      C  , ,���U������U���N�������N����������U���      C  , ,���9������9���N�������N����������9���      C  , ,����������������S�������S���������      C  , ,��ۉ�����ۉ�������3�������3�����ۉ���      C  , ,���m������m��������������������m���      C  , ,���Q������Q����������������������Q���      C  , ,���1������1����������������������1���      C  , ,���������������Ϳ������Ϳ���������      C  , ,���1���<���1�������������������<���1���<      C  , ,������<���������Ϳ������Ϳ���<������<      C  , ,���1������1���N�������N����������1���      C  , ,������������N��Ϳ���N��Ϳ���������      C  , ,��������������N��У���N��У����������      C  , ,��������������N��Ӈ���N��Ӈ����������      C  , ,��������������N���k���N���k����������      C  , ,��إ�����إ���N���O���N���O�����إ���      C  , ,��ۉ�����ۉ���N���3���N���3�����ۉ���      C  , ,���m������m���N������N���������m���      C  , ,���Q������Q���N�������N����������Q���      C  , ,�������<����������У������У���<�������<      C  , ,�������<����������Ӈ������Ӈ���<�������<      C  , ,�������<�����������k�������k���<�������<      C  , ,��إ���<��إ�������O�������O���<��إ���<      C  , ,��ۉ���<��ۉ�������3�������3���<��ۉ���<      C  , ,���m���<���m�����������������<���m���<      C  , ,���Q���<���Q�������������������<���Q���<      C  , ,�����������������У������У����������      C  , ,�����������������Ӈ������Ӈ����������      C  , ,������������������k�������k����������      C  , ,��إ�����إ�������O�������O�����إ���      C  , ,��إ���l��إ������O������O���l��إ���l      C  , ,��ۉ���l��ۉ������3������3���l��ۉ���l      C  , ,���m���l���m���������������l���m���l      C  , ,���Q���l���Q�����������������l���Q���l      C  , ,���1���l���1�����������������l���1���l      C  , ,������l��������Ϳ�����Ϳ���l������l      C  , ,���1������1��������������������1���      C  , ,��������������Ϳ�����Ϳ���������      C  , ,����������������У�����У����������      C  , ,����������������Ӈ�����Ӈ����������      C  , ,�����������������k������k����������      C  , ,��إ�����إ������O������O�����إ���      C  , ,��ۉ�����ۉ������3������3�����ۉ���      C  , ,���m������m������������������m���      C  , ,���Q������Q��������������������Q���      C  , ,�������l���������У�����У���l�������l      C  , ,�������l���������Ӈ�����Ӈ���l�������l      C  , ,��ˣ������ˣ������M������M������ˣ����      C  , ,��·������·������1������1������·����      C  , ,���k�������k�������������������k����      C  , ,���O�������O���������������������O����      C  , ,���3�������3���������������������3����      C  , ,�����������������������������������      C  , ,�����������������ݥ�����ݥ������������      C  , ,��������������������������������������      C  , ,������������������m������m������������      C  , ,�������l����������k������k���l�������l      C  , ,���������������������������������      C  , ,�����������������o������o����������      C  , ,���������������S������S���������      C  , ,�����������������7������7����������      C  , ,���q������q������������������q���      C  , ,���U������U��������������������U���      C  , ,���9������9��������������������9���      C  , ,�������l�������������������l�������l      C  , ,�������l����������o������o���l�������l      C  , ,������l���������S������S���l������l      C  , ,�������l����������7������7���l�������l      C  , ,���q���l���q���������������l���q���l      C  , ,���U���l���U�����������������l���U���l      C  , ,���9���l���9�����������������l���9���l      C  , ,������l��������������������l������l      C  , ,�������l�������������������l�������l      C  , ,��������������������������������      C  , ,����������������Q������Q�����������      C  , ,����������������5������5�����������      C  , ,���o�������o�������������������o����      C  , ,���S�������S���������������������S����      C  , ,���7�������7���������������������7����      C  , ,�����������������������������������      C  , ,��������������������������������������      C  , ,��������������������������������������      C  , ,������������������q������q������������      C  , ,���������������������������������      C  , ,  S����  S���G  T)���G  T)����  S����      C  , ,  Vc����  Vc���G  W���G  W����  Vc����      C  , ,  YG����  YG���G  Y����G  Y�����  YG����      C  , ,  \+����  \+���G  \����G  \�����  \+����      C  , ,  _����  _���G  _����G  _�����  _����      C  , ,  a�����  a����G  b����G  b�����  a�����      C  , ,  d�����  d����G  e����G  e�����  d�����      C  , ,  g�����  g����G  he���G  he����  g�����      C  , ,  j�����  j����G  kI���G  kI����  j�����      C  , ,  R���  R����  R�����  R����  R���      C  , ,  T����  T�����  U�����  U����  T����      C  , ,  W����  W�����  X����  X���  W����      C  , ,  Z����  Z�����  [c����  [c���  Z����      C  , ,  ]����  ]�����  ^G����  ^G���  ]����      C  , ,  `����  `�����  a+����  a+���  `����      C  , ,  ce���  ce����  d����  d���  ce���      C  , ,  fI���  fI����  f�����  f����  fI���      C  , ,  i-���  i-����  i�����  i����  i-���      C  , ,  l���  l����  l�����  l����  l���      C  , ,  R���|  R���&  R����&  R����|  R���|      C  , ,  T����|  T����&  U����&  U����|  T����|      C  , ,  W����|  W����&  X���&  X���|  W����|      C  , ,  Z����|  Z����&  [c���&  [c���|  Z����|      C  , ,  ]����|  ]����&  ^G���&  ^G���|  ]����|      C  , ,  `����|  `����&  a+���&  a+���|  `����|      C  , ,  ce���|  ce���&  d���&  d���|  ce���|      C  , ,  fI���|  fI���&  f����&  f����|  fI���|      C  , ,  i-���|  i-���&  i����&  i����|  i-���|      C  , ,  l���|  l���&  l����&  l����|  l���|      C  , ,  6�����  6����G  7A���G  7A����  6�����      C  , ,  9{����  9{���G  :%���G  :%����  9{����      C  , ,  <_����  <_���G  =	���G  =	����  <_����      C  , ,  ?C����  ?C���G  ?����G  ?�����  ?C����      C  , ,  B'����  B'���G  B����G  B�����  B'����      C  , ,  E����  E���G  E����G  E�����  E����      C  , ,  G�����  G����G  H����G  H�����  G�����      C  , ,  J�����  J����G  K}���G  K}����  J�����      C  , ,  M�����  M����G  Na���G  Na����  M�����      C  , ,  8	���|  8	���&  8����&  8����|  8	���|      C  , ,  :����|  :����&  ;����&  ;����|  :����|      C  , ,  =����|  =����&  >{���&  >{���|  =����|      C  , ,  @����|  @����&  A_���&  A_���|  @����|      C  , ,  C����|  C����&  DC���&  DC���|  C����|      C  , ,  F}���|  F}���&  G'���&  G'���|  F}���|      C  , ,  Ia���|  Ia���&  J���&  J���|  Ia���|      C  , ,  LE���|  LE���&  L����&  L����|  LE���|      C  , ,  O)���|  O)���&  O����&  O����|  O)���|      C  , ,  8	���  8	����  8�����  8����  8	���      C  , ,  :����  :�����  ;�����  ;����  :����      C  , ,  =����  =�����  >{����  >{���  =����      C  , ,  @����  @�����  A_����  A_���  @����      C  , ,  C����  C�����  DC����  DC���  C����      C  , ,  F}���  F}����  G'����  G'���  F}���      C  , ,  Ia���  Ia����  J����  J���  Ia���      C  , ,  LE���  LE����  L�����  L����  LE���      C  , ,  O)���  O)����  O�����  O����  O)���      C  , ,  P�����  P����G  QE���G  QE����  P�����      C  , ,  :�����  :�����  ;�����  ;�����  :�����      C  , ,  =�����  =�����  >{����  >{����  =�����      C  , ,  @�����  @�����  A_����  A_����  @�����      C  , ,  C�����  C�����  DC����  DC����  C�����      C  , ,  F}����  F}����  G'����  G'����  F}����      C  , ,  Ia����  Ia����  J����  J����  Ia����      C  , ,  LE����  LE����  L�����  L�����  LE����      C  , ,  O)����  O)����  O�����  O�����  O)����      C  , ,  =�����  =����V  >{���V  >{����  =�����      C  , ,  @�����  @����V  A_���V  A_����  @�����      C  , ,  C�����  C����V  DC���V  DC����  C�����      C  , ,  F}����  F}���V  G'���V  G'����  F}����      C  , ,  Ia����  Ia���V  J���V  J����  Ia����      C  , ,  LE����  LE���V  L����V  L�����  LE����      C  , ,  O)����  O)���V  O����V  O�����  O)����      C  , ,  8	����  8	���V  8����V  8�����  8	����      C  , ,  8	���D  8	����  8�����  8����D  8	���D      C  , ,  :����D  :�����  ;�����  ;����D  :����D      C  , ,  =����D  =�����  >{����  >{���D  =����D      C  , ,  @����D  @�����  A_����  A_���D  @����D      C  , ,  C����D  C�����  DC����  DC���D  C����D      C  , ,  F}���D  F}����  G'����  G'���D  F}���D      C  , ,  Ia���D  Ia����  J����  J���D  Ia���D      C  , ,  LE���D  LE����  L�����  L����D  LE���D      C  , ,  O)���D  O)����  O�����  O����D  O)���D      C  , ,  :�����  :����V  ;����V  ;�����  :�����      C  , ,  8	����  8	����  8�����  8�����  8	����      C  , ,  8	���t  8	���  8����  8����t  8	���t      C  , ,  :����t  :����  ;����  ;����t  :����t      C  , ,  =����t  =����  >{���  >{���t  =����t      C  , ,  @����t  @����  A_���  A_���t  @����t      C  , ,  C����t  C����  DC���  DC���t  C����t      C  , ,  F}���t  F}���  G'���  G'���t  F}���t      C  , ,  Ia���t  Ia���  J���  J���t  Ia���t      C  , ,  LE���t  LE���  L����  L����t  LE���t      C  , ,  O)���t  O)���  O����  O����t  O)���t      C  , ,  i-����  i-����  i�����  i�����  i-����      C  , ,  l����  l����  l�����  l�����  l����      C  , ,  ce����  ce���V  d���V  d����  ce����      C  , ,  fI����  fI���V  f����V  f�����  fI����      C  , ,  R���D  R����  R�����  R����D  R���D      C  , ,  T����D  T�����  U�����  U����D  T����D      C  , ,  W����D  W�����  X����  X���D  W����D      C  , ,  Z����D  Z�����  [c����  [c���D  Z����D      C  , ,  ]����D  ]�����  ^G����  ^G���D  ]����D      C  , ,  `����D  `�����  a+����  a+���D  `����D      C  , ,  ce���D  ce����  d����  d���D  ce���D      C  , ,  fI���D  fI����  f�����  f����D  fI���D      C  , ,  i-���D  i-����  i�����  i����D  i-���D      C  , ,  l���D  l����  l�����  l����D  l���D      C  , ,  i-����  i-���V  i����V  i�����  i-����      C  , ,  l����  l���V  l����V  l�����  l����      C  , ,  R����  R���V  R����V  R�����  R����      C  , ,  T�����  T����V  U����V  U�����  T�����      C  , ,  W�����  W����V  X���V  X����  W�����      C  , ,  Z�����  Z����V  [c���V  [c����  Z�����      C  , ,  ]�����  ]����V  ^G���V  ^G����  ]�����      C  , ,  `�����  `����V  a+���V  a+����  `�����      C  , ,  R����  R����  R�����  R�����  R����      C  , ,  T�����  T�����  U�����  U�����  T�����      C  , ,  W�����  W�����  X����  X����  W�����      C  , ,  Z�����  Z�����  [c����  [c����  Z�����      C  , ,  ]�����  ]�����  ^G����  ^G����  ]�����      C  , ,  `�����  `�����  a+����  a+����  `�����      C  , ,  ce����  ce����  d����  d����  ce����      C  , ,  fI����  fI����  f�����  f�����  fI����      C  , ,  R���t  R���  R����  R����t  R���t      C  , ,  T����t  T����  U����  U����t  T����t      C  , ,  W����t  W����  X���  X���t  W����t      C  , ,  Z����t  Z����  [c���  [c���t  Z����t      C  , ,  ]����t  ]����  ^G���  ^G���t  ]����t      C  , ,  `����t  `����  a+���  a+���t  `����t      C  , ,  ce���t  ce���  d���  d���t  ce���t      C  , ,  fI���t  fI���  f����  f����t  fI���t      C  , ,  i-���t  i-���  i����  i����t  i-���t      C  , ,  l���t  l���  l����  l����t  l���t      C  , ,  !����  !����  �����  �����  !����      C  , ,  !���D  !����  �����  ����D  !���D      C  , ,  !���|  !���&  ����&  ����|  !���|      C  , ,  !���t  !���  ����  ����t  !���t      C  , ,  !���  !����  �����  ����  !���      C  , ,  !����  !���V  ����V  �����  !����      C  , ,  &����|  &����&  '[���&  '[���|  &����|      C  , ,  )����|  )����&  *?���&  *?���|  )����|      C  , ,  ,y���|  ,y���&  -#���&  -#���|  ,y���|      C  , ,  /]���|  /]���&  0���&  0���|  /]���|      C  , ,  2A���|  2A���&  2����&  2����|  2A���|      C  , ,  5%���|  5%���&  5����&  5����|  5%���|      C  , ,  �����  ����G  =���G  =����  �����      C  , ,  w����  w���G   !���G   !����  w����      C  , ,  "[����  "[���G  #���G  #����  "[����      C  , ,  %?����  %?���G  %����G  %�����  %?����      C  , ,  (#����  (#���G  (����G  (�����  (#����      C  , ,  +����  +���G  +����G  +�����  +����      C  , ,  -�����  -����G  .����G  .�����  -�����      C  , ,  0�����  0����G  1y���G  1y����  0�����      C  , ,  3�����  3����G  4]���G  4]����  3�����      C  , ,  ���|  ���&  ����&  ����|  ���|      C  , ,   ����|   ����&  !����&  !����|   ����|      C  , ,  ���  ����  �����  ����  ���      C  , ,   ����   �����  !�����  !����   ����      C  , ,  #����  #�����  $w����  $w���  #����      C  , ,  &����  &�����  '[����  '[���  &����      C  , ,  )����  )�����  *?����  *?���  )����      C  , ,  ,y���  ,y����  -#����  -#���  ,y���      C  , ,  /]���  /]����  0����  0���  /]���      C  , ,  2A���  2A����  2�����  2����  2A���      C  , ,  5%���  5%����  5�����  5����  5%���      C  , ,  #����|  #����&  $w���&  $w���|  #����|      C  , ,  Y���|  Y���&  ���&  ���|  Y���|      C  , ,  =���|  =���&  ����&  ����|  =���|      C  , ,  �����  ����G  9���G  9����  �����      C  , ,  ���|  ���&  ����&  ����|  ���|      C  , ,  ���  ����  �����  ����  ���      C  , ,  ���|  ���&  ����&  ����|  ���|      C  , ,  ���  ����  �����  ����  ���      C  , ,  ����  �����  �����  ����  ����      C  , ,  s����  s���G  ���G  ����  s����      C  , ,  W����  W���G  	���G  	����  W����      C  , ,  	����  	�����  
s����  
s���  	����      C  , ,  ����  �����  W����  W���  ����      C  , ,  ����  �����  ;����  ;���  ����      C  , ,  u���  u����  ����  ���  u���      C  , ,  Y���  Y����  ����  ���  Y���      C  , ,  =���  =����  �����  ����  =���      C  , ,  ;����  ;���G  ����G  �����  ;����      C  , ,  ����  ���G  ����G  �����  ����      C  , ,  ����  ���G  ����G  �����  ����      C  , ,  ����|  ����&  ����&  ����|  ����|      C  , ,  	����|  	����&  
s���&  
s���|  	����|      C  , ,  �����  ����G  ����G  �����  �����      C  , ,  �����  ����G  u���G  u����  �����      C  , ,  �����  ����G  Y���G  Y����  �����      C  , ,  ����|  ����&  W���&  W���|  ����|      C  , ,  ����|  ����&  ;���&  ;���|  ����|      C  , ,  u���|  u���&  ���&  ���|  u���|      C  , ,  �����  ����V  ;���V  ;����  �����      C  , ,  u����  u���V  ���V  ����  u����      C  , ,  Y����  Y���V  ���V  ����  Y����      C  , ,  =����  =���V  ����V  �����  =����      C  , ,  �����  ����V  ����V  �����  �����      C  , ,  ����D  �����  �����  ����D  ����D      C  , ,  	����D  	�����  
s����  
s���D  	����D      C  , ,  ����  ���V  ����V  �����  ����      C  , ,  ���t  ���  ����  ����t  ���t      C  , ,  ���t  ���  ����  ����t  ���t      C  , ,  ����t  ����  ����  ����t  ����t      C  , ,  	����t  	����  
s���  
s���t  	����t      C  , ,  ����t  ����  W���  W���t  ����t      C  , ,  ����t  ����  ;���  ;���t  ����t      C  , ,  u���t  u���  ���  ���t  u���t      C  , ,  Y���t  Y���  ���  ���t  Y���t      C  , ,  =���t  =���  ����  ����t  =���t      C  , ,  ����D  �����  W����  W���D  ����D      C  , ,  ����D  �����  ;����  ;���D  ����D      C  , ,  u���D  u����  ����  ���D  u���D      C  , ,  Y���D  Y����  ����  ���D  Y���D      C  , ,  =���D  =����  �����  ����D  =���D      C  , ,  ���D  ����  �����  ����D  ���D      C  , ,  ���D  ����  �����  ����D  ���D      C  , ,  	�����  	����V  
s���V  
s����  	�����      C  , ,  ����  ����  �����  �����  ����      C  , ,  ����  ����  �����  �����  ����      C  , ,  �����  �����  �����  �����  �����      C  , ,  	�����  	�����  
s����  
s����  	�����      C  , ,  �����  �����  W����  W����  �����      C  , ,  �����  �����  ;����  ;����  �����      C  , ,  u����  u����  ����  ����  u����      C  , ,  Y����  Y����  ����  ����  Y����      C  , ,  =����  =����  �����  �����  =����      C  , ,  �����  ����V  W���V  W����  �����      C  , ,  ����  ���V  ����V  �����  ����      C  , ,  #����D  #�����  $w����  $w���D  #����D      C  , ,  &����D  &�����  '[����  '[���D  &����D      C  , ,  )����D  )�����  *?����  *?���D  )����D      C  , ,  ,y���D  ,y����  -#����  -#���D  ,y���D      C  , ,  /]���D  /]����  0����  0���D  /]���D      C  , ,  2A���D  2A����  2�����  2����D  2A���D      C  , ,  5%���D  5%����  5�����  5����D  5%���D      C  , ,  ���t  ���  ����  ����t  ���t      C  , ,   ����t   ����  !����  !����t   ����t      C  , ,  #����t  #����  $w���  $w���t  #����t      C  , ,  &����t  &����  '[���  '[���t  &����t      C  , ,  )����t  )����  *?���  *?���t  )����t      C  , ,  ,y���t  ,y���  -#���  -#���t  ,y���t      C  , ,  /]���t  /]���  0���  0���t  /]���t      C  , ,  2A���t  2A���  2����  2����t  2A���t      C  , ,  5%���t  5%���  5����  5����t  5%���t      C  , ,   �����   �����  !�����  !�����   �����      C  , ,  #�����  #�����  $w����  $w����  #�����      C  , ,  &�����  &�����  '[����  '[����  &�����      C  , ,  )�����  )�����  *?����  *?����  )�����      C  , ,  ,y����  ,y����  -#����  -#����  ,y����      C  , ,  /]����  /]����  0����  0����  /]����      C  , ,  2A����  2A����  2�����  2�����  2A����      C  , ,  5%����  5%����  5�����  5�����  5%����      C  , ,  5%����  5%���V  5����V  5�����  5%����      C  , ,  #�����  #����V  $w���V  $w����  #�����      C  , ,  &�����  &����V  '[���V  '[����  &�����      C  , ,  )�����  )����V  *?���V  *?����  )�����      C  , ,  ,y����  ,y���V  -#���V  -#����  ,y����      C  , ,  /]����  /]���V  0���V  0����  /]����      C  , ,  2A����  2A���V  2����V  2�����  2A����      C  , ,  ����  ����  �����  �����  ����      C  , ,  ���D  ����  �����  ����D  ���D      C  , ,  ����  ���V  ����V  �����  ����      C  , ,   �����   ����V  !����V  !�����   �����      C  , ,   ����D   �����  !�����  !����D   ����D      C  , ,  !���l  !���  ����  ����l  !���l      C  , ,  !���  !���N  ����N  ����  !���      C  , ,  ����  ���~  ����~  �����  ����      C  , ,  ����  ���~  ����~  �����  ����      C  , ,  �����  ����~  ����~  �����  �����      C  , ,  	�����  	����~  
s���~  
s����  	�����      C  , ,  �����  ����~  W���~  W����  �����      C  , ,  �����  ����~  ;���~  ;����  �����      C  , ,  u����  u���~  ���~  ����  u����      C  , ,  Y����  Y���~  ���~  ����  Y����      C  , ,  =����  =���~  ����~  �����  =����      C  , ,  !����  !���~  ����~  �����  !����      C  , ,  ����  ���~  ����~  �����  ����      C  , ,   �����   ����~  !����~  !�����   �����      C  , ,  #�����  #����~  $w���~  $w����  #�����      C  , ,  &�����  &����~  '[���~  '[����  &�����      C  , ,  )�����  )����~  *?���~  *?����  )�����      C  , ,  ,y����  ,y���~  -#���~  -#����  ,y����      C  , ,  /]����  /]���~  0���~  0����  /]����      C  , ,  2A����  2A���~  2����~  2�����  2A����      C  , ,  5%����  5%���~  5����~  5�����  5%����      C  , ,  !���  !���  ����  ����  !���      C  , ,  !���<  !����  �����  ����<  !���<      C  , ,  !���  !����  �����  ����  !���      C  , ,  )����  )����N  *?���N  *?���  )����      C  , ,  ,y���  ,y���N  -#���N  -#���  ,y���      C  , ,  /]���  /]���N  0���N  0���  /]���      C  , ,  2A���  2A���N  2����N  2����  2A���      C  , ,  5%���  5%���N  5����N  5����  5%���      C  , ,  ���  ���N  ����N  ����  ���      C  , ,   ����   ����N  !����N  !����   ����      C  , ,  #����  #����N  $w���N  $w���  #����      C  , ,  ���<  ����  �����  ����<  ���<      C  , ,   ����<   �����  !�����  !����<   ����<      C  , ,  #����<  #�����  $w����  $w���<  #����<      C  , ,  &����<  &�����  '[����  '[���<  &����<      C  , ,  )����<  )�����  *?����  *?���<  )����<      C  , ,  ,y���<  ,y����  -#����  -#���<  ,y���<      C  , ,  /]���<  /]����  0����  0���<  /]���<      C  , ,  2A���<  2A����  2�����  2����<  2A���<      C  , ,  5%���<  5%����  5�����  5����<  5%���<      C  , ,  &����  &����N  '[���N  '[���  &����      C  , ,  ���  ����  �����  ����  ���      C  , ,   ����   �����  !�����  !����   ����      C  , ,  #����  #�����  $w����  $w���  #����      C  , ,  &����  &�����  '[����  '[���  &����      C  , ,  )����  )�����  *?����  *?���  )����      C  , ,  ,y���  ,y����  -#����  -#���  ,y���      C  , ,  /]���  /]����  0����  0���  /]���      C  , ,  2A���  2A����  2�����  2����  2A���      C  , ,  5%���  5%����  5�����  5����  5%���      C  , ,  ����  ����N  ;���N  ;���  ����      C  , ,  u���  u���N  ���N  ���  u���      C  , ,  Y���  Y���N  ���N  ���  Y���      C  , ,  =���  =���N  ����N  ����  =���      C  , ,  ���  ���N  ����N  ����  ���      C  , ,  ���  ���N  ����N  ����  ���      C  , ,  ����  ����N  ����N  ����  ����      C  , ,  ���<  ����  �����  ����<  ���<      C  , ,  ���  ����  �����  ����  ���      C  , ,  ���  ����  �����  ����  ���      C  , ,  ����  �����  �����  ����  ����      C  , ,  	����  	�����  
s����  
s���  	����      C  , ,  ����  �����  W����  W���  ����      C  , ,  ����  �����  ;����  ;���  ����      C  , ,  u���  u����  ����  ���  u���      C  , ,  Y���  Y����  ����  ���  Y���      C  , ,  =���  =����  �����  ����  =���      C  , ,  ���<  ����  �����  ����<  ���<      C  , ,  ����<  �����  �����  ����<  ����<      C  , ,  	����<  	�����  
s����  
s���<  	����<      C  , ,  ����<  �����  W����  W���<  ����<      C  , ,  ����<  �����  ;����  ;���<  ����<      C  , ,  u���<  u����  ����  ���<  u���<      C  , ,  Y���<  Y����  ����  ���<  Y���<      C  , ,  =���<  =����  �����  ����<  =���<      C  , ,  	����  	����N  
s���N  
s���  	����      C  , ,  ����  ����N  W���N  W���  ����      C  , ,  u���l  u���  ���  ���l  u���l      C  , ,  Y���l  Y���  ���  ���l  Y���l      C  , ,  =���l  =���  ����  ����l  =���l      C  , ,  ���l  ���  ����  ����l  ���l      C  , ,  ���l  ���  ����  ����l  ���l      C  , ,  ����l  ����  ����  ����l  ����l      C  , ,  ���  ���  ����  ����  ���      C  , ,  ���  ���  ����  ����  ���      C  , ,  ����  ����  ����  ����  ����      C  , ,  	����  	����  
s���  
s���  	����      C  , ,  ����  ����  W���  W���  ����      C  , ,  ����  ����  ;���  ;���  ����      C  , ,  u���  u���  ���  ���  u���      C  , ,  Y���  Y���  ���  ���  Y���      C  , ,  =���  =���  ����  ����  =���      C  , ,  	����l  	����  
s���  
s���l  	����l      C  , ,  ����l  ����  W���  W���l  ����l      C  , ,  ����l  ����  ;���  ;���l  ����l      C  , ,  �����  ����  9���  9����  �����      C  , ,  s����  s���  ���  ����  s����      C  , ,  W����  W���  	���  	����  W����      C  , ,  ;����  ;���  ����  �����  ;����      C  , ,  ����  ���  ����  �����  ����      C  , ,  ����  ���  ����  �����  ����      C  , ,  �����  ����  ����  �����  �����      C  , ,  �����  ����  u���  u����  �����      C  , ,  �����  ����  Y���  Y����  �����      C  , ,  #����  #����  $w���  $w���  #����      C  , ,  &����  &����  '[���  '[���  &����      C  , ,  )����  )����  *?���  *?���  )����      C  , ,  ,y���  ,y���  -#���  -#���  ,y���      C  , ,  /]���  /]���  0���  0���  /]���      C  , ,  2A���  2A���  2����  2����  2A���      C  , ,  5%���  5%���  5����  5����  5%���      C  , ,  &����l  &����  '[���  '[���l  &����l      C  , ,  )����l  )����  *?���  *?���l  )����l      C  , ,  ,y���l  ,y���  -#���  -#���l  ,y���l      C  , ,  /]���l  /]���  0���  0���l  /]���l      C  , ,  2A���l  2A���  2����  2����l  2A���l      C  , ,  5%���l  5%���  5����  5����l  5%���l      C  , ,  ���l  ���  ����  ����l  ���l      C  , ,   ����l   ����  !����  !����l   ����l      C  , ,  #����l  #����  $w���  $w���l  #����l      C  , ,  ���  ���  ����  ����  ���      C  , ,   ����   ����  !����  !����   ����      C  , ,  �����  ����  =���  =����  �����      C  , ,  w����  w���   !���   !����  w����      C  , ,  "[����  "[���  #���  #����  "[����      C  , ,  %?����  %?���  %����  %�����  %?����      C  , ,  (#����  (#���  (����  (�����  (#����      C  , ,  +����  +���  +����  +�����  +����      C  , ,  -�����  -����  .����  .�����  -�����      C  , ,  0�����  0����  1y���  1y����  0�����      C  , ,  3�����  3����  4]���  4]����  3�����      C  , ,  l����  l���~  l����~  l�����  l����      C  , ,  8	����  8	���~  8����~  8�����  8	����      C  , ,  :�����  :����~  ;����~  ;�����  :�����      C  , ,  =�����  =����~  >{���~  >{����  =�����      C  , ,  @�����  @����~  A_���~  A_����  @�����      C  , ,  C�����  C����~  DC���~  DC����  C�����      C  , ,  F}����  F}���~  G'���~  G'����  F}����      C  , ,  Ia����  Ia���~  J���~  J����  Ia����      C  , ,  LE����  LE���~  L����~  L�����  LE����      C  , ,  O)����  O)���~  O����~  O�����  O)����      C  , ,  R����  R���~  R����~  R�����  R����      C  , ,  T�����  T����~  U����~  U�����  T�����      C  , ,  W�����  W����~  X���~  X����  W�����      C  , ,  Z�����  Z����~  [c���~  [c����  Z�����      C  , ,  ]�����  ]����~  ^G���~  ^G����  ]�����      C  , ,  `�����  `����~  a+���~  a+����  `�����      C  , ,  ce����  ce���~  d���~  d����  ce����      C  , ,  fI����  fI���~  f����~  f�����  fI����      C  , ,  i-����  i-���~  i����~  i�����  i-����      C  , ,  i-���  i-����  i�����  i����  i-���      C  , ,  l���  l����  l�����  l����  l���      C  , ,  R���<  R����  R�����  R����<  R���<      C  , ,  T����<  T�����  U�����  U����<  T����<      C  , ,  W����<  W�����  X����  X���<  W����<      C  , ,  Z����<  Z�����  [c����  [c���<  Z����<      C  , ,  ]����<  ]�����  ^G����  ^G���<  ]����<      C  , ,  `����<  `�����  a+����  a+���<  `����<      C  , ,  ce���<  ce����  d����  d���<  ce���<      C  , ,  fI���<  fI����  f�����  f����<  fI���<      C  , ,  i-���<  i-����  i�����  i����<  i-���<      C  , ,  l���<  l����  l�����  l����<  l���<      C  , ,  R���  R���N  R����N  R����  R���      C  , ,  T����  T����N  U����N  U����  T����      C  , ,  W����  W����N  X���N  X���  W����      C  , ,  Z����  Z����N  [c���N  [c���  Z����      C  , ,  ]����  ]����N  ^G���N  ^G���  ]����      C  , ,  `����  `����N  a+���N  a+���  `����      C  , ,  ce���  ce���N  d���N  d���  ce���      C  , ,  fI���  fI���N  f����N  f����  fI���      C  , ,  i-���  i-���N  i����N  i����  i-���      C  , ,  l���  l���N  l����N  l����  l���      C  , ,  R���  R����  R�����  R����  R���      C  , ,  T����  T�����  U�����  U����  T����      C  , ,  W����  W�����  X����  X���  W����      C  , ,  Z����  Z�����  [c����  [c���  Z����      C  , ,  ]����  ]�����  ^G����  ^G���  ]����      C  , ,  `����  `�����  a+����  a+���  `����      C  , ,  ce���  ce����  d����  d���  ce���      C  , ,  fI���  fI����  f�����  f����  fI���      C  , ,  =����  =�����  >{����  >{���  =����      C  , ,  @����  @�����  A_����  A_���  @����      C  , ,  C����  C�����  DC����  DC���  C����      C  , ,  F}���  F}����  G'����  G'���  F}���      C  , ,  Ia���  Ia����  J����  J���  Ia���      C  , ,  LE���  LE����  L�����  L����  LE���      C  , ,  O)���  O)����  O�����  O����  O)���      C  , ,  :����  :����N  ;����N  ;����  :����      C  , ,  =����  =����N  >{���N  >{���  =����      C  , ,  @����  @����N  A_���N  A_���  @����      C  , ,  C����  C����N  DC���N  DC���  C����      C  , ,  F}���  F}���N  G'���N  G'���  F}���      C  , ,  Ia���  Ia���N  J���N  J���  Ia���      C  , ,  LE���  LE���N  L����N  L����  LE���      C  , ,  O)���  O)���N  O����N  O����  O)���      C  , ,  8	���  8	���N  8����N  8����  8	���      C  , ,  8	���  8	����  8�����  8����  8	���      C  , ,  8	���<  8	����  8�����  8����<  8	���<      C  , ,  :����<  :�����  ;�����  ;����<  :����<      C  , ,  =����<  =�����  >{����  >{���<  =����<      C  , ,  @����<  @�����  A_����  A_���<  @����<      C  , ,  C����<  C�����  DC����  DC���<  C����<      C  , ,  F}���<  F}����  G'����  G'���<  F}���<      C  , ,  Ia���<  Ia����  J����  J���<  Ia���<      C  , ,  LE���<  LE����  L�����  L����<  LE���<      C  , ,  O)���<  O)����  O�����  O����<  O)���<      C  , ,  :����  :�����  ;�����  ;����  :����      C  , ,  :����  :����  ;����  ;����  :����      C  , ,  =����  =����  >{���  >{���  =����      C  , ,  @����  @����  A_���  A_���  @����      C  , ,  C����  C����  DC���  DC���  C����      C  , ,  F}���  F}���  G'���  G'���  F}���      C  , ,  Ia���  Ia���  J���  J���  Ia���      C  , ,  LE���  LE���  L����  L����  LE���      C  , ,  O)���  O)���  O����  O����  O)���      C  , ,  8	���  8	���  8����  8����  8	���      C  , ,  8	���l  8	���  8����  8����l  8	���l      C  , ,  :����l  :����  ;����  ;����l  :����l      C  , ,  =����l  =����  >{���  >{���l  =����l      C  , ,  @����l  @����  A_���  A_���l  @����l      C  , ,  C����l  C����  DC���  DC���l  C����l      C  , ,  F}���l  F}���  G'���  G'���l  F}���l      C  , ,  Ia���l  Ia���  J���  J���l  Ia���l      C  , ,  LE���l  LE���  L����  L����l  LE���l      C  , ,  O)���l  O)���  O����  O����l  O)���l      C  , ,  6�����  6����  7A���  7A����  6�����      C  , ,  9{����  9{���  :%���  :%����  9{����      C  , ,  <_����  <_���  =	���  =	����  <_����      C  , ,  ?C����  ?C���  ?����  ?�����  ?C����      C  , ,  B'����  B'���  B����  B�����  B'����      C  , ,  E����  E���  E����  E�����  E����      C  , ,  G�����  G����  H����  H�����  G�����      C  , ,  J�����  J����  K}���  K}����  J�����      C  , ,  M�����  M����  Na���  Na����  M�����      C  , ,  P�����  P����  QE���  QE����  P�����      C  , ,  ce���  ce���  d���  d���  ce���      C  , ,  fI���  fI���  f����  f����  fI���      C  , ,  R���l  R���  R����  R����l  R���l      C  , ,  T����l  T����  U����  U����l  T����l      C  , ,  W����l  W����  X���  X���l  W����l      C  , ,  Z����l  Z����  [c���  [c���l  Z����l      C  , ,  ]����l  ]����  ^G���  ^G���l  ]����l      C  , ,  `����l  `����  a+���  a+���l  `����l      C  , ,  ce���l  ce���  d���  d���l  ce���l      C  , ,  fI���l  fI���  f����  f����l  fI���l      C  , ,  i-���l  i-���  i����  i����l  i-���l      C  , ,  l���l  l���  l����  l����l  l���l      C  , ,  i-���  i-���  i����  i����  i-���      C  , ,  l���  l���  l����  l����  l���      C  , ,  R���  R���  R����  R����  R���      C  , ,  T����  T����  U����  U����  T����      C  , ,  W����  W����  X���  X���  W����      C  , ,  Z����  Z����  [c���  [c���  Z����      C  , ,  ]����  ]����  ^G���  ^G���  ]����      C  , ,  `����  `����  a+���  a+���  `����      C  , ,  S����  S���  T)���  T)����  S����      C  , ,  Vc����  Vc���  W���  W����  Vc����      C  , ,  YG����  YG���  Y����  Y�����  YG����      C  , ,  \+����  \+���  \����  \�����  \+����      C  , ,  _����  _���  _����  _�����  _����      C  , ,  a�����  a����  b����  b�����  a�����      C  , ,  d�����  d����  e����  e�����  d�����      C  , ,  g�����  g����  he���  he����  g�����      C  , ,  j�����  j����  kI���  kI����  j�����      D   ,���3  U���3  ;   �  ;   �  U���3  U      D   ,���3   ����3  �   �  �   �   ����3   �      D   ,���3������3���e   ����e   �������3���      D   ,���3�������3���   ����   ��������3����      D   ,  6  U  6  ;  7�  ;  7�  U  6  U      D   ,   �  !   �  �  �  �  �  !   �  !      D   ,  �  !  �  �  �  �  �  !  �  !      D   ,  �  !  �  �  �  �  �  !  �  !      D   ,  	�  !  	�  �  
�  �  
�  !  	�  !      D   ,  �  !  �  �  u  �  u  !  �  !      D   ,  s  !  s  �  Y  �  Y  !  s  !      D   ,  W  !  W  �  =  �  =  !  W  !      D   ,  ;  !  ;  �  !  �  !  !  ;  !      D   ,    !    �    �    !    !      D   ,    !    �  �  �  �  !    !      D   ,  �  !  �  �  �  �  �  !  �  !      D   ,   �  !   �  �  !�  �  !�  !   �  !      D   ,  #�  !  #�  �  $�  �  $�  !  #�  !      D   ,  &�  !  &�  �  'y  �  'y  !  &�  !      D   ,  )w  !  )w  �  *]  �  *]  !  )w  !      D   ,  ,[  !  ,[  �  -A  �  -A  !  ,[  !      D   ,  /?  !  /?  �  0%  �  0%  !  /?  !      D   ,  2#  !  2#  �  3	  �  3	  !  2#  !      D   ,  5  !  5  �  5�  �  5�  !  5  !      D   ,  7�  !  7�  �  8�  �  8�  !  7�  !      D   ,  :�  !  :�  �  ;�  �  ;�  !  :�  !      D   ,  =�  !  =�  �  >�  �  >�  !  =�  !      D   ,  @�  !  @�  �  A}  �  A}  !  @�  !      D   ,  C{  !  C{  �  Da  �  Da  !  C{  !      D   ,  F_  !  F_  �  GE  �  GE  !  F_  !      D   ,  IC  !  IC  �  J)  �  J)  !  IC  !      D   ,  L'  !  L'  �  M  �  M  !  L'  !      D   ,  O  !  O  �  O�  �  O�  !  O  !      D   ,  Q�  !  Q�  �  R�  �  R�  !  Q�  !      D   ,  T�  !  T�  �  U�  �  U�  !  T�  !      D   ,  W�  !  W�  �  X�  �  X�  !  W�  !      D   ,  Z�  !  Z�  �  [�  �  [�  !  Z�  !      D   ,  ]  !  ]  �  ^e  �  ^e  !  ]  !      D   ,  `c  !  `c  �  aI  �  aI  !  `c  !      D   ,  cG  !  cG  �  d-  �  d-  !  cG  !      D   ,  f+  !  f+  �  g  �  g  !  f+  !      D   ,  i  !  i  �  i�  �  i�  !  i  !      D   ,  k�  !  k�  �  l�  �  l�  !  k�  !      D   ,  6   �  6  �  7�  �  7�   �  6   �      D   ,  A�  U  A�  ;  CI  ;  CI  U  A�  U      D   ,  D�  U  D�  ;  F-  ;  F-  U  D�  U      D   ,  Gw  U  Gw  ;  I  ;  I  U  Gw  U      D   ,  J[  U  J[  ;  K�  ;  K�  U  J[  U      D   ,  M?  U  M?  ;  N�  ;  N�  U  M?  U      D   ,  P#  U  P#  ;  Q�  ;  Q�  U  P#  U      D   ,  S  U  S  ;  T�  ;  T�  U  S  U      D   ,  U�  U  U�  ;  W�  ;  W�  U  U�  U      D   ,  X�  U  X�  ;  Zi  ;  Zi  U  X�  U      D   ,  [�  U  [�  ;  ]M  ;  ]M  U  [�  U      D   ,  ^�  U  ^�  ;  `1  ;  `1  U  ^�  U      D   ,  a{  U  a{  ;  c  ;  c  U  a{  U      D   ,  d_  U  d_  ;  e�  ;  e�  U  d_  U      D   ,  gC  U  gC  ;  h�  ;  h�  U  gC  U      D   ,  j'  U  j'  ;  k�  ;  k�  U  j'  U      D   ,  9  U  9  ;  :�  ;  :�  U  9  U      D   ,  ;�  U  ;�  ;  =�  ;  =�  U  ;�  U      D   ,  >�  U  >�  ;  @e  ;  @e  U  >�  U      D   ,  0W  U  0W  ;  1�  ;  1�  U  0W  U      D   ,  3;  U  3;  ;  4�  ;  4�  U  3;  U      D   ,  
�  U  
�  ;  ]  ;  ]  U  
�  U      D   ,  �  U  �  ;  A  ;  A  U  �  U      D   ,  �  U  �  ;  %  ;  %  U  �  U      D   ,  o  U  o  ;  	  ;  	  U  o  U      D   ,  S  U  S  ;  �  ;  �  U  S  U      D   ,  7  U  7  ;  �  ;  �  U  7  U      D   ,    U    ;  �  ;  �  U    U      D   ,  �  U  �  ;   �  ;   �  U  �  U      D   ,  !�  U  !�  ;  #}  ;  #}  U  !�  U      D   ,  $�  U  $�  ;  &a  ;  &a  U  $�  U      D   ,  '�  U  '�  ;  )E  ;  )E  U  '�  U      D   ,  *�  U  *�  ;  ,)  ;  ,)  U  *�  U      D   ,    U    ;  �  ;  �  U    U      D   ,  -s  U  -s  ;  /  ;  /  U  -s  U      D   ,  �  U  �  ;  �  ;  �  U  �  U      D   ,  �  U  �  ;  	y  ;  	y  U  �  U      D   ,  
�   �  
�  �  ]  �  ]   �  
�   �      D   ,  �   �  �  �  A  �  A   �  �   �      D   ,  �   �  �  �  %  �  %   �  �   �      D   ,  o   �  o  �  	  �  	   �  o   �      D   ,  S   �  S  �  �  �  �   �  S   �      D   ,  7   �  7  �  �  �  �   �  7   �      D   ,     �    �  �  �  �   �     �      D   ,  �   �  �  �   �  �   �   �  �   �      D   ,  !�   �  !�  �  #}  �  #}   �  !�   �      D   ,  $�   �  $�  �  &a  �  &a   �  $�   �      D   ,  '�   �  '�  �  )E  �  )E   �  '�   �      D   ,  *�   �  *�  �  ,)  �  ,)   �  *�   �      D   ,  -s   �  -s  �  /  �  /   �  -s   �      D   ,  0W   �  0W  �  1�  �  1�   �  0W   �      D   ,  3;   �  3;  �  4�  �  4�   �  3;   �      D   ,     �    �  �  �  �   �     �      D   ,  �   �  �  �  �  �  �   �  �   �      D   ,  �   �  �  �  	y  �  	y   �  �   �      D   ,  >�   �  >�  �  @e  �  @e   �  >�   �      D   ,  A�   �  A�  �  CI  �  CI   �  A�   �      D   ,  D�   �  D�  �  F-  �  F-   �  D�   �      D   ,  Gw   �  Gw  �  I  �  I   �  Gw   �      D   ,  J[   �  J[  �  K�  �  K�   �  J[   �      D   ,  M?   �  M?  �  N�  �  N�   �  M?   �      D   ,  P#   �  P#  �  Q�  �  Q�   �  P#   �      D   ,  S   �  S  �  T�  �  T�   �  S   �      D   ,  U�   �  U�  �  W�  �  W�   �  U�   �      D   ,  X�   �  X�  �  Zi  �  Zi   �  X�   �      D   ,  [�   �  [�  �  ]M  �  ]M   �  [�   �      D   ,  ^�   �  ^�  �  `1  �  `1   �  ^�   �      D   ,  a{   �  a{  �  c  �  c   �  a{   �      D   ,  d_   �  d_  �  e�  �  e�   �  d_   �      D   ,  gC   �  gC  �  h�  �  h�   �  gC   �      D   ,  j'   �  j'  �  k�  �  k�   �  j'   �      D   ,  9   �  9  �  :�  �  :�   �  9   �      D   ,  ;�   �  ;�  �  =�  �  =�   �  ;�   �      D   ,���G  U���G  ;����  ;����  U���G  U      D   ,���'  !���'  ����  ����  !���'  !      D   ,���G   ����G  �����  �����   ����G   �      D   ,���  !���  �����  �����  !���  !      D   ,����  !����  �����  �����  !����  !      D   ,����  !����  �����  �����  !����  !      D   ,����  !����  �����  �����  !����  !      D   ,����  !����  �����  �����  !����  !      D   ,���  !���  ����e  ����e  !���  !      D   ,���c  !���c  ����I  ����I  !���c  !      D   ,���G  !���G  ����-  ����-  !���G  !      D   ,���+  !���+  ����  ����  !���+  !      D   ,���  !���  �����  �����  !���  !      D   ,����  !����  �����  �����  !����  !      D   ,����  !����  �����  �����  !����  !      D   ,����  !����  �����  �����  !����  !      D   ,����  !����  �����  �����  !����  !      D   ,����  !����  ����i  ����i  !����  !      D   ,���g  !���g  ����M  ����M  !���g  !      D   ,���K  !���K  ����1  ����1  !���K  !      D   ,���/  !���/  ����  ����  !���/  !      D   ,���  !���  �����  �����  !���  !      D   ,����  !����  �����  �����  !����  !      D   ,����  !����  �����  �����  !����  !      D   ,��ҿ  !��ҿ  ���ӥ  ���ӥ  !��ҿ  !      D   ,��գ  !��գ  ���։  ���։  !��գ  !      D   ,��؇  !��؇  ����m  ����m  !��؇  !      D   ,���k  !���k  ����Q  ����Q  !���k  !      D   ,���O  !���O  ����5  ����5  !���O  !      D   ,���3  !���3  ����  ����  !���3  !      D   ,���  !���  �����  �����  !���  !      D   ,����  !����  �����  �����  !����  !      D   ,����  !����  �����  �����  !����  !      D   ,����  !����  ����  ����  !����  !      D   ,���  !���  �����  �����  !���  !      D   ,���  !���  ����q  ����q  !���  !      D   ,���o  !���o  ����U  ����U  !���o  !      D   ,���S  !���S  ����9  ����9  !���S  !      D   ,���7  !���7  ����  ����  !���7  !      D   ,���  !���  ����  ����  !���  !      D   ,����  U����  ;���q  ;���q  U����  U      D   ,��ֻ  U��ֻ  ;���U  ;���U  U��ֻ  U      D   ,��ٟ  U��ٟ  ;���9  ;���9  U��ٟ  U      D   ,��܃  U��܃  ;���  ;���  U��܃  U      D   ,���g  U���g  ;���  ;���  U���g  U      D   ,���K  U���K  ;����  ;����  U���K  U      D   ,���/  U���/  ;����  ;����  U���/  U      D   ,���  U���  ;���  ;���  U���  U      D   ,����  U����  ;���  ;���  U����  U      D   ,����  U����  ;���u  ;���u  U����  U      D   ,���  U���  ;���Y  ;���Y  U���  U      D   ,���  U���  ;���=  ;���=  U���  U      D   ,����  U����  ;���!  ;���!  U����  U      D   ,���k  U���k  ;���  ;���  U���k  U      D   ,���O  U���O  ;����  ;����  U���O  U      D   ,���+  U���+  ;����  ;����  U���+  U      D   ,���  U���  ;��ϩ  ;��ϩ  U���  U      D   ,����  U����  ;��ҍ  ;��ҍ  U����  U      D   ,����  U����  ;���i  ;���i  U����  U      D   ,����  U����  ;���M  ;���M  U����  U      D   ,����  U����  ;���1  ;���1  U����  U      D   ,���{  U���{  ;���  ;���  U���{  U      D   ,���_  U���_  ;����  ;����  U���_  U      D   ,���?  U���?  ;����  ;����  U���?  U      D   ,���C  U���C  ;����  ;����  U���C  U      D   ,���'  U���'  ;����  ;����  U���'  U      D   ,���  U���  ;����  ;����  U���  U      D   ,����  U����  ;����  ;����  U����  U      D   ,����  U����  ;���m  ;���m  U����  U      D   ,����  U����  ;���Q  ;���Q  U����  U      D   ,����  U����  ;���5  ;���5  U����  U      D   ,���  U���  ;���  ;���  U���  U      D   ,���c  U���c  ;����  ;����  U���c  U      D   ,���#  U���#  ;����  ;����  U���#  U      D   ,���  U���  ;����  ;����  U���  U      D   ,����  U����  ;����  ;����  U����  U      D   ,����   �����  ����M  ����M   �����   �      D   ,����   �����  ����1  ����1   �����   �      D   ,���{   ����{  ����  ����   ����{   �      D   ,���_   ����_  �����  �����   ����_   �      D   ,���C   ����C  �����  �����   ����C   �      D   ,���'   ����'  �����  �����   ����'   �      D   ,���   ����  �����  �����   ����   �      D   ,����   �����  �����  �����   �����   �      D   ,����   �����  ����m  ����m   �����   �      D   ,����   �����  ����Q  ����Q   �����   �      D   ,����   �����  ����5  ����5   �����   �      D   ,���   ����  ����  ����   ����   �      D   ,���c   ����c  �����  �����   ����c   �      D   ,���?   ����?  �����  �����   ����?   �      D   ,���#   ����#  �����  �����   ����#   �      D   ,���   ����  �����  �����   ����   �      D   ,����   �����  �����  �����   �����   �      D   ,����   �����  ����i  ����i   �����   �      D   ,��ֻ   ���ֻ  ����U  ����U   ���ֻ   �      D   ,��ٟ   ���ٟ  ����9  ����9   ���ٟ   �      D   ,��܃   ���܃  ����  ����   ���܃   �      D   ,���g   ����g  ����  ����   ����g   �      D   ,���K   ����K  �����  �����   ����K   �      D   ,���/   ����/  �����  �����   ����/   �      D   ,���   ����  ����  ����   ����   �      D   ,����   �����  ����  ����   �����   �      D   ,����   �����  ����u  ����u   �����   �      D   ,���   ����  ����Y  ����Y   ����   �      D   ,���   ����  ����=  ����=   ����   �      D   ,����   �����  ����!  ����!   �����   �      D   ,���k   ����k  ����  ����   ����k   �      D   ,���O   ����O  �����  �����   ����O   �      D   ,���+   ����+  �����  �����   ����+   �      D   ,���   ����  ���ϩ  ���ϩ   ����   �      D   ,����   �����  ���ҍ  ���ҍ   �����   �      D   ,����   �����  ����q  ����q   �����   �      D   ,���G������G���e�������e����������G���      D   ,���'���K���'�����������������K���'���K      D   ,������K����������������������K������K      D   ,�������K�����������������������K�������K      D   ,�������K�����������������������K�������K      D   ,�������K�����������������������K�������K      D   ,�������K�����������������������K�������K      D   ,������K����������e�������e���K������K      D   ,���c���K���c�������I�������I���K���c���K      D   ,���G���K���G�������-�������-���K���G���K      D   ,���+���K���+�����������������K���+���K      D   ,������K����������������������K������K      D   ,�������K�����������������������K�������K      D   ,�������K�����������������������K�������K      D   ,�������K�����������������������K�������K      D   ,�������K�����������������������K�������K      D   ,�������K�����������i�������i���K�������K      D   ,���g���K���g�������M�������M���K���g���K      D   ,���K���K���K�������1�������1���K���K���K      D   ,���/���K���/�����������������K���/���K      D   ,������K����������������������K������K      D   ,�������K�����������������������K�������K      D   ,�������K�����������������������K�������K      D   ,��ҿ���K��ҿ������ӥ������ӥ���K��ҿ���K      D   ,��գ���K��գ������։������։���K��գ���K      D   ,��؇���K��؇�������m�������m���K��؇���K      D   ,���k���K���k�������Q�������Q���K���k���K      D   ,���O���K���O�������5�������5���K���O���K      D   ,���3���K���3�����������������K���3���K      D   ,������K����������������������K������K      D   ,�������K�����������������������K�������K      D   ,�������K�����������������������K�������K      D   ,�������K���������������������K�������K      D   ,������K����������������������K������K      D   ,������K����������q�������q���K������K      D   ,���o���K���o�������U�������U���K���o���K      D   ,���S���K���S�������9�������9���K���S���K      D   ,���7���K���7�����������������K���7���K      D   ,������K��������������������K������K      D   ,���G�������G���������������������G����      D   ,��������������e���q���e���q����������      D   ,��ֻ�����ֻ���e���U���e���U�����ֻ���      D   ,��ٟ�����ٟ���e���9���e���9�����ٟ���      D   ,��܃�����܃���e������e��������܃���      D   ,���g������g���e������e���������g���      D   ,���K������K���e�������e����������K���      D   ,���/������/���e�������e����������/���      D   ,������������e������e������������      D   ,��������������e������e�������������      D   ,��������������e���u���e���u����������      D   ,������������e���Y���e���Y���������      D   ,������������e���=���e���=���������      D   ,��������������e���!���e���!����������      D   ,���k������k���e������e���������k���      D   ,���O������O���e�������e����������O���      D   ,���+������+���e�������e����������+���      D   ,������������e��ϩ���e��ϩ���������      D   ,��������������e��ҍ���e��ҍ����������      D   ,���'������'���e�������e����������'���      D   ,������������e�������e�������������      D   ,��������������e�������e��������������      D   ,��������������e���m���e���m����������      D   ,��������������e���Q���e���Q����������      D   ,��������������e���5���e���5����������      D   ,������������e������e������������      D   ,���c������c���e�������e����������c���      D   ,������������e�������e�������������      D   ,��������������e�������e��������������      D   ,��������������e���i���e���i����������      D   ,���?������?���e�������e����������?���      D   ,��������������e���M���e���M����������      D   ,��������������e���1���e���1����������      D   ,���{������{���e������e���������{���      D   ,���_������_���e�������e����������_���      D   ,���C������C���e�������e����������C���      D   ,���#������#���e�������e����������#���      D   ,�����������������������������������      D   ,��������������������������������������      D   ,������������������i������i������������      D   ,������������������M������M������������      D   ,������������������1������1������������      D   ,���{�������{�������������������{����      D   ,���_�������_���������������������_����      D   ,���C�������C���������������������C����      D   ,���'�������'���������������������'����      D   ,�����������������������������������      D   ,��������������������������������������      D   ,������������������m������m������������      D   ,������������������Q������Q������������      D   ,������������������5������5������������      D   ,���������������������������������      D   ,���c�������c���������������������c����      D   ,���?�������?���������������������?����      D   ,���#�������#���������������������#����      D   ,���������������ϩ�����ϩ�����������      D   ,�����������������ҍ�����ҍ������������      D   ,������������������q������q������������      D   ,��ֻ������ֻ������U������U������ֻ����      D   ,��ٟ������ٟ������9������9������ٟ����      D   ,��܃������܃������������������܃����      D   ,���g�������g�������������������g����      D   ,���K�������K���������������������K����      D   ,���/�������/���������������������/����      D   ,���������������������������������      D   ,������������������������������������      D   ,������������������u������u������������      D   ,����������������Y������Y�����������      D   ,����������������=������=�����������      D   ,������������������!������!������������      D   ,���k�������k�������������������k����      D   ,���O�������O���������������������O����      D   ,���+�������+���������������������+����      D   ,  ����K  �����  �����  ����K  ����K      D   ,  ����K  �����  �����  ����K  ����K      D   ,  	����K  	�����  
�����  
����K  	����K      D   ,  ����K  �����  u����  u���K  ����K      D   ,  s���K  s����  Y����  Y���K  s���K      D   ,  W���K  W����  =����  =���K  W���K      D   ,  ;���K  ;����  !����  !���K  ;���K      D   ,  ���K  ����  ����  ���K  ���K      D   ,  ���K  ����  �����  ����K  ���K      D   ,  ����K  �����  �����  ����K  ����K      D   ,   ����K   �����  !�����  !����K   ����K      D   ,  #����K  #�����  $�����  $����K  #����K      D   ,  &����K  &�����  'y����  'y���K  &����K      D   ,  )w���K  )w����  *]����  *]���K  )w���K      D   ,  ,[���K  ,[����  -A����  -A���K  ,[���K      D   ,  /?���K  /?����  0%����  0%���K  /?���K      D   ,  2#���K  2#����  3	����  3	���K  2#���K      D   ,  5���K  5����  5�����  5����K  5���K      D   ,  7����K  7�����  8�����  8����K  7����K      D   ,  :����K  :�����  ;�����  ;����K  :����K      D   ,  =����K  =�����  >�����  >����K  =����K      D   ,  @����K  @�����  A}����  A}���K  @����K      D   ,  C{���K  C{����  Da����  Da���K  C{���K      D   ,  F_���K  F_����  GE����  GE���K  F_���K      D   ,  IC���K  IC����  J)����  J)���K  IC���K      D   ,  L'���K  L'����  M����  M���K  L'���K      D   ,  O���K  O����  O�����  O����K  O���K      D   ,  Q����K  Q�����  R�����  R����K  Q����K      D   ,  T����K  T�����  U�����  U����K  T����K      D   ,  W����K  W�����  X�����  X����K  W����K      D   ,  Z����K  Z�����  [�����  [����K  Z����K      D   ,  ]���K  ]����  ^e����  ^e���K  ]���K      D   ,  `c���K  `c����  aI����  aI���K  `c���K      D   ,  cG���K  cG����  d-����  d-���K  cG���K      D   ,  f+���K  f+����  g����  g���K  f+���K      D   ,  i���K  i����  i�����  i����K  i���K      D   ,  k����K  k�����  l�����  l����K  k����K      D   ,  6���  6���e  7����e  7����  6���      D   ,   ����K   �����  �����  ����K   ����K      D   ,  6����  6���  7����  7�����  6����      D   ,  >����  >����e  @e���e  @e���  >����      D   ,  A����  A����e  CI���e  CI���  A����      D   ,  D����  D����e  F-���e  F-���  D����      D   ,  Gw���  Gw���e  I���e  I���  Gw���      D   ,  J[���  J[���e  K����e  K����  J[���      D   ,  M?���  M?���e  N����e  N����  M?���      D   ,  P#���  P#���e  Q����e  Q����  P#���      D   ,  S���  S���e  T����e  T����  S���      D   ,  U����  U����e  W����e  W����  U����      D   ,  X����  X����e  Zi���e  Zi���  X����      D   ,  [����  [����e  ]M���e  ]M���  [����      D   ,  ^����  ^����e  `1���e  `1���  ^����      D   ,  a{���  a{���e  c���e  c���  a{���      D   ,  d_���  d_���e  e����e  e����  d_���      D   ,  gC���  gC���e  h����e  h����  gC���      D   ,  j'���  j'���e  k����e  k����  j'���      D   ,  9���  9���e  :����e  :����  9���      D   ,  ;����  ;����e  =����e  =����  ;����      D   ,  ����  ����e  %���e  %���  ����      D   ,  o���  o���e  	���e  	���  o���      D   ,  S���  S���e  ����e  ����  S���      D   ,  7���  7���e  ����e  ����  7���      D   ,  ���  ���e  ����e  ����  ���      D   ,  ����  ����e   ����e   ����  ����      D   ,  !����  !����e  #}���e  #}���  !����      D   ,  $����  $����e  &a���e  &a���  $����      D   ,  '����  '����e  )E���e  )E���  '����      D   ,  *����  *����e  ,)���e  ,)���  *����      D   ,  -s���  -s���e  /���e  /���  -s���      D   ,  0W���  0W���e  1����e  1����  0W���      D   ,  3;���  3;���e  4����e  4����  3;���      D   ,  ����  ����e  ����e  ����  ����      D   ,  ����  ����e  	y���e  	y���  ����      D   ,  ���  ���e  ����e  ����  ���      D   ,  
����  
����e  ]���e  ]���  
����      D   ,  ����  ����e  A���e  A���  ����      D   ,  �����  ����  ����  �����  �����      D   ,  �����  ����  	y���  	y����  �����      D   ,  
�����  
����  ]���  ]����  
�����      D   ,  �����  ����  A���  A����  �����      D   ,  �����  ����  %���  %����  �����      D   ,  o����  o���  	���  	����  o����      D   ,  S����  S���  ����  �����  S����      D   ,  7����  7���  ����  �����  7����      D   ,  ����  ���  ����  �����  ����      D   ,  �����  ����   ����   �����  �����      D   ,  !�����  !����  #}���  #}����  !�����      D   ,  $�����  $����  &a���  &a����  $�����      D   ,  '�����  '����  )E���  )E����  '�����      D   ,  *�����  *����  ,)���  ,)����  *�����      D   ,  -s����  -s���  /���  /����  -s����      D   ,  0W����  0W���  1����  1�����  0W����      D   ,  3;����  3;���  4����  4�����  3;����      D   ,  ����  ���  ����  �����  ����      D   ,  9����  9���  :����  :�����  9����      D   ,  ;�����  ;����  =����  =�����  ;�����      D   ,  >�����  >����  @e���  @e����  >�����      D   ,  A�����  A����  CI���  CI����  A�����      D   ,  D�����  D����  F-���  F-����  D�����      D   ,  Gw����  Gw���  I���  I����  Gw����      D   ,  J[����  J[���  K����  K�����  J[����      D   ,  M?����  M?���  N����  N�����  M?����      D   ,  P#����  P#���  Q����  Q�����  P#����      D   ,  S����  S���  T����  T�����  S����      D   ,  U�����  U����  W����  W�����  U�����      D   ,  X�����  X����  Zi���  Zi����  X�����      D   ,  [�����  [����  ]M���  ]M����  [�����      D   ,  ^�����  ^����  `1���  `1����  ^�����      D   ,  a{����  a{���  c���  c����  a{����      D   ,  d_����  d_���  e����  e�����  d_����      D   ,  gC����  gC���  h����  h�����  gC����      D   ,  j'����  j'���  k����  k�����  j'����     �     "�     " "sky130_fd_pr__nfet_01v8_8HUREQ    �   ,���}������}  �  �  �  �������}���      A   ,���&  !���&  �  �  �  �  !���&  !      A   ,���&���'���&����  �����  ����'���&���'      A  , ,���(  ����(  ?  �  ?  �  ����(  �      A  , ,���(���k���(  �����  ��������k���(���k      A  , ,  .���k  .  �  �  �  ����k  .���k      A  , ,���(�������(���k  ����k  ��������(����      ^   ,���  ���  �  U  �  U  ���        ^   ,����������  ���O  ���O�����������      ^   ,  �����  �    U    U����  �����      ^   ,������D�������  U����  U���D������D      ]  , ,���  ����  V  W  V  W  ����  �      ]  , ,������������\  W���\  W���������      B   ,���9  G���9  �����  �����  G���9  G      B   ,���  G���  �����  �����  G���  G      B   ,����  G����  ����  ����  G����  G      B   ,���#  G���#  ����m  ����m  G���#  G      B   ,���q  G���q  �����  �����  G���q  G      B   ,����  G����  ����	  ����	  G����  G      B   ,���  G���  ����W  ����W  G���  G      B   ,���[  G���[  �   �  �   �  G���[  G      B   ,  �  G  �  �  �  �  �  G  �  G      B   ,  �  G  �  �  A  �  A  G  �  G      B   ,  E  G  E  �  �  �  �  G  E  G      B   ,  �  G  �  �  	�  �  	�  G  �  G      B   ,  
�  G  
�  �  +  �  +  G  
�  G      B   ,  /  G  /  �  y  �  y  G  /  G      B   ,  }  G  }  �  �  �  �  G  }  G      B   ,���H  ����H  G���t  G���t  ����H  �      B   ,���  ����  G����  G����  ����  �      B   ,����  �����  G���  G���  �����  �      B   ,���2  ����2  G���^  G���^  ����2  �      B   ,����  �����  G����  G����  �����  �      B   ,����  �����  G����  G����  �����  �      B   ,���  ����  G���H  G���H  ����  �      B   ,���j  ����j  G   �  G   �  ����j  �      B   ,  �  �  �  G  �  G  �  �  �  �      B   ,    �    G  2  G  2  �    �      B   ,  T  �  T  G  �  G  �  �  T  �      B   ,  �  �  �  G  	�  G  	�  �  �  �      B   ,  
�  �  
�  G    G    �  
�  �      B   ,  >  �  >  G  j  G  j  �  >  �      B   ,  �  �  �  G  �  G  �  �  �  �      B   ,���9   i���9  �����  �����   i���9   i      B   ,���   i���  �����  �����   i���   i      B   ,����   i����  ����  ����   i����   i      B   ,���#   i���#  ����m  ����m   i���#   i      B   ,���q   i���q  �����  �����   i���q   i      B   ,����   i����  ����	  ����	   i����   i      B   ,���   i���  ����W  ����W   i���   i      B   ,���[   i���[  �   �  �   �   i���[   i      B   ,  �   i  �  �  �  �  �   i  �   i      B   ,  �   i  �  �  A  �  A   i  �   i      B   ,  E   i  E  �  �  �  �   i  E   i      B   ,  �   i  �  �  	�  �  	�   i  �   i      B   ,  
�   i  
�  �  +  �  +   i  
�   i      B   ,  /   i  /  �  y  �  y   i  /   i      B   ,  }   i  }  �  �  �  �   i  }   i      B   ,���9���M���9�������������������M���9���M      B   ,������M����������������������M������M      B   ,�������M���������������������M�������M      B   ,���#���M���#�������m�������m���M���#���M      B   ,���q���M���q�������������������M���q���M      B   ,�������M�����������	�������	���M�������M      B   ,������M����������W�������W���M������M      B   ,���[���M���[����   �����   ����M���[���M      B   ,  ����M  �����  �����  ����M  ����M      B   ,  ����M  �����  A����  A���M  ����M      B   ,  E���M  E����  �����  ����M  E���M      B   ,  ����M  �����  	�����  	����M  ����M      B   ,  
����M  
�����  +����  +���M  
����M      B   ,  /���M  /����  y����  y���M  /���M      B   ,  }���M  }����  �����  ����M  }���M      B   ,���H������H���M���t���M���t������H���      B   ,������������M�������M�������������      B   ,��������������M������M�������������      B   ,���2������2���M���^���M���^������2���      B   ,��������������M�������M��������������      B   ,��������������M�������M��������������      B   ,������������M���H���M���H���������      B   ,���j������j���M   ����M   �������j���      B   ,  ����  ����M  ����M  ����  ����      B   ,  ���  ���M  2���M  2���  ���      B   ,  T���  T���M  ����M  ����  T���      B   ,  ����  ����M  	����M  	����  ����      B   ,  
����  
����M  ���M  ���  
����      B   ,  >���  >���M  j���M  j���  >���      B   ,  ����  ����M  ����M  ����  ����      B   ,���9���o���9�����������������o���9���o      B   ,������o��������������������o������o      B   ,�������o�������������������o�������o      B   ,���#���o���#������m������m���o���#���o      B   ,���q���o���q�����������������o���q���o      B   ,�������o����������	������	���o�������o      B   ,������o���������W������W���o������o      B   ,���[���o���[���   ����   ����o���[���o      B   ,  ����o  ����  ����  ����o  ����o      B   ,  ����o  ����  A���  A���o  ����o      B   ,  E���o  E���  ����  ����o  E���o      B   ,  ����o  ����  	����  	����o  ����o      B   ,  
����o  
����  +���  +���o  
����o      B   ,  /���o  /���  y���  y���o  /���o      B   ,  }���o  }���  ����  ����o  }���o      B  , ,����  �����  ?   U  ?   U  �����  �      B  , ,����   �����  c   U  c   U   �����   �      B  , ,���(�������(   U����   U�����������(����      B  , ,  .����  .   U  �   U  �����  .����      B  , ,���������������G   U���G   U������������      B  , ,���������������k   U���k   U������������      B  , ,  �  �  �  ?  M  ?  M  �  �  �      B  , ,  �  �  �  ?  	�  ?  	�  �  �  �      B  , ,  
K  �  
K  ?  
�  ?  
�  �  
K  �      B  , ,  �  �  �  ?  I  ?  I  �  �  �      B  , ,  �  �  �  ?  �  ?  �  �  �  �      B  , ,  G  �  G  ?  �  ?  �  �  G  �      B  , ,  �  �  �  ?  E  ?  E  �  �  �      B  , ,  �  �  �  ?  �  ?  �  �  �  �      B  , ,  .  G  .  �  �  �  �  G  .  G      B  , ,   �  N   �  �  |  �  |  N   �  N      B  , ,     N     �  �  �  �  N     N      B  , ,  n  N  n  �    �    N  n  N      B  , ,  �  N  �  �  f  �  f  N  �  N      B  , ,  

  N  

  �  
�  �  
�  N  

  N      B  , ,  X  N  X  �    �    N  X  N      B  , ,  �  N  �  �  P  �  P  N  �  N      B  , ,  �  N  �  �  �  �  �  N  �  N      B  , ,  .  �  .  �  �  �  �  �  .  �      B  , ,   �  
�   �  �  |  �  |  
�   �  
�      B  , ,     
�     �  �  �  �  
�     
�      B  , ,  n  
�  n  �    �    
�  n  
�      B  , ,  �  
�  �  �  f  �  f  
�  �  
�      B  , ,  

  
�  

  �  
�  �  
�  
�  

  
�      B  , ,  X  
�  X  �    �    
�  X  
�      B  , ,  �  
�  �  �  P  �  P  
�  �  
�      B  , ,  �  
�  �  �  �  �  �  
�  �  
�      B  , ,  .  �  .  I  �  I  �  �  .  �      B  , ,   �  	�   �  
P  |  
P  |  	�   �  	�      B  , ,     	�     
P  �  
P  �  	�     	�      B  , ,  n  	�  n  
P    
P    	�  n  	�      B  , ,  �  	�  �  
P  f  
P  f  	�  �  	�      B  , ,  

  	�  

  
P  
�  
P  
�  	�  

  	�      B  , ,  X  	�  X  
P    
P    	�  X  	�      B  , ,  �  	�  �  
P  P  
P  P  	�  �  	�      B  , ,  �  	�  �  
P  �  
P  �  	�  �  	�      B  , ,  .  
K  .  
�  �  
�  �  
K  .  
K      B  , ,   �  R   �  �  |  �  |  R   �  R      B  , ,     R     �  �  �  �  R     R      B  , ,  n  R  n  �    �    R  n  R      B  , ,  �  R  �  �  f  �  f  R  �  R      B  , ,  

  R  

  �  
�  �  
�  R  

  R      B  , ,  X  R  X  �    �    R  X  R      B  , ,  �  R  �  �  P  �  P  R  �  R      B  , ,  �  R  �  �  �  �  �  R  �  R      B  , ,  .  �  .  	�  �  	�  �  �  .  �      B  , ,   �  �   �  �  |  �  |  �   �  �      B  , ,     �     �  �  �  �  �     �      B  , ,  n  �  n  �    �    �  n  �      B  , ,  �  �  �  �  f  �  f  �  �  �      B  , ,  

  �  

  �  
�  �  
�  �  

  �      B  , ,  X  �  X  �    �    �  X  �      B  , ,  �  �  �  �  P  �  P  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  .  �  .  M  �  M  �  �  .  �      B  , ,   �  �   �  T  |  T  |  �   �  �      B  , ,     �     T  �  T  �  �     �      B  , ,  n  �  n  T    T    �  n  �      B  , ,  �  �  �  T  f  T  f  �  �  �      B  , ,  

  �  

  T  
�  T  
�  �  

  �      B  , ,  X  �  X  T    T    �  X  �      B  , ,  �  �  �  T  P  T  P  �  �  �      B  , ,  �  �  �  T  �  T  �  �  �  �      B  , ,  .  O  .  �  �  �  �  O  .  O      B  , ,   �  V   �     |     |  V   �  V      B  , ,     V        �     �  V     V      B  , ,  n  V  n            V  n  V      B  , ,  �  V  �     f     f  V  �  V      B  , ,  

  V  

     
�     
�  V  

  V      B  , ,  X  V  X            V  X  V      B  , ,  �  V  �     P     P  V  �  V      B  , ,  �  V  �     �     �  V  �  V      B  , ,  .  �  .  �  �  �  �  �  .  �      B  , ,   �     �  �  |  �  |     �        B  , ,          �  �  �  �             B  , ,  n    n  �    �      n        B  , ,  �    �  �  f  �  f    �        B  , ,  

    

  �  
�  �  
�    

        B  , ,  X    X  �    �      X        B  , ,  �    �  �  P  �  P    �        B  , ,  �    �  �  �  �  �    �        B  , ,  .  �  .  Q  �  Q  �  �  .  �      B  , ,  .  S  .  �  �  �  �  S  .  S      B  , ,   �  �   �  ?  �  ?  �  �   �  �      B  , ,  �   �  �  c  �  c  �   �  �   �      B  , ,  G   �  G  c  �  c  �   �  G   �      B  , ,  �   �  �  c  ?  c  ?   �  �   �      B  , ,  �   �  �  c  	�  c  	�   �  �   �      B  , ,  1   �  1  c  �  c  �   �  1   �      B  , ,     �    c  )  c  )   �     �      B  , ,  �   �  �  c  w  c  w   �  �   �      B  , ,  .   �  .  �  �  �  �   �  .   �      B  , ,  S  �  S  ?  �  ?  �  �  S  �      B  , ,  �  �  �  ?  Q  ?  Q  �  �  �      B  , ,  �  �  �  ?  �  ?  �  �  �  �      B  , ,  O  �  O  ?  �  ?  �  �  O  �      B  , ,���(  ����(  M����  M����  ����(  �      B  , ,���b  ����b  ����  ����  ����b  �      B  , ,���  ����  ����Z  ����Z  ����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,���L  ����L  �����  �����  ����L  �      B  , ,����  �����  ����D  ����D  �����  �      B  , ,����  �����  �����  �����  �����  �      B  , ,���6  ����6  �����  �����  ����6  �      B  , ,����  �����  ����.  ����.  �����  �      B  , ,���L  
����L  �����  �����  
����L  
�      B  , ,����  
�����  ����D  ����D  
�����  
�      B  , ,����  
�����  �����  �����  
�����  
�      B  , ,���6  
����6  �����  �����  
����6  
�      B  , ,����  
�����  ����.  ����.  
�����  
�      B  , ,���  ����  ?����  ?����  ����  �      B  , ,���W  ����W  ?���  ?���  ����W  �      B  , ,���g  ����g  ?���  ?���  ����g  �      B  , ,���(  G���(  �����  �����  G���(  G      B  , ,���(  O���(  �����  �����  O���(  O      B  , ,���b  ����b  T���  T���  ����b  �      B  , ,���  ����  T���Z  T���Z  ����  �      B  , ,����  �����  T���  T���  �����  �      B  , ,���L  ����L  T����  T����  ����L  �      B  , ,����  �����  T���D  T���D  �����  �      B  , ,����  �����  T����  T����  �����  �      B  , ,���6  ����6  T����  T����  ����6  �      B  , ,����  �����  T���.  T���.  �����  �      B  , ,���  ����  ?���e  ?���e  ����  �      B  , ,���(  ����(  �����  �����  ����(  �      B  , ,���b  N���b  ����  ����  N���b  N      B  , ,���  N���  ����Z  ����Z  N���  N      B  , ,����  N����  ����  ����  N����  N      B  , ,���(  
K���(  
�����  
�����  
K���(  
K      B  , ,���b  	����b  
P���  
P���  	����b  	�      B  , ,���  	����  
P���Z  
P���Z  	����  	�      B  , ,����  	�����  
P���  
P���  	�����  	�      B  , ,���(  ����(  �����  �����  ����(  �      B  , ,���b  V���b   ���   ���  V���b  V      B  , ,���  V���   ���Z   ���Z  V���  V      B  , ,����  V����   ���   ���  V����  V      B  , ,���L  V���L   ����   ����  V���L  V      B  , ,����  V����   ���D   ���D  V����  V      B  , ,����  V����   ����   ����  V����  V      B  , ,���6  V���6   ����   ����  V���6  V      B  , ,����  V����   ���.   ���.  V����  V      B  , ,���L  	����L  
P����  
P����  	����L  	�      B  , ,����  	�����  
P���D  
P���D  	�����  	�      B  , ,����  	�����  
P����  
P����  	�����  	�      B  , ,���6  	����6  
P����  
P����  	����6  	�      B  , ,����  	�����  
P���.  
P���.  	�����  	�      B  , ,���L  N���L  �����  �����  N���L  N      B  , ,����  N����  ����D  ����D  N����  N      B  , ,����  N����  �����  �����  N����  N      B  , ,���6  N���6  �����  �����  N���6  N      B  , ,���(  ����(  Q����  Q����  ����(  �      B  , ,���b  ���b  ����  ����  ���b        B  , ,���  ���  ����Z  ����Z  ���        B  , ,����  ����  ����  ����  ����        B  , ,���L  ���L  �����  �����  ���L        B  , ,����  ����  ����D  ����D  ����        B  , ,����  ����  �����  �����  ����        B  , ,���6  ���6  �����  �����  ���6        B  , ,����  ����  ����.  ����.  ����        B  , ,����  N����  ����.  ����.  N����  N      B  , ,���  ����  ?���  ?���  ����  �      B  , ,���c  ����c  ?���  ?���  ����c  �      B  , ,���  ����  ?���a  ?���a  ����  �      B  , ,���  ����  ?����  ?����  ����  �      B  , ,���(  ����(  	�����  	�����  ����(  �      B  , ,���b  R���b  ����  ����  R���b  R      B  , ,���  R���  ����Z  ����Z  R���  R      B  , ,����  R����  ����  ����  R����  R      B  , ,���(  S���(  �����  �����  S���(  S      B  , ,���L  R���L  �����  �����  R���L  R      B  , ,���(   ����(  �����  �����   ����(   �      B  , ,���   ����  c���3  c���3   ����   �      B  , ,����   �����  c���  c���   �����   �      B  , ,���%   ����%  c����  c����   ����%   �      B  , ,���s   ����s  c���  c���   ����s   �      B  , ,����   �����  c���k  c���k   �����   �      B  , ,���   ����  c����  c����   ����   �      B  , ,���]   ����]  c���  c���   ����]   �      B  , ,����  R����  ����D  ����D  R����  R      B  , ,����  R����  �����  �����  R����  R      B  , ,���6  R���6  �����  �����  R���6  R      B  , ,����  R����  ����.  ����.  R����  R      B  , ,���_  ����_  ?���	  ?���	  ����_  �      B  , ,����  �����  ?���]  ?���]  �����  �      B  , ,���  ����  ?����  ?����  ����  �      B  , ,���[  ����[  ?���  ?���  ����[  �      B  , ,����  �����  ?���Y  ?���Y  �����  �      B  , ,���(  ����(  I����  I����  ����(  �      B  , ,���b  
����b  ����  ����  
����b  
�      B  , ,���  
����  ����Z  ����Z  
����  
�      B  , ,����  
�����  ����  ����  
�����  
�      B  , ,���������������G������G���������������      B  , ,���%�������%���G�������G�����������%����      B  , ,���s�������s���G������G����������s����      B  , ,���������������G���k���G���k������������      B  , ,�������������G�������G���������������      B  , ,���]�������]���G������G����������]����      B  , ,���(���W���(�����������������W���(���W      B  , ,���(������(����������������������(���      B  , ,���(�������(���Y�������Y�����������(����      B  , ,���b���T���b�����������������T���b���T      B  , ,������T����������Z�������Z���T������T      B  , ,�������T���������������������T�������T      B  , ,���L���T���L�������������������T���L���T      B  , ,�������T�����������D�������D���T�������T      B  , ,�������T�����������������������T�������T      B  , ,���6���T���6�������������������T���6���T      B  , ,�������T�����������.�������.���T�������T      B  , ,���(���[���(�����������������[���(���[      B  , ,���b��� ���b����������������� ���b���       B  , ,������ ����������Z�������Z��� ������       B  , ,������� ��������������������� �������       B  , ,���L��� ���L������������������� ���L���       B  , ,������� �����������D�������D��� �������       B  , ,������� ����������������������� �������       B  , ,���6��� ���6������������������� ���6���       B  , ,������� �����������.�������.��� �������       B  , ,���(������(����������������������(���      B  , ,���b�������b���V������V����������b����      B  , ,�������������V���Z���V���Z�����������      B  , ,���������������V������V���������������      B  , ,���L�������L���V�������V�����������L����      B  , ,���������������V���D���V���D������������      B  , ,���������������V�������V����������������      B  , ,���6�������6���V�������V�����������6����      B  , ,���������������V���.���V���.������������      B  , ,���(�������(���]�������]�����������(����      B  , ,���b���X���b���������������X���b���X      B  , ,������X���������Z������Z���X������X      B  , ,�������X�������������������X�������X      B  , ,���L���X���L�����������������X���L���X      B  , ,�������X����������D������D���X�������X      B  , ,�������X���������������������X�������X      B  , ,���6���X���6�����������������X���6���X      B  , ,�������X����������.������.���X�������X      B  , ,���(���_���(���	�������	�������_���(���_      B  , ,���b������b��������������������b���      B  , ,����������������Z�������Z���������      B  , ,�����������������������������������      B  , ,���L������L����������������������L���      B  , ,������������������D�������D����������      B  , ,�������������������������������������      B  , ,���6������6����������������������6���      B  , ,������������������.�������.����������      B  , ,���(������(����������������������(���      B  , ,���b�������b���Z������Z����������b����      B  , ,�������������Z���Z���Z���Z�����������      B  , ,���������������Z������Z���������������      B  , ,���L�������L���Z�������Z�����������L����      B  , ,���������������Z���D���Z���D������������      B  , ,���������������Z�������Z����������������      B  , ,���6�������6���Z�������Z�����������6����      B  , ,���������������Z���.���Z���.������������      B  , ,���(������(���a�������a����������(���      B  , ,���b���\���b���������������\���b���\      B  , ,������\���������Z������Z���\������\      B  , ,�������\�������������������\�������\      B  , ,���L���\���L�����������������\���L���\      B  , ,�������\����������D������D���\�������\      B  , ,�������\���������������������\�������\      B  , ,���6���\���6�����������������\���6���\      B  , ,�������\����������.������.���\�������\      B  , ,���(���c���(�����������������c���(���c      B  , ,���b������b������������������b���      B  , ,���������������Z������Z���������      B  , ,���������������������������������      B  , ,���L������L��������������������L���      B  , ,�����������������D������D����������      B  , ,�����������������������������������      B  , ,���6������6��������������������6���      B  , ,�����������������.������.����������      B  , ,���(������(��������������������(���      B  , ,���g�������g���k������k����������g����      B  , ,�������������k���e���k���e�����������      B  , ,�������������k������k��������������      B  , ,���c�������c���k������k����������c����      B  , ,�������������k���a���k���a�����������      B  , ,�������������k�������k���������������      B  , ,���_�������_���k���	���k���	�������_����      B  , ,���������������k���]���k���]������������      B  , ,�������������k�������k���������������      B  , ,���[�������[���k������k����������[����      B  , ,���������������k���Y���k���Y������������      B  , ,�������������k�������k���������������      B  , ,���W�������W���k������k����������W����      B  , ,�������������G���3���G���3�����������      B  , ,  ����   �����  P����  P���   ����       B  , ,  ����   �����  �����  ����   ����       B  , ,  .���[  .���  ����  ����[  .���[      B  , ,   ����   �����  |����  |���   ����      B  , ,   ���   ����  �����  ����   ���      B  , ,  n���  n����  ����  ���  n���      B  , ,  ����  �����  f����  f���  ����      B  , ,  

���  

����  
�����  
����  

���      B  , ,  X���  X����  ����  ���  X���      B  , ,  ����  �����  P����  P���  ����      B  , ,  ����  �����  �����  ����  ����      B  , ,  .���_  .���	  ����	  ����_  .���_      B  , ,   ����T   �����  |����  |���T   ����T      B  , ,   ���T   ����  �����  ����T   ���T      B  , ,  n���T  n����  ����  ���T  n���T      B  , ,  ����T  �����  f����  f���T  ����T      B  , ,  

���T  

����  
�����  
����T  

���T      B  , ,  X���T  X����  ����  ���T  X���T      B  , ,  ����T  �����  P����  P���T  ����T      B  , ,  ����T  �����  �����  ����T  ����T      B  , ,  .����  .���Y  ����Y  �����  .����      B  , ,   �����   ����Z  |���Z  |����   �����      B  , ,   ����   ���Z  ����Z  �����   ����      B  , ,  n����  n���Z  ���Z  ����  n����      B  , ,  �����  ����Z  f���Z  f����  �����      B  , ,  

����  

���Z  
����Z  
�����  

����      B  , ,  X����  X���Z  ���Z  ����  X����      B  , ,  �����  ����Z  P���Z  P����  �����      B  , ,  �����  ����Z  ����Z  �����  �����      B  , ,  .���  .����  �����  ����  .���      B  , ,   �����   ����V  |���V  |����   �����      B  , ,   ����   ���V  ����V  �����   ����      B  , ,  n����  n���V  ���V  ����  n����      B  , ,  �����  ����V  f���V  f����  �����      B  , ,  

����  

���V  
����V  
�����  

����      B  , ,  X����  X���V  ���V  ����  X����      B  , ,  �����  ����V  P���V  P����  �����      B  , ,  �����  ����V  ����V  �����  �����      B  , ,  .���  .����  �����  ����  .���      B  , ,   ����\   ����  |���  |���\   ����\      B  , ,   ���\   ���  ����  ����\   ���\      B  , ,  n���\  n���  ���  ���\  n���\      B  , ,  ����\  ����  f���  f���\  ����\      B  , ,  

���\  

���  
����  
����\  

���\      B  , ,  X���\  X���  ���  ���\  X���\      B  , ,  ����\  ����  P���  P���\  ����\      B  , ,  ����\  ����  ����  ����\  ����\      B  , ,  .���  .���a  ����a  ����  .���      B  , ,  G����  G���G  ����G  �����  G����      B  , ,  �����  ����G  ?���G  ?����  �����      B  , ,  �����  ����G  	����G  	�����  �����      B  , ,  1����  1���G  ����G  �����  1����      B  , ,  ����  ���G  )���G  )����  ����      B  , ,  �����  ����G  w���G  w����  �����      B  , ,  .���W  .���  ����  ����W  .���W      B  , ,  �����  ����G  ����G  �����  �����      B  , ,  .���  .����  �����  ����  .���      B  , ,   ����   ����  |���  |���   ����      B  , ,   ���   ���  ����  ����   ���      B  , ,  n���  n���  ���  ���  n���      B  , ,  ����  ����  f���  f���  ����      B  , ,  

���  

���  
����  
����  

���      B  , ,  X���  X���  ���  ���  X���      B  , ,  ����  ����  P���  P���  ����      B  , ,  ����  ����  ����  ����  ����      B  , ,  .���c  .���  ����  ����c  .���c      B  , ,   ����X   ����  |���  |���X   ����X      B  , ,  .���  .���  ����  ����  .���      B  , ,   ���X   ���  ����  ����X   ���X      B  , ,  n���X  n���  ���  ���X  n���X      B  , ,  ����X  ����  f���  f���X  ����X      B  , ,  

���X  

���  
����  
����X  

���X      B  , ,  X���X  X���  ���  ���X  X���X      B  , ,  ����X  ����  P���  P���X  ����X      B  , ,  ����X  ����  ����  ����X  ����X      B  , ,  .����  .���]  ����]  �����  .����      B  , ,   ����    �����  |����  |���    ����       B  , ,   ���    ����  �����  ����    ���       B  , ,  n���   n����  ����  ���   n���       B  , ,  ����   �����  f����  f���   ����       B  , ,  

���   

����  
�����  
����   

���       B  , ,  X���   X����  ����  ���   X���       B  , ,   �����   ����k  ����k  �����   �����      B  , ,  S����  S���k  ����k  �����  S����      B  , ,  �����  ����k  Q���k  Q����  �����      B  , ,  �����  ����k  ����k  �����  �����      B  , ,  O����  O���k  ����k  �����  O����      B  , ,  �����  ����k  M���k  M����  �����      B  , ,  �����  ����k  	����k  	�����  �����      B  , ,  
K����  
K���k  
����k  
�����  
K����      B  , ,  �����  ����k  I���k  I����  �����      B  , ,  �����  ����k  ����k  �����  �����      B  , ,  G����  G���k  ����k  �����  G����      B  , ,  �����  ����k  E���k  E����  �����      B  , ,  �����  ����k  ����k  �����  �����      _   ,���%���9���%  �  �  �  ����9���%���9      C   ,���(  ����(  ?  �  ?  �  ����(  �      C   ,���(���k���(  �����  ��������k���(���k      C   ,���b  ���b  ����  ����  ���b        C   ,���  ���  ����Z  ����Z  ���        C   ,����  ����  ����  ����  ����        C   ,���L  ���L  �����  �����  ���L        C   ,����  ����  ����D  ����D  ����        C   ,����  ����  �����  �����  ����        C   ,���6  ���6  �����  �����  ���6        C   ,����  ����  ����.  ����.  ����        C   ,   �     �  �  |  �  |     �        C   ,          �  �  �  �             C   ,  n    n  �    �      n        C   ,  �    �  �  f  �  f    �        C   ,  

    

  �  
�  �  
�    

        C   ,  X    X  �    �      X        C   ,  �    �  �  P  �  P    �        C   ,  �    �  �  �  �  �    �        C   ,���9   ����9  c����  c����   ����9   �      C   ,���   ����  c����  c����   ����   �      C   ,����   �����  c���  c���   �����   �      C   ,���#   ����#  c���m  c���m   ����#   �      C   ,���q   ����q  c����  c����   ����q   �      C   ,����   �����  c���	  c���	   �����   �      C   ,���   ����  c���W  c���W   ����   �      C   ,���[   ����[  c   �  c   �   ����[   �      C   ,  �   �  �  c  �  c  �   �  �   �      C   ,  �   �  �  c  A  c  A   �  �   �      C   ,  E   �  E  c  �  c  �   �  E   �      C   ,  �   �  �  c  	�  c  	�   �  �   �      C   ,  
�   �  
�  c  +  c  +   �  
�   �      C   ,  /   �  /  c  y  c  y   �  /   �      C   ,  }   �  }  c  �  c  �   �  }   �      C   ,���9�������9���G�������G�����������9����      C   ,�������������G�������G���������������      C   ,���������������G������G���������������      C   ,���#�������#���G���m���G���m�������#����      C   ,���q�������q���G�������G�����������q����      C   ,���������������G���	���G���	������������      C   ,�������������G���W���G���W�����������      C   ,���[�������[���G   ����G   ��������[����      C   ,  �����  ����G  ����G  �����  �����      C   ,  �����  ����G  A���G  A����  �����      C   ,  E����  E���G  ����G  �����  E����      C   ,  �����  ����G  	����G  	�����  �����      C   ,  
�����  
����G  +���G  +����  
�����      C   ,  /����  /���G  y���G  y����  /����      C   ,  }����  }���G  ����G  �����  }����      C   ,���b������b��������������������b���      C   ,����������������Z�������Z���������      C   ,�����������������������������������      C   ,���L������L����������������������L���      C   ,������������������D�������D����������      C   ,�������������������������������������      C   ,���6������6����������������������6���      C   ,������������������.�������.����������      C   ,   ����   �����  |����  |���   ����      C   ,   ���   ����  �����  ����   ���      C   ,  n���  n����  ����  ���  n���      C   ,  ����  �����  f����  f���  ����      C   ,  

���  

����  
�����  
����  

���      C   ,  X���  X����  ����  ���  X���      C   ,  ����  �����  P����  P���  ����      C   ,  ����  �����  �����  ����  ����      C   ,  .���k  .  �  �  �  ����k  .���k      C   ,���(�������(���k  ����k  ��������(����      C  , ,����   �����  c   U  c   U   �����   �      C  , ,���������������G   U���G   U������������      C  , ,  n  �  n  >    >    �  n  �      C  , ,  �  �  �  >  f  >  f  �  �  �      C  , ,  

  �  

  >  
�  >  
�  �  

  �      C  , ,  X  �  X  >    >    �  X  �      C  , ,  �  �  �  >  P  >  P  �  �  �      C  , ,  �  �  �  >  �  >  �  �  �  �      C  , ,   �  ,   �  �  |  �  |  ,   �  ,      C  , ,     ,     �  �  �  �  ,     ,      C  , ,  n  ,  n  �    �    ,  n  ,      C  , ,  �  ,  �  �  f  �  f  ,  �  ,      C  , ,  

  ,  

  �  
�  �  
�  ,  

  ,      C  , ,  X  ,  X  �    �    ,  X  ,      C  , ,  �  ,  �  �  P  �  P  ,  �  ,      C  , ,  �  ,  �  �  �  �  �  ,  �  ,      C  , ,   �  	�   �  
n  |  
n  |  	�   �  	�      C  , ,     	�     
n  �  
n  �  	�     	�      C  , ,  n  	�  n  
n    
n    	�  n  	�      C  , ,  �  	�  �  
n  f  
n  f  	�  �  	�      C  , ,  

  	�  

  
n  
�  
n  
�  	�  

  	�      C  , ,  X  	�  X  
n    
n    	�  X  	�      C  , ,  �  	�  �  
n  P  
n  P  	�  �  	�      C  , ,  �  	�  �  
n  �  
n  �  	�  �  	�      C  , ,   �  \   �  	  |  	  |  \   �  \      C  , ,     \     	  �  	  �  \     \      C  , ,  n  \  n  	    	    \  n  \      C  , ,  �  \  �  	  f  	  f  \  �  \      C  , ,  

  \  

  	  
�  	  
�  \  

  \      C  , ,  X  \  X  	    	    \  X  \      C  , ,  �  \  �  	  P  	  P  \  �  \      C  , ,  �  \  �  	  �  	  �  \  �  \      C  , ,   �  �   �  �  |  �  |  �   �  �      C  , ,     �     �  �  �  �  �     �      C  , ,  n  �  n  �    �    �  n  �      C  , ,  �  �  �  �  f  �  f  �  �  �      C  , ,  

  �  

  �  
�  �  
�  �  

  �      C  , ,  X  �  X  �    �    �  X  �      C  , ,  �  �  �  �  P  �  P  �  �  �      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,   �  �   �  6  |  6  |  �   �  �      C  , ,     �     6  �  6  �  �     �      C  , ,  n  �  n  6    6    �  n  �      C  , ,  �  �  �  6  f  6  f  �  �  �      C  , ,  

  �  

  6  
�  6  
�  �  

  �      C  , ,  X  �  X  6    6    �  X  �      C  , ,  �  �  �  6  P  6  P  �  �  �      C  , ,  �  �  �  6  �  6  �  �  �  �      C  , ,   �  $   �  �  |  �  |  $   �  $      C  , ,     $     �  �  �  �  $     $      C  , ,  n  $  n  �    �    $  n  $      C  , ,  �  $  �  �  f  �  f  $  �  $      C  , ,  

  $  

  �  
�  �  
�  $  

  $      C  , ,  X  $  X  �    �    $  X  $      C  , ,  �  $  �  �  P  �  P  $  �  $      C  , ,  �  $  �  �  �  �  �  $  �  $      C  , ,   �  �   �  f  |  f  |  �   �  �      C  , ,     �     f  �  f  �  �     �      C  , ,  n  �  n  f    f    �  n  �      C  , ,  �  �  �  f  f  f  f  �  �  �      C  , ,  

  �  

  f  
�  f  
�  �  

  �      C  , ,  X  �  X  f    f    �  X  �      C  , ,  �  �  �  f  P  f  P  �  �  �      C  , ,  �  �  �  f  �  f  �  �  �  �      C  , ,   �  �   �  >  |  >  |  �   �  �      C  , ,  �   �  �  c  �  c  �   �  �   �      C  , ,  G   �  G  c  �  c  �   �  G   �      C  , ,  �   �  �  c  ?  c  ?   �  �   �      C  , ,  �   �  �  c  	�  c  	�   �  �   �      C  , ,  1   �  1  c  �  c  �   �  1   �      C  , ,     �    c  )  c  )   �     �      C  , ,  �   �  �  c  w  c  w   �  �   �      C  , ,     �     >  �  >  �  �     �      C  , ,���  	����  
n���Z  
n���Z  	����  	�      C  , ,����  	�����  
n���  
n���  	�����  	�      C  , ,���L  	����L  
n����  
n����  	����L  	�      C  , ,����  	�����  
n���D  
n���D  	�����  	�      C  , ,����  	�����  
n����  
n����  	�����  	�      C  , ,���6  	����6  
n����  
n����  	����6  	�      C  , ,����  	�����  
n���.  
n���.  	�����  	�      C  , ,���b  ����b  6���  6���  ����b  �      C  , ,���  ����  6���Z  6���Z  ����  �      C  , ,����  �����  6���  6���  �����  �      C  , ,���L  ����L  6����  6����  ����L  �      C  , ,����  �����  6���D  6���D  �����  �      C  , ,����  �����  6����  6����  �����  �      C  , ,���6  ����6  6����  6����  ����6  �      C  , ,����  �����  6���.  6���.  �����  �      C  , ,���b  ,���b  ����  ����  ,���b  ,      C  , ,���  ,���  ����Z  ����Z  ,���  ,      C  , ,����  ,����  ����  ����  ,����  ,      C  , ,���L  ,���L  �����  �����  ,���L  ,      C  , ,����  ,����  ����D  ����D  ,����  ,      C  , ,����  ,����  �����  �����  ,����  ,      C  , ,���6  ,���6  �����  �����  ,���6  ,      C  , ,����  ,����  ����.  ����.  ,����  ,      C  , ,���b  $���b  ����  ����  $���b  $      C  , ,���  $���  ����Z  ����Z  $���  $      C  , ,����  $����  ����  ����  $����  $      C  , ,���L  $���L  �����  �����  $���L  $      C  , ,����  $����  ����D  ����D  $����  $      C  , ,����  $����  �����  �����  $����  $      C  , ,���6  $���6  �����  �����  $���6  $      C  , ,����  $����  ����.  ����.  $����  $      C  , ,���b  \���b  	���  	���  \���b  \      C  , ,���  \���  	���Z  	���Z  \���  \      C  , ,����  \����  	���  	���  \����  \      C  , ,���L  \���L  	����  	����  \���L  \      C  , ,����  \����  	���D  	���D  \����  \      C  , ,����  \����  	����  	����  \����  \      C  , ,���6  \���6  	����  	����  \���6  \      C  , ,����  \����  	���.  	���.  \����  \      C  , ,���b  ����b  f���  f���  ����b  �      C  , ,���  ����  f���Z  f���Z  ����  �      C  , ,����  �����  f���  f���  �����  �      C  , ,���L  ����L  f����  f����  ����L  �      C  , ,����  �����  f���D  f���D  �����  �      C  , ,����  �����  f����  f����  �����  �      C  , ,���6  ����6  f����  f����  ����6  �      C  , ,����  �����  f���.  f���.  �����  �      C  , ,���b  ����b  >���  >���  ����b  �      C  , ,���  ����  >���Z  >���Z  ����  �      C  , ,����  �����  >���  >���  �����  �      C  , ,���L  ����L  >����  >����  ����L  �      C  , ,����  �����  >���D  >���D  �����  �      C  , ,����  �����  >����  >����  �����  �      C  , ,���6  ����6  >����  >����  ����6  �      C  , ,����  �����  >���.  >���.  �����  �      C  , ,���   ����  c���3  c���3   ����   �      C  , ,����   �����  c���  c���   �����   �      C  , ,���%   ����%  c����  c����   ����%   �      C  , ,���s   ����s  c���  c���   ����s   �      C  , ,����   �����  c���k  c���k   �����   �      C  , ,���   ����  c����  c����   ����   �      C  , ,���]   ����]  c���  c���   ����]   �      C  , ,���b  ����b  ����  ����  ����b  �      C  , ,���  ����  ����Z  ����Z  ����  �      C  , ,����  �����  ����  ����  �����  �      C  , ,���L  ����L  �����  �����  ����L  �      C  , ,����  �����  ����D  ����D  �����  �      C  , ,����  �����  �����  �����  �����  �      C  , ,���6  ����6  �����  �����  ����6  �      C  , ,����  �����  ����.  ����.  �����  �      C  , ,���b  	����b  
n���  
n���  	����b  	�      C  , ,���������������G������G���������������      C  , ,���%�������%���G�������G�����������%����      C  , ,���s�������s���G������G����������s����      C  , ,���������������G���k���G���k������������      C  , ,�������������G�������G���������������      C  , ,���]�������]���G������G����������]����      C  , ,�������������G���3���G���3�����������      C  , ,���b�������b���D������D����������b����      C  , ,�������������D���Z���D���Z�����������      C  , ,���������������D������D���������������      C  , ,���L�������L���D�������D�����������L����      C  , ,���������������D���D���D���D������������      C  , ,���������������D�������D����������������      C  , ,���6�������6���D�������D�����������6����      C  , ,���������������D���.���D���.������������      C  , ,���b���2���b�����������������2���b���2      C  , ,������2����������Z�������Z���2������2      C  , ,�������2���������������������2�������2      C  , ,���L���2���L�������������������2���L���2      C  , ,�������2�����������D�������D���2�������2      C  , ,�������2�����������������������2�������2      C  , ,���6���2���6�������������������2���6���2      C  , ,�������2�����������.�������.���2�������2      C  , ,���b�������b���t������t����������b����      C  , ,�������������t���Z���t���Z�����������      C  , ,���������������t������t���������������      C  , ,���L�������L���t�������t�����������L����      C  , ,���������������t���D���t���D������������      C  , ,���������������t�������t����������������      C  , ,���6�������6���t�������t�����������6����      C  , ,���������������t���.���t���.������������      C  , ,���b���b���b���������������b���b���b      C  , ,������b���������Z������Z���b������b      C  , ,�������b�������������������b�������b      C  , ,���L���b���L�����������������b���L���b      C  , ,�������b����������D������D���b�������b      C  , ,�������b���������������������b�������b      C  , ,���6���b���6�����������������b���6���b      C  , ,�������b����������.������.���b�������b      C  , ,���b�������b���������������������b����      C  , ,�����������������Z�������Z�����������      C  , ,��������������������������������������      C  , ,���L�������L�����������������������L����      C  , ,�������������������D�������D������������      C  , ,����������������������������������������      C  , ,���6�������6�����������������������6����      C  , ,�������������������.�������.������������      C  , ,���b�������b���<������<����������b����      C  , ,�������������<���Z���<���Z�����������      C  , ,���������������<������<���������������      C  , ,���L�������L���<�������<�����������L����      C  , ,���������������<���D���<���D������������      C  , ,���������������<�������<����������������      C  , ,���6�������6���<�������<�����������6����      C  , ,���������������<���.���<���.������������      C  , ,���b���*���b�����������������*���b���*      C  , ,������*����������Z�������Z���*������*      C  , ,�������*���������������������*�������*      C  , ,���L���*���L�������������������*���L���*      C  , ,�������*�����������D�������D���*�������*      C  , ,�������*�����������������������*�������*      C  , ,���6���*���6�������������������*���6���*      C  , ,�������*�����������.�������.���*�������*      C  , ,���b�������b���l������l����������b����      C  , ,�������������l���Z���l���Z�����������      C  , ,���������������l������l���������������      C  , ,���L�������L���l�������l�����������L����      C  , ,���������������l���D���l���D������������      C  , ,���������������l�������l����������������      C  , ,���6�������6���l�������l�����������6����      C  , ,���������������l���.���l���.������������      C  , ,   ���b   ���  ����  ����b   ���b      C  , ,  n���b  n���  ���  ���b  n���b      C  , ,  ����b  ����  f���  f���b  ����b      C  , ,  

���b  

���  
����  
����b  

���b      C  , ,  X���b  X���  ���  ���b  X���b      C  , ,  ����b  ����  P���  P���b  ����b      C  , ,  ����b  ����  ����  ����b  ����b      C  , ,   ���2   ����  �����  ����2   ���2      C  , ,  n���2  n����  ����  ���2  n���2      C  , ,  ����2  �����  f����  f���2  ����2      C  , ,  

���2  

����  
�����  
����2  

���2      C  , ,  X���2  X����  ����  ���2  X���2      C  , ,  ����2  �����  P����  P���2  ����2      C  , ,  ����2  �����  �����  ����2  ����2      C  , ,   ����   ���D  ����D  �����   ����      C  , ,   �����   �����  |����  |����   �����      C  , ,   ����   ����  �����  �����   ����      C  , ,  n����  n����  ����  ����  n����      C  , ,  �����  �����  f����  f����  �����      C  , ,  

����  

����  
�����  
�����  

����      C  , ,  X����  X����  ����  ����  X����      C  , ,  �����  �����  P����  P����  �����      C  , ,  �����  �����  �����  �����  �����      C  , ,  n����  n���D  ���D  ����  n����      C  , ,  �����  ����D  f���D  f����  �����      C  , ,  

����  

���D  
����D  
�����  

����      C  , ,  X����  X���D  ���D  ����  X����      C  , ,  �����  ����D  P���D  P����  �����      C  , ,  �����  ����D  ����D  �����  �����      C  , ,  G����  G���G  ����G  �����  G����      C  , ,   �����   ����t  |���t  |����   �����      C  , ,   �����   ����<  |���<  |����   �����      C  , ,   ����   ���<  ����<  �����   ����      C  , ,  n����  n���<  ���<  ����  n����      C  , ,  �����  ����<  f���<  f����  �����      C  , ,  

����  

���<  
����<  
�����  

����      C  , ,  X����  X���<  ���<  ����  X����      C  , ,  �����  ����<  P���<  P����  �����      C  , ,  �����  ����<  ����<  �����  �����      C  , ,   ����   ���t  ����t  �����   ����      C  , ,  n����  n���t  ���t  ����  n����      C  , ,  �����  ����t  f���t  f����  �����      C  , ,  

����  

���t  
����t  
�����  

����      C  , ,  X����  X���t  ���t  ����  X����      C  , ,  �����  ����t  P���t  P����  �����      C  , ,  �����  ����t  ����t  �����  �����      C  , ,  �����  ����G  ?���G  ?����  �����      C  , ,   ����*   �����  |����  |���*   ����*      C  , ,   ���*   ����  �����  ����*   ���*      C  , ,  n���*  n����  ����  ���*  n���*      C  , ,  ����*  �����  f����  f���*  ����*      C  , ,  

���*  

����  
�����  
����*  

���*      C  , ,  X���*  X����  ����  ���*  X���*      C  , ,  ����*  �����  P����  P���*  ����*      C  , ,  ����*  �����  �����  ����*  ����*      C  , ,  �����  ����G  	����G  	�����  �����      C  , ,  1����  1���G  ����G  �����  1����      C  , ,  ����  ���G  )���G  )����  ����      C  , ,  �����  ����G  w���G  w����  �����      C  , ,  �����  ����G  ����G  �����  �����      C  , ,   �����   ����D  |���D  |����   �����      C  , ,   ����2   �����  |����  |���2   ����2      C  , ,   ����b   ����  |���  |���b   ����b      C  , ,   �����   ����l  |���l  |����   �����      C  , ,   ����   ���l  ����l  �����   ����      C  , ,  n����  n���l  ���l  ����  n����      C  , ,  �����  ����l  f���l  f����  �����      C  , ,  

����  

���l  
����l  
�����  

����      C  , ,  X����  X���l  ���l  ����  X����      C  , ,  �����  ����l  P���l  P����  �����      C  , ,  �����  ����l  ����l  �����  �����      D   ,���D  !���D  ����*  ����*  !���D  !      D   ,���  !���  ����x  ����x  !���  !      D   ,����  !����  �����  �����  !����  !      D   ,���.  !���.  ����  ����  !���.  !      D   ,���|  !���|  ����b  ����b  !���|  !      D   ,����  !����  �����  �����  !����  !      D   ,���  !���  �����  �����  !���  !      D   ,���f  !���f  ����L  ����L  !���f  !      D   ,   �  !   �  �  �  �  �  !   �  !      D   ,    !    �  �  �  �  !    !      D   ,  P  !  P  �  6  �  6  !  P  !      D   ,  �  !  �  �  �  �  �  !  �  !      D   ,  	�  !  	�  �  
�  �  
�  !  	�  !      D   ,  :  !  :  �     �     !  :  !      D   ,  �  !  �  �  n  �  n  !  �  !      D   ,  �  !  �  �  �  �  �  !  �  !      D   ,���M   ����M  ����o  ����o   ����M   �      D   ,���   ����  ����  ����   ����   �      D   ,����   �����  ����  ����   �����   �      D   ,���7   ����7  ����Y  ����Y   ����7   �      D   ,����   �����  �����  �����   �����   �      D   ,����   �����  �����  �����   �����   �      D   ,���!   ����!  ����C  ����C   ����!   �      D   ,���o   ����o  �   �  �   �   ����o   �      D   ,  �   �  �  �  �  �  �   �  �   �      D   ,     �    �  -  �  -   �     �      D   ,  Y   �  Y  �  {  �  {   �  Y   �      D   ,  �   �  �  �  	�  �  	�   �  �   �      D   ,  
�   �  
�  �    �     �  
�   �      D   ,  C   �  C  �  e  �  e   �  C   �      D   ,  �   �  �  �  �  �  �   �  �   �      D   ,���M������M���e���o���e���o������M���      D   ,������������e������e������������      D   ,��������������e������e�������������      D   ,���7������7���e���Y���e���Y������7���      D   ,��������������e�������e��������������      D   ,��������������e�������e��������������      D   ,���!������!���e���C���e���C������!���      D   ,���o������o���e   ����e   �������o���      D   ,  ����  ����e  ����e  ����  ����      D   ,  ���  ���e  -���e  -���  ���      D   ,  Y���  Y���e  {���e  {���  Y���      D   ,  ����  ����e  	����e  	����  ����      D   ,  
����  
����e  ���e  ���  
����      D   ,  C���  C���e  e���e  e���  C���      D   ,  ����  ����e  ����e  ����  ����      D   ,���D���'���D�������*�������*���'���D���'      D   ,������'����������x�������x���'������'      D   ,�������'�����������������������'�������'      D   ,���.���'���.�����������������'���.���'      D   ,���|���'���|�������b�������b���'���|���'      D   ,�������'�����������������������'�������'      D   ,������'����������������������'������'      D   ,���f���'���f�������L�������L���'���f���'      D   ,   ����'   �����  �����  ����'   ����'      D   ,  ���'  ����  �����  ����'  ���'      D   ,  P���'  P����  6����  6���'  P���'      D   ,  ����'  �����  �����  ����'  ����'      D   ,  	����'  	�����  
�����  
����'  	����'      D   ,  :���'  :����   ����   ���'  :���'      D   ,  ����'  �����  n����  n���'  ����'      D   ,  ����'  �����  �����  ����'  ����'     �     "�     " &sky130_fd_pr__cap_mim_m3_1_BLS9H9     �   ,����������  @  "�  @  "������������      F   ,����������  @  %�  @  %������������      G   ,�������w����  �  �  �  ����w�������w      G   ,  #�����  #�    %�    %�����  #�����      F  , ,    �    �  �  �  �  �    �      F  , ,    d    ,  �  ,  �  d    d      F  , ,    �    �  �  �  �  �    �      F  , ,    D      �    �  D    D      F  , ,    �    |  �  |  �  �    �      F  , ,    $    �  �  �  �  $    $      F  , ,    �    \  �  \  �  �    �      F  , ,        �  �  �  �            F  , ,    t    <  �  <  �  t    t      F  , ,    �    �  �  �  �  �    �      F  , ,    T      �    �  T    T      F  , ,    	�    
�  �  
�  �  	�    	�      F  , ,    4    �  �  �  �  4    4      F  , ,    �    l  �  l  �  �    �      F  , ,        �  �  �  �            F  , ,    �    L  �  L  �  �    �      F  , ,    �    �  �  �  �  �    �      F  , ,     d    ,  �  ,  �   d     d      F  , ,  $�����  $�   d  %I   d  %I����  $�����      F  , ,  ����  ����  �����  �����  ����      F  , ,  ���D  ���  ����  ����D  ���D      F  , ,  ����  ���|  ����|  �����  ����      F  , ,  ���$  ����  �����  ����$  ���$      F  , ,  ����  ���\  ����\  �����  ����      F  , ,  ���  ����  �����  ����  ���      F  , ,  ���t  ���<  ����<  ����t  ���t      F  , ,  ����  ����  �����  �����  ����      F  , ,  ���T  ���  ����  ����T  ���T      F  , ,  ����  ���  ����  �����  ����      F  , ,  ���4  ����  �����  ����4  ���4      F  , ,  ���  ���l  ����l  ����  ���      F  , ,  ���  ����  �����  ����  ���      F  , ,  ���  ���L  ����L  ����  ���      F  , ,  ����  ���  ����  �����  ����      F  , ,  ���d  ���,  ����,  ����d  ���d      F  , ,  ����  ���  ����  �����  ����      F  , ,  ���D  ���  ����  ����D  ���D      F  , ,  �  t  �  <  f  <  f  t  �  t      F  , ,  .  t  .  <  �  <  �  t  .  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  N  t  N  <    <    t  N  t      F  , ,  �  t  �  <  	�  <  	�  t  �  t      F  , ,  
n  t  
n  <  6  <  6  t  
n  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  �  t  �  <  V  <  V  t  �  t      F  , ,    t    <  �  <  �  t    t      F  , ,  �  t  �  <  v  <  v  t  �  t      F  , ,  >  t  >  <    <    t  >  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  ^  t  ^  <  &  <  &  t  ^  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  ~  t  ~  <  F  <  F  t  ~  t      F  , ,    t    <  �  <  �  t    t      F  , ,  �  t  �  <  f  <  f  t  �  t      F  , ,  .  t  .  <  �  <  �  t  .  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  �  D  �    �    �  D  �  D      F  , ,  ~  D  ~    F    F  D  ~  D      F  , ,    D      �    �  D    D      F  , ,  �  D  �    f    f  D  �  D      F  , ,  .  D  .    �    �  D  .  D      F  , ,  �  D  �    �    �  D  �  D      F  , ,  $�  |  $�  D  %I  D  %I  |  $�  |      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  ^  �  ^  |  &  |  &  �  ^  �      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  ~  �  ~  |  F  |  F  �  ~  �      F  , ,    �    |  �  |  �  �    �      F  , ,  �  �  �  |  f  |  f  �  �  �      F  , ,  .  �  .  |  �  |  �  �  .  �      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  $�  �  $�  �  %I  �  %I  �  $�  �      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  ^  $  ^  �  &  �  &  $  ^  $      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  ~  $  ~  �  F  �  F  $  ~  $      F  , ,    $    �  �  �  �  $    $      F  , ,  �  $  �  �  f  �  f  $  �  $      F  , ,  .  $  .  �  �  �  �  $  .  $      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  $�  \  $�  $  %I  $  %I  \  $�  \      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  ^  �  ^  \  &  \  &  �  ^  �      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  ~  �  ~  \  F  \  F  �  ~  �      F  , ,    �    \  �  \  �  �    �      F  , ,  �  �  �  \  f  \  f  �  �  �      F  , ,  .  �  .  \  �  \  �  �  .  �      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  $�  �  $�  �  %I  �  %I  �  $�  �      F  , ,  �    �  �  �  �  �    �        F  , ,  ^    ^  �  &  �  &    ^        F  , ,  �    �  �  �  �  �    �        F  , ,  ~    ~  �  F  �  F    ~        F  , ,        �  �  �  �            F  , ,  �    �  �  f  �  f    �        F  , ,  .    .  �  �  �  �    .        F  , ,  �    �  �  �  �  �    �        F  , ,  $�  <  $�    %I    %I  <  $�  <      F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  ~  d  ~  ,  F  ,  F  d  ~  d      F  , ,    d    ,  �  ,  �  d    d      F  , ,  �  d  �  ,  f  ,  f  d  �  d      F  , ,  .  d  .  ,  �  ,  �  d  .  d      F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  $�  �  $�  d  %I  d  %I  �  $�  �      F  , ,  $�  L  $�    %I    %I  L  $�  L      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  ^  �  ^  �  &  �  &  �  ^  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  ~  �  ~  �  F  �  F  �  ~  �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  f  �  f  �  �  �      F  , ,  .  �  .  �  �  �  �  �  .  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  $�    $�  �  %I  �  %I    $�        F  , ,  �  D  �    �    �  D  �  D      F  , ,  ^  D  ^    &    &  D  ^  D      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  ^  �  ^  �  &  �  &  �  ^  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  ~  �  ~  �  F  �  F  �  ~  �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  f  �  f  �  �  �      F  , ,  .  �  .  �  �  �  �  �  .  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  $�  ,  $�  �  %I  �  %I  ,  $�  ,      F  , ,  $�  �  $�  �  %I  �  %I  �  $�  �      F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  ^  d  ^  ,  &  ,  &  d  ^  d      F  , ,  .  �  .  \  �  \  �  �  .  �      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  N  �  N  \    \    �  N  �      F  , ,  �  �  �  \  	�  \  	�  �  �  �      F  , ,  
n  �  
n  \  6  \  6  �  
n  �      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  �  �  �  \  V  \  V  �  �  �      F  , ,    �    \  �  \  �  �    �      F  , ,  �  �  �  \  v  \  v  �  �  �      F  , ,  >  �  >  \    \    �  >  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  N  �  N  �    �    �  N  �      F  , ,  �  �  �  �  	�  �  	�  �  �  �      F  , ,  
n  �  
n  �  6  �  6  �  
n  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  .  �  .  �  �  �  �  �  .  �      F  , ,  �  �  �  |  f  |  f  �  �  �      F  , ,  .  �  .  |  �  |  �  �  .  �      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  �  �  �  �  	�  �  	�  �  �  �      F  , ,  �    �  �  f  �  f    �        F  , ,  .    .  �  �  �  �    .        F  , ,  �    �  �  �  �  �    �        F  , ,  N    N  �    �      N        F  , ,  �    �  �  	�  �  	�    �        F  , ,  
n    
n  �  6  �  6    
n        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  V  �  V    �        F  , ,        �  �  �  �            F  , ,  �    �  �  v  �  v    �        F  , ,  >    >  �    �      >        F  , ,  N  �  N  |    |    �  N  �      F  , ,  �  �  �  |  	�  |  	�  �  �  �      F  , ,  
n  �  
n  |  6  |  6  �  
n  �      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  �  �  �  |  V  |  V  �  �  �      F  , ,    �    |  �  |  �  �    �      F  , ,  �  �  �  |  v  |  v  �  �  �      F  , ,  >  �  >  |    |    �  >  �      F  , ,  �  �  �  �  V  �  V  �  �  �      F  , ,  
n  �  
n  �  6  �  6  �  
n  �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  f  �  f  �  �  �      F  , ,  �  D  �    f    f  D  �  D      F  , ,  .  D  .    �    �  D  .  D      F  , ,  �  D  �    �    �  D  �  D      F  , ,  N  D  N          D  N  D      F  , ,  �  D  �    	�    	�  D  �  D      F  , ,  
n  D  
n    6    6  D  
n  D      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  $  �  �  f  �  f  $  �  $      F  , ,  .  $  .  �  �  �  �  $  .  $      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  N  $  N  �    �    $  N  $      F  , ,  �  $  �  �  	�  �  	�  $  �  $      F  , ,  
n  $  
n  �  6  �  6  $  
n  $      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  �  $  �  �  V  �  V  $  �  $      F  , ,    $    �  �  �  �  $    $      F  , ,  �  $  �  �  v  �  v  $  �  $      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  V  �  V  �  �  �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  v  �  v  �  �  �      F  , ,  >  �  >  �    �    �  >  �      F  , ,  >  $  >  �    �    $  >  $      F  , ,  �  D  �    �    �  D  �  D      F  , ,  �  D  �    V    V  D  �  D      F  , ,    D      �    �  D    D      F  , ,  �  D  �    v    v  D  �  D      F  , ,  >  D  >          D  >  D      F  , ,  �  �  �  �  v  �  v  �  �  �      F  , ,  >  �  >  �    �    �  >  �      F  , ,  �  �  �  �  f  �  f  �  �  �      F  , ,  .  �  .  �  �  �  �  �  .  �      F  , ,  �  d  �  ,  f  ,  f  d  �  d      F  , ,  .  d  .  ,  �  ,  �  d  .  d      F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  N  d  N  ,    ,    d  N  d      F  , ,  �  d  �  ,  	�  ,  	�  d  �  d      F  , ,  
n  d  
n  ,  6  ,  6  d  
n  d      F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  �  d  �  ,  V  ,  V  d  �  d      F  , ,    d    ,  �  ,  �  d    d      F  , ,  �  d  �  ,  v  ,  v  d  �  d      F  , ,  >  d  >  ,    ,    d  >  d      F  , ,  N  �  N  �    �    �  N  �      F  , ,  �  �  �  \  f  \  f  �  �  �      F  , ,  N  	�  N  
�    
�    	�  N  	�      F  , ,  �  	�  �  
�  	�  
�  	�  	�  �  	�      F  , ,  
n  	�  
n  
�  6  
�  6  	�  
n  	�      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  �  	�  �  
�  V  
�  V  	�  �  	�      F  , ,    	�    
�  �  
�  �  	�    	�      F  , ,  �  	�  �  
�  v  
�  v  	�  �  	�      F  , ,  >  	�  >  
�    
�    	�  >  	�      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  4  �  �  f  �  f  4  �  4      F  , ,  .  4  .  �  �  �  �  4  .  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  N  4  N  �    �    4  N  4      F  , ,  �  4  �  �  	�  �  	�  4  �  4      F  , ,  
n  4  
n  �  6  �  6  4  
n  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  �  4  �  �  V  �  V  4  �  4      F  , ,    4    �  �  �  �  4    4      F  , ,  �  4  �  �  v  �  v  4  �  4      F  , ,  >  4  >  �    �    4  >  4      F  , ,  N  �  N  �    �    �  N  �      F  , ,  �  �  �  l  f  l  f  �  �  �      F  , ,  .  �  .  l  �  l  �  �  .  �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  N  �  N  l    l    �  N  �      F  , ,  �  �  �  l  	�  l  	�  �  �  �      F  , ,  
n  �  
n  l  6  l  6  �  
n  �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  �  �  �  l  V  l  V  �  �  �      F  , ,    �    l  �  l  �  �    �      F  , ,  �  �  �  l  v  l  v  �  �  �      F  , ,  >  �  >  l    l    �  >  �      F  , ,  �  �  �  �  	�  �  	�  �  �  �      F  , ,  �    �  �  f  �  f    �        F  , ,  .    .  �  �  �  �    .        F  , ,  �    �  �  �  �  �    �        F  , ,  N    N  �    �      N        F  , ,  �    �  �  	�  �  	�    �        F  , ,  
n    
n  �  6  �  6    
n        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  V  �  V    �        F  , ,        �  �  �  �            F  , ,  �    �  �  v  �  v    �        F  , ,  >    >  �    �      >        F  , ,  
n  �  
n  �  6  �  6  �  
n  �      F  , ,  �  �  �  L  f  L  f  �  �  �      F  , ,  .  �  .  L  �  L  �  �  .  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  N  �  N  L    L    �  N  �      F  , ,  �  �  �  L  	�  L  	�  �  �  �      F  , ,  
n  �  
n  L  6  L  6  �  
n  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  �  �  �  L  V  L  V  �  �  �      F  , ,    �    L  �  L  �  �    �      F  , ,  �  �  �  L  v  L  v  �  �  �      F  , ,  >  �  >  L    L    �  >  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  f  �  f  �  �  �      F  , ,  .  �  .  �  �  �  �  �  .  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  N  �  N  �    �    �  N  �      F  , ,  �  �  �  �  	�  �  	�  �  �  �      F  , ,  
n  �  
n  �  6  �  6  �  
n  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  V  �  V  �  �  �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  v  �  v  �  �  �      F  , ,  >  �  >  �    �    �  >  �      F  , ,  �  �  �  �  V  �  V  �  �  �      F  , ,  �   d  �  ,  f  ,  f   d  �   d      F  , ,  .   d  .  ,  �  ,  �   d  .   d      F  , ,  �   d  �  ,  �  ,  �   d  �   d      F  , ,  N   d  N  ,    ,     d  N   d      F  , ,  �   d  �  ,  	�  ,  	�   d  �   d      F  , ,  
n   d  
n  ,  6  ,  6   d  
n   d      F  , ,  �   d  �  ,  �  ,  �   d  �   d      F  , ,  �   d  �  ,  V  ,  V   d  �   d      F  , ,     d    ,  �  ,  �   d     d      F  , ,  �   d  �  ,  v  ,  v   d  �   d      F  , ,  >   d  >  ,    ,     d  >   d      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  v  �  v  �  �  �      F  , ,  >  �  >  �    �    �  >  �      F  , ,  �  �  �  �  f  �  f  �  �  �      F  , ,  �  T  �    f    f  T  �  T      F  , ,  .  T  .    �    �  T  .  T      F  , ,  �  T  �    �    �  T  �  T      F  , ,  N  T  N          T  N  T      F  , ,  �  T  �    	�    	�  T  �  T      F  , ,  
n  T  
n    6    6  T  
n  T      F  , ,  �  T  �    �    �  T  �  T      F  , ,  �  T  �    V    V  T  �  T      F  , ,    T      �    �  T    T      F  , ,  �  T  �    v    v  T  �  T      F  , ,  >  T  >          T  >  T      F  , ,  .  �  .  �  �  �  �  �  .  �      F  , ,  �  	�  �  
�  f  
�  f  	�  �  	�      F  , ,  .  	�  .  
�  �  
�  �  	�  .  	�      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  ~  �  ~  �  F  �  F  �  ~  �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  f  �  f  �  �  �      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  ^  4  ^  �  &  �  &  4  ^  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  ~  4  ~  �  F  �  F  4  ~  4      F  , ,    4    �  �  �  �  4    4      F  , ,  �  4  �  �  f  �  f  4  �  4      F  , ,  .  4  .  �  �  �  �  4  .  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  ^  �  ^  L  &  L  &  �  ^  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  ~  �  ~  L  F  L  F  �  ~  �      F  , ,    �    L  �  L  �  �    �      F  , ,  �  �  �  L  f  L  f  �  �  �      F  , ,  .  �  .  L  �  L  �  �  .  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  $�  �  $�  �  %I  �  %I  �  $�  �      F  , ,  $�  l  $�  4  %I  4  %I  l  $�  l      F  , ,  .  �  .  �  �  �  �  �  .  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  $�    $�  �  %I  �  %I    $�        F  , ,  $�  �  $�  t  %I  t  %I  �  $�  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  T  �    �    �  T  �  T      F  , ,  ^  T  ^    &    &  T  ^  T      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  ^  	�  ^  
�  &  
�  &  	�  ^  	�      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  ~  	�  ~  
�  F  
�  F  	�  ~  	�      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  ^  �  ^  �  &  �  &  �  ^  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  ~  �  ~  �  F  �  F  �  ~  �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  f  �  f  �  �  �      F  , ,  .  �  .  �  �  �  �  �  .  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  $�  ,  $�  �  %I  �  %I  ,  $�  ,      F  , ,    	�    
�  �  
�  �  	�    	�      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  ^  �  ^  l  &  l  &  �  ^  �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  ~  �  ~  l  F  l  F  �  ~  �      F  , ,    �    l  �  l  �  �    �      F  , ,  �  �  �  l  f  l  f  �  �  �      F  , ,  .  �  .  l  �  l  �  �  .  �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  $�  �  $�  �  %I  �  %I  �  $�  �      F  , ,  �  	�  �  
�  f  
�  f  	�  �  	�      F  , ,  .  	�  .  
�  �  
�  �  	�  .  	�      F  , ,  �   d  �  ,  �  ,  �   d  �   d      F  , ,  ^   d  ^  ,  &  ,  &   d  ^   d      F  , ,  �   d  �  ,  �  ,  �   d  �   d      F  , ,  ~   d  ~  ,  F  ,  F   d  ~   d      F  , ,     d    ,  �  ,  �   d     d      F  , ,  �   d  �  ,  f  ,  f   d  �   d      F  , ,  .   d  .  ,  �  ,  �   d  .   d      F  , ,  �   d  �  ,  �  ,  �   d  �   d      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  $�  �  $�  	�  %I  	�  %I  �  $�  �      F  , ,  �  T  �    �    �  T  �  T      F  , ,  ~  T  ~    F    F  T  ~  T      F  , ,    T      �    �  T    T      F  , ,  �  T  �    f    f  T  �  T      F  , ,  .  T  .    �    �  T  .  T      F  , ,  �  T  �    �    �  T  �  T      F  , ,  $�  
�  $�  T  %I  T  %I  
�  $�  
�      F  , ,  ^  �  ^  �  &  �  &  �  ^  �      F  , ,  �    �  �  �  �  �    �        F  , ,  ^    ^  �  &  �  &    ^        F  , ,  �    �  �  �  �  �    �        F  , ,  ~    ~  �  F  �  F    ~        F  , ,        �  �  �  �            F  , ,  �    �  �  f  �  f    �        F  , ,  .    .  �  �  �  �    .        F  , ,  �    �  �  �  �  �    �        F  , ,  $�  L  $�    %I    %I  L  $�  L      F  , ,���  t���  <����  <����  t���  t      F  , ,��ޮ  t��ޮ  <���v  <���v  t��ޮ  t      F  , ,���>  t���>  <���  <���  t���>  t      F  , ,����  t����  <���  <���  t����  t      F  , ,���^  t���^  <���&  <���&  t���^  t      F  , ,����  t����  <���  <���  t����  t      F  , ,���~  t���~  <���F  <���F  t���~  t      F  , ,���  t���  <����  <����  t���  t      F  , ,���  t���  <���f  <���f  t���  t      F  , ,���.  t���.  <����  <����  t���.  t      F  , ,���  t���  <���  <���  t���  t      F  , ,���N  t���N  <���  <���  t���N  t      F  , ,����  t����  <���  <���  t����  t      F  , ,���n  t���n  <���6  <���6  t���n  t      F  , ,����  t����  <����  <����  t����  t      F  , ,���  t���  <���V  <���V  t���  t      F  , ,���  t���  <����  <����  t���  t      F  , ,����  t����  <���v  <���v  t����  t      F  , ,���>  t���>  <���  <���  t���>  t      F  , ,����  t����  <����  <����  t����  t      F  , ,���^  t���^  <���&  <���&  t���^  t      F  , ,����  t����  <����  <����  t����  t      F  , ,���~  t���~  <   F  <   F  t���~  t      F  , ,���  $���  �����  �����  $���  $      F  , ,����  $����  ����v  ����v  $����  $      F  , ,���>  $���>  ����  ����  $���>  $      F  , ,����  $����  �����  �����  $����  $      F  , ,���^  $���^  ����&  ����&  $���^  $      F  , ,����  $����  �����  �����  $����  $      F  , ,���~  $���~  �   F  �   F  $���~  $      F  , ,����  �����  ����v  ����v  �����  �      F  , ,���>  ����>  ����  ����  ����>  �      F  , ,����  �����  �����  �����  �����  �      F  , ,���^  ����^  ����&  ����&  ����^  �      F  , ,����  �����  �����  �����  �����  �      F  , ,���~  ����~  �   F  �   F  ����~  �      F  , ,����  �����  �����  �����  �����  �      F  , ,���^  ����^  ����&  ����&  ����^  �      F  , ,����  d����  ,���  ,���  d����  d      F  , ,����  �����  \���  \���  �����  �      F  , ,���n  ����n  \���6  \���6  ����n  �      F  , ,����  �����  \����  \����  �����  �      F  , ,���  ����  \���V  \���V  ����  �      F  , ,���  ����  \����  \����  ����  �      F  , ,����  �����  \���v  \���v  �����  �      F  , ,���>  ����>  \���  \���  ����>  �      F  , ,����  �����  \����  \����  �����  �      F  , ,���^  ����^  \���&  \���&  ����^  �      F  , ,����  �����  \����  \����  �����  �      F  , ,���~  ����~  \   F  \   F  ����~  �      F  , ,���n  d���n  ,���6  ,���6  d���n  d      F  , ,����  d����  ,����  ,����  d����  d      F  , ,���  d���  ,���V  ,���V  d���  d      F  , ,���  d���  ,����  ,����  d���  d      F  , ,����  d����  ,���v  ,���v  d����  d      F  , ,���>  d���>  ,���  ,���  d���>  d      F  , ,����  D����  ���  ���  D����  D      F  , ,���n  D���n  ���6  ���6  D���n  D      F  , ,����  D����  ����  ����  D����  D      F  , ,����  ����  ����  ����  ����        F  , ,���n  ���n  ����6  ����6  ���n        F  , ,����  ����  �����  �����  ����        F  , ,���  ���  ����V  ����V  ���        F  , ,���  ���  �����  �����  ���        F  , ,����  ����  ����v  ����v  ����        F  , ,���>  ���>  ����  ����  ���>        F  , ,����  ����  �����  �����  ����        F  , ,���^  ���^  ����&  ����&  ���^        F  , ,����  ����  �����  �����  ����        F  , ,���~  ���~  �   F  �   F  ���~        F  , ,���  D���  ���V  ���V  D���  D      F  , ,���  D���  ����  ����  D���  D      F  , ,����  D����  ���v  ���v  D����  D      F  , ,���>  D���>  ���  ���  D���>  D      F  , ,����  D����  ����  ����  D����  D      F  , ,���^  D���^  ���&  ���&  D���^  D      F  , ,����  D����  ����  ����  D����  D      F  , ,���~  D���~     F     F  D���~  D      F  , ,����  d����  ,����  ,����  d����  d      F  , ,���^  d���^  ,���&  ,���&  d���^  d      F  , ,����  d����  ,����  ,����  d����  d      F  , ,���~  d���~  ,   F  ,   F  d���~  d      F  , ,����  �����  �����  �����  �����  �      F  , ,���~  ����~  �   F  �   F  ����~  �      F  , ,���n  ����n  |���6  |���6  ����n  �      F  , ,����  �����  |����  |����  �����  �      F  , ,���  ����  |���V  |���V  ����  �      F  , ,���  ����  |����  |����  ����  �      F  , ,����  �����  |���v  |���v  �����  �      F  , ,���>  ����>  |���  |���  ����>  �      F  , ,����  �����  |����  |����  �����  �      F  , ,���^  ����^  |���&  |���&  ����^  �      F  , ,����  �����  |����  |����  �����  �      F  , ,���~  ����~  |   F  |   F  ����~  �      F  , ,���  ����  ����V  ����V  ����  �      F  , ,���  ����  �����  �����  ����  �      F  , ,����  �����  ����v  ����v  �����  �      F  , ,���>  ����>  ����  ����  ����>  �      F  , ,����  �����  ����  ����  �����  �      F  , ,���n  ����n  ����6  ����6  ����n  �      F  , ,����  �����  �����  �����  �����  �      F  , ,���  ����  ����V  ����V  ����  �      F  , ,���  ����  �����  �����  ����  �      F  , ,����  $����  ����  ����  $����  $      F  , ,���n  $���n  ����6  ����6  $���n  $      F  , ,����  $����  �����  �����  $����  $      F  , ,���  $���  ����V  ����V  $���  $      F  , ,����  �����  ����  ����  �����  �      F  , ,���n  ����n  ����6  ����6  ����n  �      F  , ,����  �����  �����  �����  �����  �      F  , ,����  �����  |���  |���  �����  �      F  , ,���  D���  ����  ����  D���  D      F  , ,���  D���  ���f  ���f  D���  D      F  , ,���.  D���.  ����  ����  D���.  D      F  , ,���  D���  ���  ���  D���  D      F  , ,���N  D���N  ���  ���  D���N  D      F  , ,��ޮ  $��ޮ  ����v  ����v  $��ޮ  $      F  , ,���>  $���>  ����  ����  $���>  $      F  , ,����  $����  ����  ����  $����  $      F  , ,���  ���  �����  �����  ���        F  , ,��ޮ  ��ޮ  ����v  ����v  ��ޮ        F  , ,���>  ���>  ����  ����  ���>        F  , ,����  ����  ����  ����  ����        F  , ,���^  ���^  ����&  ����&  ���^        F  , ,����  ����  ����  ����  ����        F  , ,���~  ���~  ����F  ����F  ���~        F  , ,���  ���  �����  �����  ���        F  , ,���  ���  ����f  ����f  ���        F  , ,���.  ���.  �����  �����  ���.        F  , ,���  ���  ����  ����  ���        F  , ,���N  ���N  ����  ����  ���N        F  , ,���^  $���^  ����&  ����&  $���^  $      F  , ,����  $����  ����  ����  $����  $      F  , ,���~  $���~  ����F  ����F  $���~  $      F  , ,���  d���  ,����  ,����  d���  d      F  , ,��ޮ  d��ޮ  ,���v  ,���v  d��ޮ  d      F  , ,���>  d���>  ,���  ,���  d���>  d      F  , ,����  d����  ,���  ,���  d����  d      F  , ,���^  d���^  ,���&  ,���&  d���^  d      F  , ,����  d����  ,���  ,���  d����  d      F  , ,���~  d���~  ,���F  ,���F  d���~  d      F  , ,���  d���  ,����  ,����  d���  d      F  , ,���  d���  ,���f  ,���f  d���  d      F  , ,���.  d���.  ,����  ,����  d���.  d      F  , ,���  d���  ,���  ,���  d���  d      F  , ,���N  d���N  ,���  ,���  d���N  d      F  , ,���  $���  �����  �����  $���  $      F  , ,���  ����  \����  \����  ����  �      F  , ,��ޮ  ���ޮ  \���v  \���v  ���ޮ  �      F  , ,���>  ����>  \���  \���  ����>  �      F  , ,����  �����  \���  \���  �����  �      F  , ,���^  ����^  \���&  \���&  ����^  �      F  , ,����  �����  \���  \���  �����  �      F  , ,���~  ����~  \���F  \���F  ����~  �      F  , ,���  ����  \����  \����  ����  �      F  , ,���  ����  \���f  \���f  ����  �      F  , ,���  ����  �����  �����  ����  �      F  , ,��ޮ  ���ޮ  ����v  ����v  ���ޮ  �      F  , ,���>  ����>  ����  ����  ����>  �      F  , ,����  �����  ����  ����  �����  �      F  , ,���^  ����^  ����&  ����&  ����^  �      F  , ,����  �����  ����  ����  �����  �      F  , ,���~  ����~  ����F  ����F  ����~  �      F  , ,���.  ����.  \����  \����  ����.  �      F  , ,���  ����  \���  \���  ����  �      F  , ,���N  ����N  \���  \���  ����N  �      F  , ,���  $���  ����f  ����f  $���  $      F  , ,���.  $���.  �����  �����  $���.  $      F  , ,���  $���  ����  ����  $���  $      F  , ,���N  $���N  ����  ����  $���N  $      F  , ,����  �����  ����  ����  �����  �      F  , ,���~  ����~  ����F  ����F  ����~  �      F  , ,���  ����  �����  �����  ����  �      F  , ,���  ����  ����f  ����f  ����  �      F  , ,���.  ����.  �����  �����  ����.  �      F  , ,���  ����  ����  ����  ����  �      F  , ,���N  ����N  ����  ����  ����N  �      F  , ,���  ����  �����  �����  ����  �      F  , ,��ޮ  ���ޮ  ����v  ����v  ���ޮ  �      F  , ,���>  ����>  ����  ����  ����>  �      F  , ,����  �����  ����  ����  �����  �      F  , ,���^  ����^  ����&  ����&  ����^  �      F  , ,���  $���  �����  �����  $���  $      F  , ,���  D���  ����  ����  D���  D      F  , ,��ޮ  D��ޮ  ���v  ���v  D��ޮ  D      F  , ,���>  D���>  ���  ���  D���>  D      F  , ,���  ����  �����  �����  ����  �      F  , ,���  ����  ����f  ����f  ����  �      F  , ,���.  ����.  �����  �����  ����.  �      F  , ,���  ����  ����  ����  ����  �      F  , ,���N  ����N  ����  ����  ����N  �      F  , ,����  D����  ���  ���  D����  D      F  , ,���^  D���^  ���&  ���&  D���^  D      F  , ,����  D����  ���  ���  D����  D      F  , ,���  ����  |����  |����  ����  �      F  , ,��ޮ  ���ޮ  |���v  |���v  ���ޮ  �      F  , ,���>  ����>  |���  |���  ����>  �      F  , ,����  �����  |���  |���  �����  �      F  , ,���^  ����^  |���&  |���&  ����^  �      F  , ,����  �����  |���  |���  �����  �      F  , ,���~  ����~  |���F  |���F  ����~  �      F  , ,���  ����  |����  |����  ����  �      F  , ,���  ����  |���f  |���f  ����  �      F  , ,���.  ����.  |����  |����  ����.  �      F  , ,���  ����  |���  |���  ����  �      F  , ,���N  ����N  |���  |���  ����N  �      F  , ,���~  D���~  ���F  ���F  D���~  D      F  , ,���.  T���.  ����  ����  T���.  T      F  , ,���  T���  ���  ���  T���  T      F  , ,���N  T���N  ���  ���  T���N  T      F  , ,���.  ����.  �����  �����  ����.  �      F  , ,���  ����  ����  ����  ����  �      F  , ,���N  ����N  ����  ����  ����N  �      F  , ,���~  ����~  ����F  ����F  ����~  �      F  , ,���  ����  �����  �����  ����  �      F  , ,���  ����  ����f  ����f  ����  �      F  , ,���~  4���~  ����F  ����F  4���~  4      F  , ,���  4���  �����  �����  4���  4      F  , ,���  4���  ����f  ����f  4���  4      F  , ,���.  4���.  �����  �����  4���.  4      F  , ,���  4���  ����  ����  4���  4      F  , ,���N  4���N  ����  ����  4���N  4      F  , ,���~  T���~  ���F  ���F  T���~  T      F  , ,���  T���  ����  ����  T���  T      F  , ,���  T���  ���f  ���f  T���  T      F  , ,���~  	����~  
����F  
����F  	����~  	�      F  , ,���  	����  
�����  
�����  	����  	�      F  , ,���  	����  
����f  
����f  	����  	�      F  , ,���.  	����.  
�����  
�����  	����.  	�      F  , ,���  	����  
����  
����  	����  	�      F  , ,���N  	����N  
����  
����  	����N  	�      F  , ,����  4����  ����  ����  4����  4      F  , ,���^  4���^  ����&  ����&  4���^  4      F  , ,����  4����  ����  ����  4����  4      F  , ,����  �����  ����  ����  �����  �      F  , ,���^  ����^  ����&  ����&  ����^  �      F  , ,����  �����  ����  ����  �����  �      F  , ,���  ����  �����  �����  ����  �      F  , ,��ޮ  ���ޮ  ����v  ����v  ���ޮ  �      F  , ,���>  ����>  ����  ����  ����>  �      F  , ,���  T���  ����  ����  T���  T      F  , ,��ޮ  T��ޮ  ���v  ���v  T��ޮ  T      F  , ,���>  T���>  ���  ���  T���>  T      F  , ,���  	����  
�����  
�����  	����  	�      F  , ,��ޮ  	���ޮ  
����v  
����v  	���ޮ  	�      F  , ,���>  	����>  
����  
����  	����>  	�      F  , ,����  	�����  
����  
����  	�����  	�      F  , ,���^  	����^  
����&  
����&  	����^  	�      F  , ,����  	�����  
����  
����  	�����  	�      F  , ,����  T����  ���  ���  T����  T      F  , ,���^  T���^  ���&  ���&  T���^  T      F  , ,����  T����  ���  ���  T����  T      F  , ,���  4���  �����  �����  4���  4      F  , ,��ޮ  4��ޮ  ����v  ����v  4��ޮ  4      F  , ,���>  4���>  ����  ����  4���>  4      F  , ,����  ����  ����  ����  ����        F  , ,���^  ���^  ����&  ����&  ���^        F  , ,����  ����  ����  ����  ����        F  , ,���  ����  �����  �����  ����  �      F  , ,��ޮ  ���ޮ  ����v  ����v  ���ޮ  �      F  , ,���>  ����>  ����  ����  ����>  �      F  , ,����  �����  ����  ����  �����  �      F  , ,���^  ����^  ����&  ����&  ����^  �      F  , ,����  �����  ����  ����  �����  �      F  , ,����  �����  l���  l���  �����  �      F  , ,���^  ����^  l���&  l���&  ����^  �      F  , ,����  �����  l���  l���  �����  �      F  , ,���  ����  l����  l����  ����  �      F  , ,��ޮ  ���ޮ  l���v  l���v  ���ޮ  �      F  , ,���>  ����>  l���  l���  ����>  �      F  , ,���  ���  �����  �����  ���        F  , ,��ޮ  ��ޮ  ����v  ����v  ��ޮ        F  , ,���>  ���>  ����  ����  ���>        F  , ,���   d���  ,����  ,����   d���   d      F  , ,��ޮ   d��ޮ  ,���v  ,���v   d��ޮ   d      F  , ,���>   d���>  ,���  ,���   d���>   d      F  , ,����   d����  ,���  ,���   d����   d      F  , ,���^   d���^  ,���&  ,���&   d���^   d      F  , ,����   d����  ,���  ,���   d����   d      F  , ,���  ����  L����  L����  ����  �      F  , ,��ޮ  ���ޮ  L���v  L���v  ���ޮ  �      F  , ,���>  ����>  L���  L���  ����>  �      F  , ,����  �����  L���  L���  �����  �      F  , ,���^  ����^  L���&  L���&  ����^  �      F  , ,����  �����  L���  L���  �����  �      F  , ,���.  ����.  L����  L����  ����.  �      F  , ,���  ����  L���  L���  ����  �      F  , ,���N  ����N  L���  L���  ����N  �      F  , ,���~  ����~  l���F  l���F  ����~  �      F  , ,���  ����  l����  l����  ����  �      F  , ,���  ����  l���f  l���f  ����  �      F  , ,���.  ����.  l����  l����  ����.  �      F  , ,���  ����  l���  l���  ����  �      F  , ,���N  ����N  l���  l���  ����N  �      F  , ,���~  ����~  ����F  ����F  ����~  �      F  , ,���  ����  �����  �����  ����  �      F  , ,���  ����  ����f  ����f  ����  �      F  , ,���~   d���~  ,���F  ,���F   d���~   d      F  , ,���   d���  ,����  ,����   d���   d      F  , ,���   d���  ,���f  ,���f   d���   d      F  , ,���.   d���.  ,����  ,����   d���.   d      F  , ,���   d���  ,���  ,���   d���   d      F  , ,���N   d���N  ,���  ,���   d���N   d      F  , ,���.  ����.  �����  �����  ����.  �      F  , ,���  ����  ����  ����  ����  �      F  , ,���N  ����N  ����  ����  ����N  �      F  , ,���~  ���~  ����F  ����F  ���~        F  , ,���  ���  �����  �����  ���        F  , ,���  ���  ����f  ����f  ���        F  , ,���.  ���.  �����  �����  ���.        F  , ,���  ���  ����  ����  ���        F  , ,���N  ���N  ����  ����  ���N        F  , ,���~  ����~  L���F  L���F  ����~  �      F  , ,���  ����  L����  L����  ����  �      F  , ,���  ����  L���f  L���f  ����  �      F  , ,���>  ���>  ����  ����  ���>        F  , ,����  ����  �����  �����  ����        F  , ,���^  ���^  ����&  ����&  ���^        F  , ,����  ����  �����  �����  ����        F  , ,���~  ���~  �   F  �   F  ���~        F  , ,����  �����  ����  ����  �����  �      F  , ,���n  ����n  ����6  ����6  ����n  �      F  , ,����  �����  �����  �����  �����  �      F  , ,���  ����  ����V  ����V  ����  �      F  , ,���  ����  �����  �����  ����  �      F  , ,����  �����  ����v  ����v  �����  �      F  , ,���>  ����>  ����  ����  ����>  �      F  , ,����  �����  �����  �����  �����  �      F  , ,���^  ����^  ����&  ����&  ����^  �      F  , ,����  �����  �����  �����  �����  �      F  , ,���~  ����~  �   F  �   F  ����~  �      F  , ,����  	�����  
����  
����  	�����  	�      F  , ,���n  	����n  
����6  
����6  	����n  	�      F  , ,����  	�����  
�����  
�����  	�����  	�      F  , ,���  	����  
����V  
����V  	����  	�      F  , ,���  	����  
�����  
�����  	����  	�      F  , ,����  	�����  
����v  
����v  	�����  	�      F  , ,���>  	����>  
����  
����  	����>  	�      F  , ,����  	�����  
�����  
�����  	�����  	�      F  , ,���^  	����^  
����&  
����&  	����^  	�      F  , ,����  	�����  
�����  
�����  	�����  	�      F  , ,���~  	����~  
�   F  
�   F  	����~  	�      F  , ,����  �����  l���  l���  �����  �      F  , ,���n  ����n  l���6  l���6  ����n  �      F  , ,����  �����  l����  l����  �����  �      F  , ,���  ����  l���V  l���V  ����  �      F  , ,���  ����  l����  l����  ����  �      F  , ,����  �����  l���v  l���v  �����  �      F  , ,���>  ����>  l���  l���  ����>  �      F  , ,����  �����  l����  l����  �����  �      F  , ,���^  ����^  l���&  l���&  ����^  �      F  , ,����  �����  l����  l����  �����  �      F  , ,���~  ����~  l   F  l   F  ����~  �      F  , ,����  4����  ����  ����  4����  4      F  , ,���n  4���n  ����6  ����6  4���n  4      F  , ,����  4����  �����  �����  4����  4      F  , ,���  4���  ����V  ����V  4���  4      F  , ,���  4���  �����  �����  4���  4      F  , ,����  4����  ����v  ����v  4����  4      F  , ,���>  4���>  ����  ����  4���>  4      F  , ,����  4����  �����  �����  4����  4      F  , ,���^  4���^  ����&  ����&  4���^  4      F  , ,����  4����  �����  �����  4����  4      F  , ,���~  4���~  �   F  �   F  4���~  4      F  , ,����   d����  ,���  ,���   d����   d      F  , ,���n   d���n  ,���6  ,���6   d���n   d      F  , ,����   d����  ,����  ,����   d����   d      F  , ,���   d���  ,���V  ,���V   d���   d      F  , ,���   d���  ,����  ,����   d���   d      F  , ,����   d����  ,���v  ,���v   d����   d      F  , ,���>   d���>  ,���  ,���   d���>   d      F  , ,����   d����  ,����  ,����   d����   d      F  , ,���^   d���^  ,���&  ,���&   d���^   d      F  , ,����   d����  ,����  ,����   d����   d      F  , ,���~   d���~  ,   F  ,   F   d���~   d      F  , ,����  �����  L���  L���  �����  �      F  , ,���n  ����n  L���6  L���6  ����n  �      F  , ,����  �����  L����  L����  �����  �      F  , ,���  ����  L���V  L���V  ����  �      F  , ,���  ����  L����  L����  ����  �      F  , ,����  �����  L���v  L���v  �����  �      F  , ,���>  ����>  L���  L���  ����>  �      F  , ,����  �����  L����  L����  �����  �      F  , ,���^  ����^  L���&  L���&  ����^  �      F  , ,����  �����  L����  L����  �����  �      F  , ,���~  ����~  L   F  L   F  ����~  �      F  , ,����  T����  ���  ���  T����  T      F  , ,���n  T���n  ���6  ���6  T���n  T      F  , ,����  T����  ����  ����  T����  T      F  , ,���  T���  ���V  ���V  T���  T      F  , ,���  T���  ����  ����  T���  T      F  , ,����  T����  ���v  ���v  T����  T      F  , ,���>  T���>  ���  ���  T���>  T      F  , ,����  T����  ����  ����  T����  T      F  , ,���^  T���^  ���&  ���&  T���^  T      F  , ,����  T����  ����  ����  T����  T      F  , ,���~  T���~     F     F  T���~  T      F  , ,����  �����  ����  ����  �����  �      F  , ,���n  ����n  ����6  ����6  ����n  �      F  , ,����  �����  �����  �����  �����  �      F  , ,���  ����  ����V  ����V  ����  �      F  , ,���  ����  �����  �����  ����  �      F  , ,����  �����  ����v  ����v  �����  �      F  , ,���>  ����>  ����  ����  ����>  �      F  , ,����  �����  �����  �����  �����  �      F  , ,���^  ����^  ����&  ����&  ����^  �      F  , ,����  �����  �����  �����  �����  �      F  , ,���~  ����~  �   F  �   F  ����~  �      F  , ,����  ����  ����  ����  ����        F  , ,���n  ���n  ����6  ����6  ���n        F  , ,����  ����  �����  �����  ����        F  , ,���  ���  ����V  ����V  ���        F  , ,���  ���  �����  �����  ���        F  , ,����  ����  ����v  ����v  ����        F  , ,�����������������������������������      F  , ,��ޮ������ޮ������v������v������ޮ����      F  , ,���>�������>�������������������>����      F  , ,������������������������������������      F  , ,���^�������^������&������&�������^����      F  , ,������������������������������������      F  , ,���~�������~������F������F�������~����      F  , ,�����������������������������������      F  , ,����������������f������f�����������      F  , ,���.�������.���������������������.����      F  , ,���������������������������������      F  , ,���N�������N�������������������N����      F  , ,������������������������������������      F  , ,���n�������n������6������6�������n����      F  , ,��������������������������������������      F  , ,����������������V������V�����������      F  , ,�����������������������������������      F  , ,������������������v������v������������      F  , ,���>�������>�������������������>����      F  , ,��������������������������������������      F  , ,���^�������^������&������&�������^����      F  , ,��������������������������������������      F  , ,���~�������~���   F���   F�������~����      F  , ,���������������|�������|����������������      F  , ,���^�������^���|���&���|���&�������^����      F  , ,���������������|�������|����������������      F  , ,���~�������~���|   F���|   F�������~����      F  , ,�������$���������������������$�������$      F  , ,���n���$���n�������6�������6���$���n���$      F  , ,�������$�����������������������$�������$      F  , ,������$����������V�������V���$������$      F  , ,������$����������������������$������$      F  , ,�������$�����������v�������v���$�������$      F  , ,���>���$���>�����������������$���>���$      F  , ,�������$�����������������������$�������$      F  , ,���^���$���^�������&�������&���$���^���$      F  , ,�������$�����������������������$�������$      F  , ,���~���$���~����   F����   F���$���~���$      F  , ,���������������\������\���������������      F  , ,���n�������n���\���6���\���6�������n����      F  , ,���������������\�������\����������������      F  , ,�������������\���V���\���V�����������      F  , ,�������������\�������\���������������      F  , ,���������������\���v���\���v������������      F  , ,���>�������>���\������\����������>����      F  , ,���������������\�������\����������������      F  , ,���^�������^���\���&���\���&�������^����      F  , ,���������������\�������\����������������      F  , ,���~�������~���\   F���\   F�������~����      F  , ,�����������������������������������      F  , ,���n������n�������6�������6������n���      F  , ,�������������������������������������      F  , ,����������������V�������V���������      F  , ,����������������������������������      F  , ,������������������v�������v����������      F  , ,���>������>��������������������>���      F  , ,�������������������������������������      F  , ,���^������^�������&�������&������^���      F  , ,�������������������������������������      F  , ,���~������~����   F����   F������~���      F  , ,�������t�������<������<������t�������t      F  , ,���n���t���n���<���6���<���6���t���n���t      F  , ,�������t�������<�������<�������t�������t      F  , ,������t������<���V���<���V���t������t      F  , ,������t������<�������<�������t������t      F  , ,�������t�������<���v���<���v���t�������t      F  , ,���>���t���>���<������<������t���>���t      F  , ,�������t�������<�������<�������t�������t      F  , ,���^���t���^���<���&���<���&���t���^���t      F  , ,�������t�������<�������<�������t�������t      F  , ,���~���t���~���<   F���<   F���t���~���t      F  , ,��������������������������������������      F  , ,���n�������n�������6�������6�������n����      F  , ,����������������������������������������      F  , ,�����������������V�������V�����������      F  , ,�������������������������������������      F  , ,�������������������v�������v������������      F  , ,���>�������>���������������������>����      F  , ,����������������������������������������      F  , ,���^�������^�������&�������&�������^����      F  , ,����������������������������������������      F  , ,���~�������~����   F����   F�������~����      F  , ,�������T�������������������T�������T      F  , ,���n���T���n������6������6���T���n���T      F  , ,�������T���������������������T�������T      F  , ,������T���������V������V���T������T      F  , ,������T��������������������T������T      F  , ,�������T����������v������v���T�������T      F  , ,���>���T���>���������������T���>���T      F  , ,�������T���������������������T�������T      F  , ,���^���T���^������&������&���T���^���T      F  , ,�������T���������������������T�������T      F  , ,���~���T���~���   F���   F���T���~���T      F  , ,���>�������>���������������������>����      F  , ,����������������������������������������      F  , ,���^�������^�������&�������&�������^����      F  , ,����������������������������������������      F  , ,���~�������~����   F����   F�������~����      F  , ,�������D�������������������D�������D      F  , ,���n���D���n������6������6���D���n���D      F  , ,�������D���������������������D�������D      F  , ,������D���������V������V���D������D      F  , ,������D��������������������D������D      F  , ,�������D����������v������v���D�������D      F  , ,���>���D���>���������������D���>���D      F  , ,�������D���������������������D�������D      F  , ,���^���D���^������&������&���D���^���D      F  , ,�������D���������������������D�������D      F  , ,���~���D���~���   F���   F���D���~���D      F  , ,���������������|������|���������������      F  , ,���n�������n���|���6���|���6�������n����      F  , ,���������������|�������|����������������      F  , ,�������������|���V���|���V�����������      F  , ,�������������|�������|���������������      F  , ,���������������|���v���|���v������������      F  , ,���>�������>���|������|����������>����      F  , ,��������������������������������������      F  , ,���n�������n�������6�������6�������n����      F  , ,����������������������������������������      F  , ,�����������������V�������V�����������      F  , ,�������������������������������������      F  , ,�������������������v�������v������������      F  , ,���~���$���~�������F�������F���$���~���$      F  , ,������$����������������������$������$      F  , ,������$����������f�������f���$������$      F  , ,���.���$���.�������������������$���.���$      F  , ,������$��������������������$������$      F  , ,���N���$���N�����������������$���N���$      F  , ,������D���������f������f���D������D      F  , ,���.���D���.�����������������D���.���D      F  , ,���~�������~�������F�������F�������~����      F  , ,���~�������~���|���F���|���F�������~����      F  , ,�������������|�������|���������������      F  , ,�������������������������������������      F  , ,���~�������~���\���F���\���F�������~����      F  , ,�������������\�������\���������������      F  , ,�������������\���f���\���f�����������      F  , ,���.�������.���\�������\�����������.����      F  , ,�������������\������\��������������      F  , ,���N�������N���\������\����������N����      F  , ,�������������|���f���|���f�����������      F  , ,���.�������.���|�������|�����������.����      F  , ,�������������|������|��������������      F  , ,�����������������f�������f�����������      F  , ,���N�������N���|������|����������N����      F  , ,������D������������������D������D      F  , ,���N���D���N���������������D���N���D      F  , ,���.�������.�����������������������.����      F  , ,�����������������������������������      F  , ,���N�������N���������������������N����      F  , ,���~���D���~������F������F���D���~���D      F  , ,������D��������������������D������D      F  , ,��ޮ������ޮ�������v�������v������ޮ����      F  , ,�������������|�������|���������������      F  , ,��ޮ������ޮ���|���v���|���v������ޮ����      F  , ,�������$���������������������$�������$      F  , ,���>�������>���|������|����������>����      F  , ,���������������|������|���������������      F  , ,���^�������^���|���&���|���&�������^����      F  , ,���������������|������|���������������      F  , ,���^���$���^�������&�������&���$���^���$      F  , ,�������$���������������������$�������$      F  , ,��������������������������������������      F  , ,�������������\�������\���������������      F  , ,��ޮ������ޮ���\���v���\���v������ޮ����      F  , ,�������������������������������������      F  , ,������D��������������������D������D      F  , ,��ޮ���D��ޮ������v������v���D��ޮ���D      F  , ,���>���D���>���������������D���>���D      F  , ,�������D�������������������D�������D      F  , ,���^�������^�������&�������&�������^����      F  , ,���^���D���^������&������&���D���^���D      F  , ,�������D�������������������D�������D      F  , ,���>�������>���\������\����������>����      F  , ,���������������\������\���������������      F  , ,��������������������������������������      F  , ,���^�������^���\���&���\���&�������^����      F  , ,���������������\������\���������������      F  , ,���>�������>���������������������>����      F  , ,������$����������������������$������$      F  , ,��ޮ���$��ޮ�������v�������v���$��ޮ���$      F  , ,���>���$���>�����������������$���>���$      F  , ,���>���T���>���������������T���>���T      F  , ,�������T�������������������T�������T      F  , ,���^���T���^������&������&���T���^���T      F  , ,�������T�������������������T�������T      F  , ,������t������<�������<�������t������t      F  , ,��ޮ���t��ޮ���<���v���<���v���t��ޮ���t      F  , ,���>���t���>���<������<������t���>���t      F  , ,����������������������������������      F  , ,��ޮ�����ޮ�������v�������v�����ޮ���      F  , ,���>������>��������������������>���      F  , ,�����������������������������������      F  , ,���^������^�������&�������&������^���      F  , ,�����������������������������������      F  , ,�������t�������<������<������t�������t      F  , ,���^���t���^���<���&���<���&���t���^���t      F  , ,�������t�������<������<������t�������t      F  , ,�������������������������������������      F  , ,��ޮ������ޮ�������v�������v������ޮ����      F  , ,���>�������>���������������������>����      F  , ,��������������������������������������      F  , ,���^�������^�������&�������&�������^����      F  , ,��������������������������������������      F  , ,������T��������������������T������T      F  , ,��ޮ���T��ޮ������v������v���T��ޮ���T      F  , ,�����������������f�������f�����������      F  , ,���.�������.�����������������������.����      F  , ,�����������������������������������      F  , ,���N�������N���������������������N����      F  , ,���~���t���~���<���F���<���F���t���~���t      F  , ,������t������<�������<�������t������t      F  , ,������t������<���f���<���f���t������t      F  , ,���~������~�������F�������F������~���      F  , ,����������������������������������      F  , ,����������������f�������f���������      F  , ,���.������.����������������������.���      F  , ,��������������������������������      F  , ,���N������N��������������������N���      F  , ,���.���t���.���<�������<�������t���.���t      F  , ,������t������<������<������t������t      F  , ,���N���t���N���<������<������t���N���t      F  , ,���~���T���~������F������F���T���~���T      F  , ,������T��������������������T������T      F  , ,������T���������f������f���T������T      F  , ,���.���T���.�����������������T���.���T      F  , ,������T������������������T������T      F  , ,���N���T���N���������������T���N���T      F  , ,���~�������~�������F�������F�������~����      F  , ,�������������������������������������      F  , ,������4����������f�������f���4������4      F  , ,���.���4���.�������������������4���.���4      F  , ,������4��������������������4������4      F  , ,���N���4���N�����������������4���N���4      F  , ,������4����������������������4������4      F  , ,������������l�������l�������������      F  , ,��ޮ�����ޮ���l���v���l���v�����ޮ���      F  , ,���>������>���l������l���������>���      F  , ,��������������l������l�������������      F  , ,���^������^���l���&���l���&������^���      F  , ,��������������l������l�������������      F  , ,���~������~���l���F���l���F������~���      F  , ,������������l�������l�������������      F  , ,������������l���f���l���f���������      F  , ,���.������.���l�������l����������.���      F  , ,������������l������l������������      F  , ,���N������N���l������l���������N���      F  , ,��ޮ���4��ޮ�������v�������v���4��ޮ���4      F  , ,����������������������������������      F  , ,��ޮ�����ޮ�������v�������v�����ޮ���      F  , ,���>������>��������������������>���      F  , ,�����������������������������������      F  , ,���^������^�������&�������&������^���      F  , ,�����������������������������������      F  , ,���~������~�������F�������F������~���      F  , ,����������������������������������      F  , ,����������������f�������f���������      F  , ,���.������.����������������������.���      F  , ,��������������������������������      F  , ,���N������N��������������������N���      F  , ,���>���4���>�����������������4���>���4      F  , ,������������L�������L�������������      F  , ,��ޮ�����ޮ���L���v���L���v�����ޮ���      F  , ,���>������>���L������L���������>���      F  , ,��������������L������L�������������      F  , ,���^������^���L���&���L���&������^���      F  , ,��������������L������L�������������      F  , ,���~������~���L���F���L���F������~���      F  , ,������������L�������L�������������      F  , ,������������L���f���L���f���������      F  , ,���.������.���L�������L����������.���      F  , ,������������L������L������������      F  , ,���N������N���L������L���������N���      F  , ,�������4���������������������4�������4      F  , ,�����������������������������������      F  , ,��ޮ������ޮ������v������v������ޮ����      F  , ,���>�������>�������������������>����      F  , ,������������������������������������      F  , ,���^�������^������&������&�������^����      F  , ,������������������������������������      F  , ,���~�������~������F������F�������~����      F  , ,�����������������������������������      F  , ,����������������f������f�����������      F  , ,���.�������.���������������������.����      F  , ,���������������������������������      F  , ,���N�������N�������������������N����      F  , ,���^���4���^�������&�������&���4���^���4      F  , ,������d������,�������,�������d������d      F  , ,��ޮ���d��ޮ���,���v���,���v���d��ޮ���d      F  , ,���>���d���>���,������,������d���>���d      F  , ,�������d�������,������,������d�������d      F  , ,���^���d���^���,���&���,���&���d���^���d      F  , ,�������d�������,������,������d�������d      F  , ,���~���d���~���,���F���,���F���d���~���d      F  , ,������d������,�������,�������d������d      F  , ,������d������,���f���,���f���d������d      F  , ,���.���d���.���,�������,�������d���.���d      F  , ,������d������,������,������d������d      F  , ,���N���d���N���,������,������d���N���d      F  , ,�������4���������������������4�������4      F  , ,�����������������������������������      F  , ,��ޮ������ޮ������v������v������ޮ����      F  , ,���>�������>�������������������>����      F  , ,������������������������������������      F  , ,���^�������^������&������&�������^����      F  , ,������������������������������������      F  , ,���~�������~������F������F�������~����      F  , ,�����������������������������������      F  , ,����������������f������f�����������      F  , ,���.�������.���������������������.����      F  , ,���������������������������������      F  , ,���N�������N�������������������N����      F  , ,���~���4���~�������F�������F���4���~���4      F  , ,������D��������������������D������D      F  , ,��ޮ���D��ޮ������v������v���D��ޮ���D      F  , ,���>���D���>���������������D���>���D      F  , ,�������D�������������������D�������D      F  , ,���^���D���^������&������&���D���^���D      F  , ,�������D�������������������D�������D      F  , ,���~���D���~������F������F���D���~���D      F  , ,������D��������������������D������D      F  , ,������D���������f������f���D������D      F  , ,���.���D���.�����������������D���.���D      F  , ,������D������������������D������D      F  , ,���N���D���N���������������D���N���D      F  , ,������4����������������������4������4      F  , ,�����������������������������������      F  , ,���n������n�������6�������6������n���      F  , ,�������������������������������������      F  , ,����������������V�������V���������      F  , ,������������������������������������      F  , ,���n�������n������6������6�������n����      F  , ,��������������������������������������      F  , ,����������������V������V�����������      F  , ,�����������������������������������      F  , ,������������������v������v������������      F  , ,���>�������>�������������������>����      F  , ,��������������������������������������      F  , ,���^�������^������&������&�������^����      F  , ,��������������������������������������      F  , ,���~�������~���   F���   F�������~����      F  , ,����������������������������������      F  , ,������������������v�������v����������      F  , ,���>������>��������������������>���      F  , ,�������������������������������������      F  , ,���^������^�������&�������&������^���      F  , ,�������������������������������������      F  , ,���~������~����   F����   F������~���      F  , ,��������������l�������l��������������      F  , ,������������l���V���l���V���������      F  , ,������������l�������l�������������      F  , ,��������������l���v���l���v����������      F  , ,���>������>���l������l���������>���      F  , ,��������������l�������l��������������      F  , ,�������d�������,������,������d�������d      F  , ,���n���d���n���,���6���,���6���d���n���d      F  , ,�������d�������,�������,�������d�������d      F  , ,������d������,���V���,���V���d������d      F  , ,������d������,�������,�������d������d      F  , ,�������d�������,���v���,���v���d�������d      F  , ,���>���d���>���,������,������d���>���d      F  , ,�������d�������,�������,�������d�������d      F  , ,���^���d���^���,���&���,���&���d���^���d      F  , ,�������d�������,�������,�������d�������d      F  , ,���~���d���~���,   F���,   F���d���~���d      F  , ,���^������^���l���&���l���&������^���      F  , ,��������������l�������l��������������      F  , ,���~������~���l   F���l   F������~���      F  , ,�������4�����������������������4�������4      F  , ,������4����������V�������V���4������4      F  , ,������4����������������������4������4      F  , ,�������4�����������v�������v���4�������4      F  , ,��������������L������L�������������      F  , ,���n������n���L���6���L���6������n���      F  , ,��������������L�������L��������������      F  , ,������������L���V���L���V���������      F  , ,������������L�������L�������������      F  , ,��������������L���v���L���v����������      F  , ,������������������������������������      F  , ,���n�������n������6������6�������n����      F  , ,��������������������������������������      F  , ,����������������V������V�����������      F  , ,�����������������������������������      F  , ,������������������v������v������������      F  , ,���>�������>�������������������>����      F  , ,��������������������������������������      F  , ,���^�������^������&������&�������^����      F  , ,��������������������������������������      F  , ,���~�������~���   F���   F�������~����      F  , ,���>������>���L������L���������>���      F  , ,��������������L�������L��������������      F  , ,���^������^���L���&���L���&������^���      F  , ,��������������L�������L��������������      F  , ,���~������~���L   F���L   F������~���      F  , ,���>���4���>�����������������4���>���4      F  , ,�������4�����������������������4�������4      F  , ,���^���4���^�������&�������&���4���^���4      F  , ,�������4�����������������������4�������4      F  , ,���~���4���~����   F����   F���4���~���4      F  , ,�������4���������������������4�������4      F  , ,���n���4���n�������6�������6���4���n���4      F  , ,��������������l������l�������������      F  , ,�������D�������������������D�������D      F  , ,���n���D���n������6������6���D���n���D      F  , ,�������D���������������������D�������D      F  , ,������D���������V������V���D������D      F  , ,������D��������������������D������D      F  , ,�������D����������v������v���D�������D      F  , ,���>���D���>���������������D���>���D      F  , ,�������D���������������������D�������D      F  , ,���^���D���^������&������&���D���^���D      F  , ,�������D���������������������D�������D      F  , ,���~���D���~���   F���   F���D���~���D      F  , ,���n������n���l���6���l���6������n���      F  , ,  ^����  ^���  &���  &����  ^����      F  , ,  �����  ����  ����  �����  �����      F  , ,  ~����  ~���  F���  F����  ~����      F  , ,  ����  ���  ����  �����  ����      F  , ,  �����  ����  f���  f����  �����      F  , ,  .����  .���  ����  �����  .����      F  , ,  �����  ����  ����  �����  �����      F  , ,  �����  ����  f���  f����  �����      F  , ,  .����  .���  ����  �����  .����      F  , ,  �����  ����  ����  �����  �����      F  , ,  N����  N���  ���  ����  N����      F  , ,  �����  ����  	����  	�����  �����      F  , ,  
n����  
n���  6���  6����  
n����      F  , ,  �����  ����  ����  �����  �����      F  , ,  �����  ����  V���  V����  �����      F  , ,  ����  ���  ����  �����  ����      F  , ,  �����  ����  v���  v����  �����      F  , ,  >����  >���  ���  ����  >����      F  , ,  �����  ����  ����  �����  �����      F  , ,  $����<  $����  %I���  %I���<  $����<      F  , ,  ����D  ����  f���  f���D  ����D      F  , ,  .���D  .���  ����  ����D  .���D      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  $����|  $����D  %I���D  %I���|  $����|      F  , ,  �����  �����  �����  �����  �����      F  , ,  ����$  �����  �����  ����$  ����$      F  , ,  ����t  ����<  ����<  ����t  ����t      F  , ,  ^���t  ^���<  &���<  &���t  ^���t      F  , ,  ����t  ����<  ����<  ����t  ����t      F  , ,  ~���t  ~���<  F���<  F���t  ~���t      F  , ,  ���t  ���<  ����<  ����t  ���t      F  , ,  ����t  ����<  f���<  f���t  ����t      F  , ,  .���t  .���<  ����<  ����t  .���t      F  , ,  ����t  ����<  ����<  ����t  ����t      F  , ,  $�����  $����t  %I���t  %I����  $�����      F  , ,  ^���$  ^����  &����  &���$  ^���$      F  , ,  ����$  �����  �����  ����$  ����$      F  , ,  ~���$  ~����  F����  F���$  ~���$      F  , ,  ���$  ����  �����  ����$  ���$      F  , ,  ����$  �����  f����  f���$  ����$      F  , ,  .���$  .����  �����  ����$  .���$      F  , ,  ����$  �����  �����  ����$  ����$      F  , ,  $����\  $����$  %I���$  %I���\  $����\      F  , ,  ^����  ^����  &����  &����  ^����      F  , ,  �����  �����  �����  �����  �����      F  , ,  ~����  ~����  F����  F����  ~����      F  , ,  ����  ����  �����  �����  ����      F  , ,  �����  �����  f����  f����  �����      F  , ,  .����  .����  �����  �����  .����      F  , ,  �����  �����  �����  �����  �����      F  , ,  $����  $�����  %I����  %I���  $����      F  , ,  �����  �����  �����  �����  �����      F  , ,  ^����  ^����  &����  &����  ^����      F  , ,  �����  �����  �����  �����  �����      F  , ,  ~����  ~����  F����  F����  ~����      F  , ,  ����  ����  �����  �����  ����      F  , ,  �����  �����  f����  f����  �����      F  , ,  .����  .����  �����  �����  .����      F  , ,  �����  �����  �����  �����  �����      F  , ,  $����  $�����  %I����  %I���  $����      F  , ,  �����  ����\  ����\  �����  �����      F  , ,  ^����  ^���\  &���\  &����  ^����      F  , ,  �����  ����\  ����\  �����  �����      F  , ,  ~����  ~���\  F���\  F����  ~����      F  , ,  ����  ���\  ����\  �����  ����      F  , ,  ����T  ����  ����  ����T  ����T      F  , ,  ^���T  ^���  &���  &���T  ^���T      F  , ,  ����T  ����  ����  ����T  ����T      F  , ,  ~���T  ~���  F���  F���T  ~���T      F  , ,  ���T  ���  ����  ����T  ���T      F  , ,  ����T  ����  f���  f���T  ����T      F  , ,  .���T  .���  ����  ����T  .���T      F  , ,  ����T  ����  ����  ����T  ����T      F  , ,  $����  $����T  %I���T  %I���  $����      F  , ,  �����  ����\  f���\  f����  �����      F  , ,  .����  .���\  ����\  �����  .����      F  , ,  �����  ����\  ����\  �����  �����      F  , ,  $�����  $�����  %I����  %I����  $�����      F  , ,  �����  ����|  ����|  �����  �����      F  , ,  ^����  ^���|  &���|  &����  ^����      F  , ,  �����  ����|  ����|  �����  �����      F  , ,  ~����  ~���|  F���|  F����  ~����      F  , ,  ����  ���|  ����|  �����  ����      F  , ,  �����  ����|  f���|  f����  �����      F  , ,  .����  .���|  ����|  �����  .����      F  , ,  �����  ����|  ����|  �����  �����      F  , ,  $�����  $�����  %I����  %I����  $�����      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  ^���D  ^���  &���  &���D  ^���D      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  ~���D  ~���  F���  F���D  ~���D      F  , ,  ���D  ���  ����  ����D  ���D      F  , ,  ����  �����  �����  ����  ����      F  , ,  ^���  ^����  &����  &���  ^���      F  , ,  ����  �����  �����  ����  ����      F  , ,  ~���  ~����  F����  F���  ~���      F  , ,  ���  ����  �����  ����  ���      F  , ,  ����  �����  f����  f���  ����      F  , ,  .���  .����  �����  ����  .���      F  , ,  ����  �����  �����  ����  ����      F  , ,  .����  .����  �����  �����  .����      F  , ,  �����  �����  �����  �����  �����      F  , ,  N����  N����  ����  ����  N����      F  , ,  �����  �����  	�����  	�����  �����      F  , ,  
n����  
n����  6����  6����  
n����      F  , ,  �����  �����  �����  �����  �����      F  , ,  �����  �����  V����  V����  �����      F  , ,  ����  ����  �����  �����  ����      F  , ,  �����  �����  v����  v����  �����      F  , ,  >����  >����  ����  ����  >����      F  , ,  ���$  ����  �����  ����$  ���$      F  , ,  ����$  �����  v����  v���$  ����$      F  , ,  >���$  >����  ����  ���$  >���$      F  , ,  N���  N����  ����  ���  N���      F  , ,  ����t  ����<  f���<  f���t  ����t      F  , ,  .���t  .���<  ����<  ����t  .���t      F  , ,  ����t  ����<  ����<  ����t  ����t      F  , ,  N���t  N���<  ���<  ���t  N���t      F  , ,  ����t  ����<  	����<  	����t  ����t      F  , ,  �����  ����|  f���|  f����  �����      F  , ,  .����  .���|  ����|  �����  .����      F  , ,  �����  ����|  ����|  �����  �����      F  , ,  N����  N���|  ���|  ����  N����      F  , ,  �����  ����|  	����|  	�����  �����      F  , ,  
n����  
n���|  6���|  6����  
n����      F  , ,  �����  ����|  ����|  �����  �����      F  , ,  �����  ����|  V���|  V����  �����      F  , ,  �����  ����\  f���\  f����  �����      F  , ,  .����  .���\  ����\  �����  .����      F  , ,  �����  ����\  ����\  �����  �����      F  , ,  N����  N���\  ���\  ����  N����      F  , ,  �����  ����\  	����\  	�����  �����      F  , ,  
n����  
n���\  6���\  6����  
n����      F  , ,  �����  ����\  ����\  �����  �����      F  , ,  �����  ����\  V���\  V����  �����      F  , ,  ����  ���\  ����\  �����  ����      F  , ,  �����  ����\  v���\  v����  �����      F  , ,  >����  >���\  ���\  ����  >����      F  , ,  
n���t  
n���<  6���<  6���t  
n���t      F  , ,  ����t  ����<  ����<  ����t  ����t      F  , ,  ����t  ����<  V���<  V���t  ����t      F  , ,  ���t  ���<  ����<  ����t  ���t      F  , ,  ����t  ����<  v���<  v���t  ����t      F  , ,  ����T  ����  f���  f���T  ����T      F  , ,  .���T  .���  ����  ����T  .���T      F  , ,  ����T  ����  ����  ����T  ����T      F  , ,  N���T  N���  ���  ���T  N���T      F  , ,  ����T  ����  	����  	����T  ����T      F  , ,  
n���T  
n���  6���  6���T  
n���T      F  , ,  ����T  ����  ����  ����T  ����T      F  , ,  ����T  ����  V���  V���T  ����T      F  , ,  ���T  ���  ����  ����T  ���T      F  , ,  ����T  ����  v���  v���T  ����T      F  , ,  >���T  >���  ���  ���T  >���T      F  , ,  >���t  >���<  ���<  ���t  >���t      F  , ,  ����  �����  	�����  	����  ����      F  , ,  
n���  
n����  6����  6���  
n���      F  , ,  ����  �����  �����  ����  ����      F  , ,  ����  �����  V����  V���  ����      F  , ,  ���  ����  �����  ����  ���      F  , ,  ����  �����  v����  v���  ����      F  , ,  >���  >����  ����  ���  >���      F  , ,  ����  �����  f����  f���  ����      F  , ,  .���  .����  �����  ����  .���      F  , ,  �����  �����  	�����  	�����  �����      F  , ,  
n����  
n����  6����  6����  
n����      F  , ,  �����  �����  �����  �����  �����      F  , ,  ����  ���|  ����|  �����  ����      F  , ,  �����  ����|  v���|  v����  �����      F  , ,  >����  >���|  ���|  ����  >����      F  , ,  �����  �����  V����  V����  �����      F  , ,  ����  ����  �����  �����  ����      F  , ,  �����  �����  v����  v����  �����      F  , ,  >����  >����  ����  ����  >����      F  , ,  ����  �����  �����  ����  ����      F  , ,  ����$  �����  f����  f���$  ����$      F  , ,  .���$  .����  �����  ����$  .���$      F  , ,  ����$  �����  �����  ����$  ����$      F  , ,  N���$  N����  ����  ���$  N���$      F  , ,  ����D  ����  	����  	����D  ����D      F  , ,  
n���D  
n���  6���  6���D  
n���D      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  ����D  ����  V���  V���D  ����D      F  , ,  ���D  ���  ����  ����D  ���D      F  , ,  ����D  ����  v���  v���D  ����D      F  , ,  >���D  >���  ���  ���D  >���D      F  , ,  ����$  �����  	�����  	����$  ����$      F  , ,  
n���$  
n����  6����  6���$  
n���$      F  , ,  ����$  �����  �����  ����$  ����$      F  , ,  ����$  �����  V����  V���$  ����$      F  , ,  �����  �����  f����  f����  �����      F  , ,  .����  .����  �����  �����  .����      F  , ,  �����  �����  �����  �����  �����      F  , ,  N����  N����  ����  ����  N����      F  , ,  ����D  ����  f���  f���D  ����D      F  , ,  .���D  .���  ����  ����D  .���D      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  N���D  N���  ���  ���D  N���D      F  , ,  �����  �����  f����  f����  �����      F  , ,  ���  ���L  ����L  ����  ���      F  , ,  ����  ����L  v���L  v���  ����      F  , ,  >���  >���L  ���L  ���  >���      F  , ,  ����  �����  �����  ����  ����      F  , ,  N���  N����  ����  ���  N���      F  , ,  ����  �����  	�����  	����  ����      F  , ,  
n���  
n����  6����  6���  
n���      F  , ,  ����d  ����,  f���,  f���d  ����d      F  , ,  .���d  .���,  ����,  ����d  .���d      F  , ,  ����d  ����,  ����,  ����d  ����d      F  , ,  N���d  N���,  ���,  ���d  N���d      F  , ,  ����d  ����,  	����,  	����d  ����d      F  , ,  
n���d  
n���,  6���,  6���d  
n���d      F  , ,  ����d  ����,  ����,  ����d  ����d      F  , ,  ����d  ����,  V���,  V���d  ����d      F  , ,  ���d  ���,  ����,  ����d  ���d      F  , ,  ����d  ����,  v���,  v���d  ����d      F  , ,  >���d  >���,  ���,  ���d  >���d      F  , ,  ����  �����  �����  ����  ����      F  , ,  ����  �����  V����  V���  ����      F  , ,  ���  ����  �����  ����  ���      F  , ,  ����  �����  v����  v���  ����      F  , ,  >���  >����  ����  ���  >���      F  , ,  ����4  �����  	�����  	����4  ����4      F  , ,  
n���4  
n����  6����  6���4  
n���4      F  , ,  ����4  �����  �����  ����4  ����4      F  , ,  ����4  �����  V����  V���4  ����4      F  , ,  ���4  ����  �����  ����4  ���4      F  , ,  ����4  �����  v����  v���4  ����4      F  , ,  >���4  >����  ����  ���4  >���4      F  , ,  ����4  �����  f����  f���4  ����4      F  , ,  .���4  .����  �����  ����4  .���4      F  , ,  ����  ����l  f���l  f���  ����      F  , ,  .���  .���l  ����l  ����  .���      F  , ,  ����  ����l  ����l  ����  ����      F  , ,  N���  N���l  ���l  ���  N���      F  , ,  ����  ����l  	����l  	����  ����      F  , ,  
n���  
n���l  6���l  6���  
n���      F  , ,  �����  ����  f���  f����  �����      F  , ,  .����  .���  ����  �����  .����      F  , ,  �����  ����  ����  �����  �����      F  , ,  N����  N���  ���  ����  N����      F  , ,  �����  ����  f���  f����  �����      F  , ,  .����  .���  ����  �����  .����      F  , ,  �����  ����  ����  �����  �����      F  , ,  N����  N���  ���  ����  N����      F  , ,  �����  ����  	����  	�����  �����      F  , ,  
n����  
n���  6���  6����  
n����      F  , ,  �����  ����  ����  �����  �����      F  , ,  �����  ����  V���  V����  �����      F  , ,  ����  ���  ����  �����  ����      F  , ,  �����  ����  v���  v����  �����      F  , ,  >����  >���  ���  ����  >����      F  , ,  �����  ����  	����  	�����  �����      F  , ,  
n����  
n���  6���  6����  
n����      F  , ,  �����  ����  ����  �����  �����      F  , ,  �����  ����  V���  V����  �����      F  , ,  ����  ���  ����  �����  ����      F  , ,  �����  ����  v���  v����  �����      F  , ,  >����  >���  ���  ����  >����      F  , ,  ����  ����l  ����l  ����  ����      F  , ,  ����  ����l  V���l  V���  ����      F  , ,  ���  ���l  ����l  ����  ���      F  , ,  ����  ����l  v���l  v���  ����      F  , ,  >���  >���l  ���l  ���  >���      F  , ,  ����4  �����  �����  ����4  ����4      F  , ,  N���4  N����  ����  ���4  N���4      F  , ,  ����  �����  f����  f���  ����      F  , ,  .���  .����  �����  ����  .���      F  , ,  ����  ����L  f���L  f���  ����      F  , ,  .���  .���L  ����L  ����  .���      F  , ,  ����  ����L  ����L  ����  ����      F  , ,  N���  N���L  ���L  ���  N���      F  , ,  ����  ����L  	����L  	����  ����      F  , ,  
n���  
n���L  6���L  6���  
n���      F  , ,  ����  ����L  ����L  ����  ����      F  , ,  ����  ����L  V���L  V���  ����      F  , ,  ����D  ����  f���  f���D  ����D      F  , ,  .���D  .���  ����  ����D  .���D      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  N���D  N���  ���  ���D  N���D      F  , ,  ����D  ����  	����  	����D  ����D      F  , ,  
n���D  
n���  6���  6���D  
n���D      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  ����D  ����  V���  V���D  ����D      F  , ,  ���D  ���  ����  ����D  ���D      F  , ,  ����D  ����  v���  v���D  ����D      F  , ,  >���D  >���  ���  ���D  >���D      F  , ,  ����4  �����  �����  ����4  ����4      F  , ,  ^���4  ^����  &����  &���4  ^���4      F  , ,  ����4  �����  �����  ����4  ����4      F  , ,  ~���4  ~����  F����  F���4  ~���4      F  , ,  ����  ����l  ����l  ����  ����      F  , ,  ^���  ^���l  &���l  &���  ^���      F  , ,  ����  ����l  ����l  ����  ����      F  , ,  ~���  ~���l  F���l  F���  ~���      F  , ,  ���  ���l  ����l  ����  ���      F  , ,  ����  ����l  f���l  f���  ����      F  , ,  ����  �����  �����  ����  ����      F  , ,  ^���  ^����  &����  &���  ^���      F  , ,  ����  �����  �����  ����  ����      F  , ,  ~���  ~����  F����  F���  ~���      F  , ,  ���  ����  �����  ����  ���      F  , ,  ����  �����  f����  f���  ����      F  , ,  .���  .����  �����  ����  .���      F  , ,  ����  �����  �����  ����  ����      F  , ,  $����L  $����  %I���  %I���L  $����L      F  , ,  .���  .���l  ����l  ����  .���      F  , ,  �����  ����  ����  �����  �����      F  , ,  ^����  ^���  &���  &����  ^����      F  , ,  �����  ����  ����  �����  �����      F  , ,  ~����  ~���  F���  F����  ~����      F  , ,  ����  ���  ����  �����  ����      F  , ,  �����  ����  f���  f����  �����      F  , ,  .����  .���  ����  �����  .����      F  , ,  �����  ����  ����  �����  �����      F  , ,  $����  $�����  %I����  %I���  $����      F  , ,  ����  ����l  ����l  ����  ����      F  , ,  $�����  $����  %I���  %I����  $�����      F  , ,  ���4  ����  �����  ����4  ���4      F  , ,  ����4  �����  f����  f���4  ����4      F  , ,  .���4  .����  �����  ����4  .���4      F  , ,  ����4  �����  �����  ����4  ����4      F  , ,  ����  ����L  ����L  ����  ����      F  , ,  ^���  ^���L  &���L  &���  ^���      F  , ,  ����  ����L  ����L  ����  ����      F  , ,  ~���  ~���L  F���L  F���  ~���      F  , ,  ���  ���L  ����L  ����  ���      F  , ,  ����d  ����,  ����,  ����d  ����d      F  , ,  ^���d  ^���,  &���,  &���d  ^���d      F  , ,  ����d  ����,  ����,  ����d  ����d      F  , ,  ~���d  ~���,  F���,  F���d  ~���d      F  , ,  ���d  ���,  ����,  ����d  ���d      F  , ,  ����d  ����,  f���,  f���d  ����d      F  , ,  .���d  .���,  ����,  ����d  .���d      F  , ,  ����d  ����,  ����,  ����d  ����d      F  , ,  $����  $����d  %I���d  %I���  $����      F  , ,  ����  ����L  f���L  f���  ����      F  , ,  .���  .���L  ����L  ����  .���      F  , ,  �����  ����  ����  �����  �����      F  , ,  ^����  ^���  &���  &����  ^����      F  , ,  �����  ����  ����  �����  �����      F  , ,  ~����  ~���  F���  F����  ~����      F  , ,  ����  ���  ����  �����  ����      F  , ,  �����  ����  f���  f����  �����      F  , ,  .����  .���  ����  �����  .����      F  , ,  �����  ����  ����  �����  �����      F  , ,  $����,  $�����  %I����  %I���,  $����,      F  , ,  ����  ����L  ����L  ����  ����      F  , ,  $����  $����  %I���  %I���  $����      F  , ,  $����l  $����4  %I���4  %I���l  $����l      F  , ,  $�����  $�����  %I����  %I����  $�����      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  ^���D  ^���  &���  &���D  ^���D      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  ~���D  ~���  F���  F���D  ~���D      F  , ,  ���D  ���  ����  ����D  ���D      F  , ,  ����D  ����  f���  f���D  ����D      F  , ,  .���D  .���  ����  ����D  .���D      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  $����|  $����D  %I���D  %I���|  $����|      F  , ,  $�����  $����  %I���  %I����  $�����      Y  , ,���������  L   �  L   ����������     �     "�     " "sky130_fd_pr__pfet_01v8_YCMRKB    �   ,���(������(  D  ;�  D  ;�������(���      A   ,����  N����    :/    :/  N����  N      A   ,����������������  :/����  :/������������      A  , ,����  �����  �  <-  �  <-  �����  �      A  , ,�����������  ����}  ����}����������      A  , ,  ;����  ;�  �  <-  �  <-���  ;����      A  , ,�������g�������  <-���  <-���g�������g      ^   ,���T  ����T  �  :�  �  :�  ����T  �      ^   ,���T���}���T���/  :����/  :����}���T���}      ]  , ,���V  r���V    <�    <�  r���V  r      ]  , ,���V������V  r����  r����������V���      ]  , ,  ;���  ;  r  <�  r  <����  ;���      ]  , ,���V�������V���  <����  <��������V����      B   ,   �  �   �  �  �  �  �  �   �  �      B   ,  �  �  �  �    �    �  �  �      B   ,    �    �  h  �  h  �    �      B   ,  l  �  l  �  �  �  �  �  l  �      B   ,  	�  �  	�  �    �    �  	�  �      B   ,    �    �  R  �  R  �    �      B   ,  V  �  V  �  �  �  �  �  V  �      B   ,  �  �  �  �  �  �  �  �  �  �      B   ,  �  �  �  �  <  �  <  �  �  �      B   ,  @  �  @  �  �  �  �  �  @  �      B   ,  �  �  �  �  �  �  �  �  �  �      B   ,  �  �  �  �  &  �  &  �  �  �      B   ,  *  �  *  �  t  �  t  �  *  �      B   ,  x  �  x  �  �  �  �  �  x  �      B   ,   �  �   �  �  "  �  "  �   �  �      B   ,  #  �  #  �  $^  �  $^  �  #  �      B   ,  %b  �  %b  �  &�  �  &�  �  %b  �      B   ,  '�  �  '�  �  (�  �  (�  �  '�  �      B   ,  )�  �  )�  �  +H  �  +H  �  )�  �      B   ,  ,L  �  ,L  �  -�  �  -�  �  ,L  �      B   ,  .�  �  .�  �  /�  �  /�  �  .�  �      B   ,  0�  �  0�  �  22  �  22  �  0�  �      B   ,  36  �  36  �  4�  �  4�  �  36  �      B   ,  5�  �  5�  �  6�  �  6�  �  5�  �      B   ,  7�  �  7�  �  9  �  9  �  7�  �      B   ,   �  �   �  �  �  �  �  �   �  �      B   ,  �  �  �  �    �    �  �  �      B   ,  -  �  -  �  Y  �  Y  �  -  �      B   ,  {  �  {  �  �  �  �  �  {  �      B   ,  	�  �  	�  �  
�  �  
�  �  	�  �      B   ,    �    �  C  �  C  �    �      B   ,  e  �  e  �  �  �  �  �  e  �      B   ,  �  �  �  �  �  �  �  �  �  �      B   ,    �    �  -  �  -  �    �      B   ,  O  �  O  �  {  �  {  �  O  �      B   ,  �  �  �  �  �  �  �  �  �  �      B   ,  �  �  �  �    �    �  �  �      B   ,  9  �  9  �  e  �  e  �  9  �      B   ,  �  �  �  �  �  �  �  �  �  �      B   ,   �  �   �  �  "  �  "  �   �  �      B   ,  ##  �  ##  �  $O  �  $O  �  ##  �      B   ,  %q  �  %q  �  &�  �  &�  �  %q  �      B   ,  '�  �  '�  �  (�  �  (�  �  '�  �      B   ,  *  �  *  �  +9  �  +9  �  *  �      B   ,  ,[  �  ,[  �  -�  �  -�  �  ,[  �      B   ,  .�  �  .�  �  /�  �  /�  �  .�  �      B   ,  0�  �  0�  �  2#  �  2#  �  0�  �      B   ,  3E  �  3E  �  4q  �  4q  �  3E  �      B   ,  5�  �  5�  �  6�  �  6�  �  5�  �      B   ,  7�  �  7�  �  9  �  9  �  7�  �      B   ,   �   i   �  �  �  �  �   i   �   i      B   ,  �   i  �  �    �     i  �   i      B   ,     i    �  h  �  h   i     i      B   ,  l   i  l  �  �  �  �   i  l   i      B   ,  	�   i  	�  �    �     i  	�   i      B   ,     i    �  R  �  R   i     i      B   ,  V   i  V  �  �  �  �   i  V   i      B   ,  �   i  �  �  �  �  �   i  �   i      B   ,  �   i  �  �  <  �  <   i  �   i      B   ,  @   i  @  �  �  �  �   i  @   i      B   ,  �   i  �  �  �  �  �   i  �   i      B   ,  �   i  �  �  &  �  &   i  �   i      B   ,  *   i  *  �  t  �  t   i  *   i      B   ,  x   i  x  �  �  �  �   i  x   i      B   ,   �   i   �  �  "  �  "   i   �   i      B   ,  #   i  #  �  $^  �  $^   i  #   i      B   ,  %b   i  %b  �  &�  �  &�   i  %b   i      B   ,  '�   i  '�  �  (�  �  (�   i  '�   i      B   ,  )�   i  )�  �  +H  �  +H   i  )�   i      B   ,  ,L   i  ,L  �  -�  �  -�   i  ,L   i      B   ,  .�   i  .�  �  /�  �  /�   i  .�   i      B   ,  0�   i  0�  �  22  �  22   i  0�   i      B   ,  36   i  36  �  4�  �  4�   i  36   i      B   ,  5�   i  5�  �  6�  �  6�   i  5�   i      B   ,  7�   i  7�  �  9  �  9   i  7�   i      B   ,����  �����  ����.  ����.  �����  �      B   ,���2  ����2  ����|  ����|  ����2  �      B   ,��ˀ  ���ˀ  �����  �����  ���ˀ  �      B   ,����  �����  ����  ����  �����  �      B   ,���  ����  ����f  ����f  ����  �      B   ,���j  ����j  ���Ӵ  ���Ӵ  ����j  �      B   ,��Ը  ���Ը  ����  ����  ���Ը  �      B   ,���  ����  ����P  ����P  ����  �      B   ,���T  ����T  ���ڞ  ���ڞ  ����T  �      B   ,��ۢ  ���ۢ  �����  �����  ���ۢ  �      B   ,����  �����  ����:  ����:  �����  �      B   ,���>  ����>  ����  ����  ����>  �      B   ,���  ����  �����  �����  ����  �      B   ,����  �����  ����$  ����$  �����  �      B   ,���(  ����(  ����r  ����r  ����(  �      B   ,���v  ����v  �����  �����  ����v  �      B   ,����  �����  ����  ����  �����  �      B   ,���  ����  ����\  ����\  ����  �      B   ,���`  ����`  ����  ����  ����`  �      B   ,���  ����  �����  �����  ����  �      B   ,����  �����  ����F  ����F  �����  �      B   ,���J  ����J  �����  �����  ����J  �      B   ,����  �����  �����  �����  �����  �      B   ,����  �����  ����0  ����0  �����  �      B   ,���4  ����4  ����~  ����~  ����4  �      B   ,����   i����  ����.  ����.   i����   i      B   ,���2   i���2  ����|  ����|   i���2   i      B   ,��ˀ   i��ˀ  �����  �����   i��ˀ   i      B   ,����   i����  ����  ����   i����   i      B   ,���   i���  ����f  ����f   i���   i      B   ,���j   i���j  ���Ӵ  ���Ӵ   i���j   i      B   ,��Ը   i��Ը  ����  ����   i��Ը   i      B   ,���   i���  ����P  ����P   i���   i      B   ,���T   i���T  ���ڞ  ���ڞ   i���T   i      B   ,��ۢ   i��ۢ  �����  �����   i��ۢ   i      B   ,����   i����  ����:  ����:   i����   i      B   ,���>   i���>  ����  ����   i���>   i      B   ,���   i���  �����  �����   i���   i      B   ,����   i����  ����$  ����$   i����   i      B   ,���(   i���(  ����r  ����r   i���(   i      B   ,���v   i���v  �����  �����   i���v   i      B   ,����   i����  ����  ����   i����   i      B   ,���   i���  ����\  ����\   i���   i      B   ,���`   i���`  ����  ����   i���`   i      B   ,���   i���  �����  �����   i���   i      B   ,����   i����  ����F  ����F   i����   i      B   ,���J   i���J  �����  �����   i���J   i      B   ,����   i����  �����  �����   i����   i      B   ,����   i����  ����0  ����0   i����   i      B   ,���4   i���4  ����~  ����~   i���4   i      B   ,����  �����  ����  ����  �����  �      B   ,���A  ����A  ����m  ����m  ����A  �      B   ,��ˏ  ���ˏ  ���̻  ���̻  ���ˏ  �      B   ,����  �����  ����	  ����	  �����  �      B   ,���+  ����+  ����W  ����W  ����+  �      B   ,���y  ����y  ���ӥ  ���ӥ  ����y  �      B   ,����  �����  �����  �����  �����  �      B   ,���  ����  ����A  ����A  ����  �      B   ,���c  ����c  ���ڏ  ���ڏ  ����c  �      B   ,��۱  ���۱  �����  �����  ���۱  �      B   ,����  �����  ����+  ����+  �����  �      B   ,���M  ����M  ����y  ����y  ����M  �      B   ,���  ����  �����  �����  ����  �      B   ,����  �����  ����  ����  �����  �      B   ,���7  ����7  ����c  ����c  ����7  �      B   ,���  ����  ����  ����  ����  �      B   ,����  �����  �����  �����  �����  �      B   ,���!  ����!  ����M  ����M  ����!  �      B   ,���o  ����o  ����  ����  ����o  �      B   ,���  ����  �����  �����  ����  �      B   ,���  ����  ����7  ����7  ����  �      B   ,���Y  ����Y  �����  �����  ����Y  �      B   ,����  �����  �����  �����  �����  �      B   ,����  �����  ����!  ����!  �����  �      B   ,���C  ����C  ����o  ����o  ����C  �      B   ,�������M�����������.�������.���M�������M      B   ,���2���M���2�������|�������|���M���2���M      B   ,��ˀ���M��ˀ�������������������M��ˀ���M      B   ,�������M���������������������M�������M      B   ,������M����������f�������f���M������M      B   ,���j���M���j������Ӵ������Ӵ���M���j���M      B   ,��Ը���M��Ը�����������������M��Ը���M      B   ,������M����������P�������P���M������M      B   ,���T���M���T������ڞ������ڞ���M���T���M      B   ,��ۢ���M��ۢ�������������������M��ۢ���M      B   ,�������M�����������:�������:���M�������M      B   ,���>���M���>�����������������M���>���M      B   ,������M����������������������M������M      B   ,�������M�����������$�������$���M�������M      B   ,���(���M���(�������r�������r���M���(���M      B   ,���v���M���v�������������������M���v���M      B   ,�������M���������������������M�������M      B   ,������M����������\�������\���M������M      B   ,���`���M���`�����������������M���`���M      B   ,������M����������������������M������M      B   ,�������M�����������F�������F���M�������M      B   ,���J���M���J�������������������M���J���M      B   ,�������M�����������������������M�������M      B   ,�������M�����������0�������0���M�������M      B   ,���4���M���4�������~�������~���M���4���M      B   ,�������_�������M������M������_�������_      B   ,���A���_���A���M���m���M���m���_���A���_      B   ,��ˏ���_��ˏ���M��̻���M��̻���_��ˏ���_      B   ,�������_�������M���	���M���	���_�������_      B   ,���+���_���+���M���W���M���W���_���+���_      B   ,���y���_���y���M��ӥ���M��ӥ���_���y���_      B   ,�������_�������M�������M�������_�������_      B   ,������_������M���A���M���A���_������_      B   ,���c���_���c���M��ڏ���M��ڏ���_���c���_      B   ,��۱���_��۱���M�������M�������_��۱���_      B   ,�������_�������M���+���M���+���_�������_      B   ,���M���_���M���M���y���M���y���_���M���_      B   ,������_������M�������M�������_������_      B   ,�������_�������M������M������_�������_      B   ,���7���_���7���M���c���M���c���_���7���_      B   ,������_������M������M������_������_      B   ,�������_�������M�������M�������_�������_      B   ,���!���_���!���M���M���M���M���_���!���_      B   ,���o���_���o���M������M������_���o���_      B   ,������_������M�������M�������_������_      B   ,������_������M���7���M���7���_������_      B   ,���Y���_���Y���M�������M�������_���Y���_      B   ,�������_�������M�������M�������_�������_      B   ,�������_�������M���!���M���!���_�������_      B   ,���C���_���C���M���o���M���o���_���C���_      B   ,��������������_���.���_���.����������      B   ,���2������2���_���|���_���|������2���      B   ,��ˀ�����ˀ���_�������_���������ˀ���      B   ,��������������_������_�������������      B   ,������������_���f���_���f���������      B   ,���j������j���_��Ӵ���_��Ӵ������j���      B   ,��Ը�����Ը���_������_��������Ը���      B   ,������������_���P���_���P���������      B   ,���T������T���_��ڞ���_��ڞ������T���      B   ,��ۢ�����ۢ���_�������_���������ۢ���      B   ,��������������_���:���_���:����������      B   ,���>������>���_������_���������>���      B   ,������������_�������_�������������      B   ,��������������_���$���_���$����������      B   ,���(������(���_���r���_���r������(���      B   ,���v������v���_�������_����������v���      B   ,��������������_������_�������������      B   ,������������_���\���_���\���������      B   ,���`������`���_������_���������`���      B   ,������������_�������_�������������      B   ,��������������_���F���_���F����������      B   ,���J������J���_�������_����������J���      B   ,��������������_�������_��������������      B   ,��������������_���0���_���0����������      B   ,���4������4���_���~���_���~������4���      B   ,   ����_   ����M  ����M  ����_   ����_      B   ,  ����_  ����M  ���M  ���_  ����_      B   ,  -���_  -���M  Y���M  Y���_  -���_      B   ,  {���_  {���M  ����M  ����_  {���_      B   ,  	����_  	����M  
����M  
����_  	����_      B   ,  ���_  ���M  C���M  C���_  ���_      B   ,  e���_  e���M  ����M  ����_  e���_      B   ,  ����_  ����M  ����M  ����_  ����_      B   ,  ���_  ���M  -���M  -���_  ���_      B   ,  O���_  O���M  {���M  {���_  O���_      B   ,  ����_  ����M  ����M  ����_  ����_      B   ,  ����_  ����M  ���M  ���_  ����_      B   ,  9���_  9���M  e���M  e���_  9���_      B   ,  ����_  ����M  ����M  ����_  ����_      B   ,   ����_   ����M  "���M  "���_   ����_      B   ,  ##���_  ##���M  $O���M  $O���_  ##���_      B   ,  %q���_  %q���M  &����M  &����_  %q���_      B   ,  '����_  '����M  (����M  (����_  '����_      B   ,  *���_  *���M  +9���M  +9���_  *���_      B   ,  ,[���_  ,[���M  -����M  -����_  ,[���_      B   ,  .����_  .����M  /����M  /����_  .����_      B   ,  0����_  0����M  2#���M  2#���_  0����_      B   ,  3E���_  3E���M  4q���M  4q���_  3E���_      B   ,  5����_  5����M  6����M  6����_  5����_      B   ,  7����_  7����M  9���M  9���_  7����_      B   ,   ����M   �����  �����  ����M   ����M      B   ,  ����M  �����  ����  ���M  ����M      B   ,  ���M  ����  h����  h���M  ���M      B   ,  l���M  l����  �����  ����M  l���M      B   ,  	����M  	�����  ����  ���M  	����M      B   ,  ���M  ����  R����  R���M  ���M      B   ,  V���M  V����  �����  ����M  V���M      B   ,  ����M  �����  �����  ����M  ����M      B   ,  ����M  �����  <����  <���M  ����M      B   ,  @���M  @����  �����  ����M  @���M      B   ,  ����M  �����  �����  ����M  ����M      B   ,  ����M  �����  &����  &���M  ����M      B   ,  *���M  *����  t����  t���M  *���M      B   ,  x���M  x����  �����  ����M  x���M      B   ,   ����M   �����  "����  "���M   ����M      B   ,  #���M  #����  $^����  $^���M  #���M      B   ,  %b���M  %b����  &�����  &����M  %b���M      B   ,  '����M  '�����  (�����  (����M  '����M      B   ,  )����M  )�����  +H����  +H���M  )����M      B   ,  ,L���M  ,L����  -�����  -����M  ,L���M      B   ,  .����M  .�����  /�����  /����M  .����M      B   ,  0����M  0�����  22����  22���M  0����M      B   ,  36���M  36����  4�����  4����M  36���M      B   ,  5����M  5�����  6�����  6����M  5����M      B   ,  7����M  7�����  9����  9���M  7����M      B   ,   ����   ����_  ����_  ����   ����      B   ,  ����  ����_  ���_  ���  ����      B   ,  ���  ���_  h���_  h���  ���      B   ,  l���  l���_  ����_  ����  l���      B   ,  	����  	����_  ���_  ���  	����      B   ,  ���  ���_  R���_  R���  ���      B   ,  V���  V���_  ����_  ����  V���      B   ,  ����  ����_  ����_  ����  ����      B   ,  ����  ����_  <���_  <���  ����      B   ,  @���  @���_  ����_  ����  @���      B   ,  ����  ����_  ����_  ����  ����      B   ,  ����  ����_  &���_  &���  ����      B   ,  *���  *���_  t���_  t���  *���      B   ,  x���  x���_  ����_  ����  x���      B   ,   ����   ����_  "���_  "���   ����      B   ,  #���  #���_  $^���_  $^���  #���      B   ,  %b���  %b���_  &����_  &����  %b���      B   ,  '����  '����_  (����_  (����  '����      B   ,  )����  )����_  +H���_  +H���  )����      B   ,  ,L���  ,L���_  -����_  -����  ,L���      B   ,  .����  .����_  /����_  /����  .����      B   ,  0����  0����_  22���_  22���  0����      B   ,  36���  36���_  4����_  4����  36���      B   ,  5����  5����_  6����_  6����  5����      B   ,  7����  7����_  9���_  9���  7����      B  , ,����  {����  %   U  %   U  {����  {      B  , ,����  '����  �   U  �   U  '����  '      B  , ,����  	�����  
}   U  
}   U  	�����  	�      B  , ,����  ����  	)   U  	)   U  ����        B  , ,����  +����  �   U  �   U  +����  +      B  , ,����  �����  �   U  �   U  �����  �      B  , ,����  �����  -   U  -   U  �����  �      B  , ,����  /����  �   U  �   U  /����  /      B  , ,�������'��������   U����   U���'�������'      B  , ,���������������}   U���}   U������������      B  , ,��������������)   U���)   U����������      B  , ,�������+��������   U����   U���+�������+      B  , ,����������������   U����   U������������      B  , ,���������������-   U���-   U������������      B  , ,�������/��������   U����   U���/�������/      B  , ,���������������   U���   U������������      B  , ,  �  �  �  �  7  �  7  �  �  �      B  , ,  �  {  �  %  K  %  K  {  �  {      B  , ,  �  '  �  �  K  �  K  '  �  '      B  , ,  �  	�  �  
}  K  
}  K  	�  �  	�      B  , ,  �    �  	)  �  	)  �    �        B  , ,  G    G  	)  �  	)  �    G        B  , ,  �    �  	)  ?  	)  ?    �        B  , ,  �    �  	)  	�  	)  	�    �        B  , ,  1    1  	)  �  	)  �    1        B  , ,        	)  )  	)  )            B  , ,  �    �  	)  w  	)  w    �        B  , ,        	)  �  	)  �            B  , ,  i    i  	)    	)      i        B  , ,  �    �  	)  a  	)  a    �        B  , ,        	)  �  	)  �            B  , ,  S    S  	)  �  	)  �    S        B  , ,  �    �  	)  K  	)  K    �        B  , ,  �    �  	)   �  	)   �    �        B  , ,  "=    "=  	)  "�  	)  "�    "=        B  , ,  $�    $�  	)  %5  	)  %5    $�        B  , ,  &�    &�  	)  '�  	)  '�    &�        B  , ,  )'    )'  	)  )�  	)  )�    )'        B  , ,  +u    +u  	)  ,  	)  ,    +u        B  , ,  -�    -�  	)  .m  	)  .m    -�        B  , ,  0    0  	)  0�  	)  0�    0        B  , ,  2_    2_  	)  3	  	)  3	    2_        B  , ,  4�    4�  	)  5W  	)  5W    4�        B  , ,  6�    6�  	)  7�  	)  7�    6�        B  , ,  9I    9I  	)  9�  	)  9�    9I        B  , ,  ;�  M  ;�  �  <-  �  <-  M  ;�  M      B  , ,  �  +  �  �  K  �  K  +  �  +      B  , ,  �  �  �  �  K  �  K  �  �  �      B  , ,  �  �  �  -  K  -  K  �  �  �      B  , ,  �  /  �  �  K  �  K  /  �  /      B  , ,  4�  {  4�  %  5W  %  5W  {  4�  {      B  , ,  6�  {  6�  %  7�  %  7�  {  6�  {      B  , ,  9I  {  9I  %  9�  %  9�  {  9I  {      B  , ,  ;�  I  ;�  �  <-  �  <-  I  ;�  I      B  , ,   5  �   5  �   �  �   �  �   5  �      B  , ,  �  '  �  �   �  �   �  '  �  '      B  , ,  "=  '  "=  �  "�  �  "�  '  "=  '      B  , ,  $�  '  $�  �  %5  �  %5  '  $�  '      B  , ,  &�  '  &�  �  '�  �  '�  '  &�  '      B  , ,  )'  '  )'  �  )�  �  )�  '  )'  '      B  , ,  +u  '  +u  �  ,  �  ,  '  +u  '      B  , ,  -�  '  -�  �  .m  �  .m  '  -�  '      B  , ,  0  '  0  �  0�  �  0�  '  0  '      B  , ,  2_  '  2_  �  3	  �  3	  '  2_  '      B  , ,  4�  '  4�  �  5W  �  5W  '  4�  '      B  , ,  6�  '  6�  �  7�  �  7�  '  6�  '      B  , ,  9I  '  9I  �  9�  �  9�  '  9I  '      B  , ,  ;�  
�  ;�  �  <-  �  <-  
�  ;�  
�      B  , ,  !�  �  !�  �  "3  �  "3  �  !�  �      B  , ,  �  	�  �  
}   �  
}   �  	�  �  	�      B  , ,  "=  	�  "=  
}  "�  
}  "�  	�  "=  	�      B  , ,  $�  	�  $�  
}  %5  
}  %5  	�  $�  	�      B  , ,  &�  	�  &�  
}  '�  
}  '�  	�  &�  	�      B  , ,  )'  	�  )'  
}  )�  
}  )�  	�  )'  	�      B  , ,  +u  	�  +u  
}  ,  
}  ,  	�  +u  	�      B  , ,  -�  	�  -�  
}  .m  
}  .m  	�  -�  	�      B  , ,  0  	�  0  
}  0�  
}  0�  	�  0  	�      B  , ,  2_  	�  2_  
}  3	  
}  3	  	�  2_  	�      B  , ,  4�  	�  4�  
}  5W  
}  5W  	�  4�  	�      B  , ,  6�  	�  6�  
}  7�  
}  7�  	�  6�  	�      B  , ,  9I  	�  9I  
}  9�  
}  9�  	�  9I  	�      B  , ,  ;�  	�  ;�  
K  <-  
K  <-  	�  ;�  	�      B  , ,  "�  �  "�  �  #�  �  #�  �  "�  �      B  , ,  $1  �  $1  �  $�  �  $�  �  $1  �      B  , ,  %�  �  %�  �  &/  �  &/  �  %�  �      B  , ,  &�  �  &�  �  '�  �  '�  �  &�  �      B  , ,  (-  �  (-  �  (�  �  (�  �  (-  �      B  , ,  )�  �  )�  �  *+  �  *+  �  )�  �      B  , ,  *�  �  *�  �  +  �  +  �  *�  �      B  , ,  ,)  �  ,)  �  ,�  �  ,�  �  ,)  �      B  , ,  -}  �  -}  �  .'  �  .'  �  -}  �      B  , ,  .�  �  .�  �  /{  �  /{  �  .�  �      B  , ,  0%  �  0%  �  0�  �  0�  �  0%  �      B  , ,  1y  �  1y  �  2#  �  2#  �  1y  �      B  , ,  2�  �  2�  �  3w  �  3w  �  2�  �      B  , ,  4!  �  4!  �  4�  �  4�  �  4!  �      B  , ,  5u  �  5u  �  6  �  6  �  5u  �      B  , ,  6�  �  6�  �  7s  �  7s  �  6�  �      B  , ,  8  �  8  �  8�  �  8�  �  8  �      B  , ,  9q  �  9q  �  :  �  :  �  9q  �      B  , ,  ;�  �  ;�  �  <-  �  <-  �  ;�  �      B  , ,  ;�  �  ;�  G  <-  G  <-  �  ;�  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  {  �  %   �  %   �  {  �  {      B  , ,  "=  {  "=  %  "�  %  "�  {  "=  {      B  , ,  $�  {  $�  %  %5  %  %5  {  $�  {      B  , ,  &�  {  &�  %  '�  %  '�  {  &�  {      B  , ,  )'  {  )'  %  )�  %  )�  {  )'  {      B  , ,  +u  {  +u  %  ,  %  ,  {  +u  {      B  , ,  -�  {  -�  %  .m  %  .m  {  -�  {      B  , ,  0  {  0  %  0�  %  0�  {  0  {      B  , ,  2_  {  2_  %  3	  %  3	  {  2_  {      B  , ,  S  	�  S  
}  �  
}  �  	�  S  	�      B  , ,  �  {  �  %  ?  %  ?  {  �  {      B  , ,  �  {  �  %  	�  %  	�  {  �  {      B  , ,  1  {  1  %  �  %  �  {  1  {      B  , ,    {    %  )  %  )  {    {      B  , ,  �  {  �  %  w  %  w  {  �  {      B  , ,  �  �  �  �  S  �  S  �  �  �      B  , ,  �  '  �  �  �  �  �  '  �  '      B  , ,  G  '  G  �  �  �  �  '  G  '      B  , ,  �  '  �  �  ?  �  ?  '  �  '      B  , ,  �  '  �  �  	�  �  	�  '  �  '      B  , ,  1  '  1  �  �  �  �  '  1  '      B  , ,    '    �  )  �  )  '    '      B  , ,  �  '  �  �  w  �  w  '  �  '      B  , ,    '    �  �  �  �  '    '      B  , ,  Q  �  Q  �  �  �  �  �  Q  �      B  , ,  i  '  i  �    �    '  i  '      B  , ,  �  '  �  �  a  �  a  '  �  '      B  , ,    '    �  �  �  �  '    '      B  , ,  S  '  S  �  �  �  �  '  S  '      B  , ,    {    %  �  %  �  {    {      B  , ,  i  {  i  %    %    {  i  {      B  , ,  �  {  �  %  a  %  a  {  �  {      B  , ,    {    %  �  %  �  {    {      B  , ,  S  {  S  %  �  %  �  {  S  {      B  , ,  �  �  �  �  ?  �  ?  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  =  �  =  �  �  �  �  �  =  �      B  , ,  �  �  �  �  ;  �  ;  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  9  �  9  �  �  �  �  �  9  �      B  , ,   U  �   U  �   �  �   �  �   U  �      B  , ,  �  {  �  %  �  %  �  {  �  {      B  , ,  G  {  G  %  �  %  �  {  G  {      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  	�  �  
}  �  
}  �  	�  �  	�      B  , ,  G  	�  G  
}  �  
}  �  	�  G  	�      B  , ,  �  	�  �  
}  ?  
}  ?  	�  �  	�      B  , ,  �  	�  �  
}  	�  
}  	�  	�  �  	�      B  , ,  1  	�  1  
}  �  
}  �  	�  1  	�      B  , ,    	�    
}  )  
}  )  	�    	�      B  , ,  �  	�  �  
}  w  
}  w  	�  �  	�      B  , ,  �  �  �  �  O  �  O  �  �  �      B  , ,    	�    
}  �  
}  �  	�    	�      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  i  	�  i  
}    
}    	�  i  	�      B  , ,  M  �  M  �  �  �  �  �  M  �      B  , ,  �  	�  �  
}  a  
}  a  	�  �  	�      B  , ,  	�  �  	�  �  
K  �  
K  �  	�  �      B  , ,    	�    
}  �  
}  �  	�    	�      B  , ,  
�  �  
�  �  �  �  �  �  
�  �      B  , ,  I  �  I  �  �  �  �  �  I  �      B  , ,  �  �  �  �  G  �  G  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  E  �  E  �  �  �  �  �  E  �      B  , ,  �  �  �  �  C  �  C  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  A  �  A  �  �  �  �  �  A  �      B  , ,  G  �  G  �  �  �  �  �  G  �      B  , ,  �  �  �  �  ?  �  ?  �  �  �      B  , ,  �  �  �  �  	�  �  	�  �  �  �      B  , ,  1  �  1  �  �  �  �  �  1  �      B  , ,    �    �  )  �  )  �    �      B  , ,  �  �  �  �  w  �  w  �  �  �      B  , ,    �    �  �  �  �  �    �      B  , ,  i  �  i  �    �    �  i  �      B  , ,  �  �  �  �  a  �  a  �  �  �      B  , ,    �    �  �  �  �  �    �      B  , ,  S  �  S  �  �  �  �  �  S  �      B  , ,  �  +  �  �  ?  �  ?  +  �  +      B  , ,  �  +  �  �  	�  �  	�  +  �  +      B  , ,  �  �  �  -  �  -  �  �  �  �      B  , ,  G  �  G  -  �  -  �  �  G  �      B  , ,  �  �  �  -  ?  -  ?  �  �  �      B  , ,  �  �  �  -  	�  -  	�  �  �  �      B  , ,  1  �  1  -  �  -  �  �  1  �      B  , ,    �    -  )  -  )  �    �      B  , ,  �  �  �  -  w  -  w  �  �  �      B  , ,    �    -  �  -  �  �    �      B  , ,  i  �  i  -    -    �  i  �      B  , ,  �  �  �  -  a  -  a  �  �  �      B  , ,    �    -  �  -  �  �    �      B  , ,  S  �  S  -  �  -  �  �  S  �      B  , ,  1  +  1  �  �  �  �  +  1  +      B  , ,    +    �  )  �  )  +    +      B  , ,  �  /  �  �  �  �  �  /  �  /      B  , ,  G  /  G  �  �  �  �  /  G  /      B  , ,  �  /  �  �  ?  �  ?  /  �  /      B  , ,  �  /  �  �  	�  �  	�  /  �  /      B  , ,  1  /  1  �  �  �  �  /  1  /      B  , ,    /    �  )  �  )  /    /      B  , ,  �  /  �  �  w  �  w  /  �  /      B  , ,    /    �  �  �  �  /    /      B  , ,  i  /  i  �    �    /  i  /      B  , ,  �  /  �  �  a  �  a  /  �  /      B  , ,    /    �  �  �  �  /    /      B  , ,  S  /  S  �  �  �  �  /  S  /      B  , ,  �  +  �  �  w  �  w  +  �  +      B  , ,   �   �   �  c  |  c  |   �   �   �      B  , ,      �     c  �  c  �   �      �      B  , ,  n   �  n  c    c     �  n   �      B  , ,  �   �  �  c  f  c  f   �  �   �      B  , ,  

   �  

  c  
�  c  
�   �  

   �      B  , ,  X   �  X  c    c     �  X   �      B  , ,  �   �  �  c  P  c  P   �  �   �      B  , ,  �   �  �  c  �  c  �   �  �   �      B  , ,  B   �  B  c  �  c  �   �  B   �      B  , ,  �   �  �  c  :  c  :   �  �   �      B  , ,  �   �  �  c  �  c  �   �  �   �      B  , ,  ,   �  ,  c  �  c  �   �  ,   �      B  , ,  z   �  z  c  $  c  $   �  z   �      B  , ,    +    �  �  �  �  +    +      B  , ,  i  +  i  �    �    +  i  +      B  , ,  �  +  �  �  a  �  a  +  �  +      B  , ,    +    �  �  �  �  +    +      B  , ,  S  +  S  �  �  �  �  +  S  +      B  , ,  �  +  �  �  �  �  �  +  �  +      B  , ,  G  +  G  �  �  �  �  +  G  +      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  4�  �  4�  -  5W  -  5W  �  4�  �      B  , ,  6�  �  6�  -  7�  -  7�  �  6�  �      B  , ,  9I  �  9I  -  9�  -  9�  �  9I  �      B  , ,  ;�  Q  ;�  �  <-  �  <-  Q  ;�  Q      B  , ,  "=  �  "=  �  "�  �  "�  �  "=  �      B  , ,  $�  �  $�  �  %5  �  %5  �  $�  �      B  , ,  &�  �  &�  �  '�  �  '�  �  &�  �      B  , ,  )'  �  )'  �  )�  �  )�  �  )'  �      B  , ,  +u  �  +u  �  ,  �  ,  �  +u  �      B  , ,  -�  �  -�  �  .m  �  .m  �  -�  �      B  , ,  0  �  0  �  0�  �  0�  �  0  �      B  , ,  2_  �  2_  �  3	  �  3	  �  2_  �      B  , ,  4�  �  4�  �  5W  �  5W  �  4�  �      B  , ,  6�  �  6�  �  7�  �  7�  �  6�  �      B  , ,  9I  �  9I  �  9�  �  9�  �  9I  �      B  , ,  ;�  �  ;�  O  <-  O  <-  �  ;�  �      B  , ,  "=  +  "=  �  "�  �  "�  +  "=  +      B  , ,  $�  +  $�  �  %5  �  %5  +  $�  +      B  , ,  �  /  �  �   �  �   �  /  �  /      B  , ,  "=  /  "=  �  "�  �  "�  /  "=  /      B  , ,  $�  /  $�  �  %5  �  %5  /  $�  /      B  , ,  &�  /  &�  �  '�  �  '�  /  &�  /      B  , ,  )'  /  )'  �  )�  �  )�  /  )'  /      B  , ,  +u  /  +u  �  ,  �  ,  /  +u  /      B  , ,  -�  /  -�  �  .m  �  .m  /  -�  /      B  , ,  0  /  0  �  0�  �  0�  /  0  /      B  , ,  2_  /  2_  �  3	  �  3	  /  2_  /      B  , ,  4�  /  4�  �  5W  �  5W  /  4�  /      B  , ,  6�  /  6�  �  7�  �  7�  /  6�  /      B  , ,  9I  /  9I  �  9�  �  9�  /  9I  /      B  , ,  ;�  �  ;�  �  <-  �  <-  �  ;�  �      B  , ,  ;�  �  ;�  S  <-  S  <-  �  ;�  �      B  , ,  &�  +  &�  �  '�  �  '�  +  &�  +      B  , ,  )'  +  )'  �  )�  �  )�  +  )'  +      B  , ,  +u  +  +u  �  ,  �  ,  +  +u  +      B  , ,  -�  +  -�  �  .m  �  .m  +  -�  +      B  , ,  0  +  0  �  0�  �  0�  +  0  +      B  , ,  2_  +  2_  �  3	  �  3	  +  2_  +      B  , ,  4�  +  4�  �  5W  �  5W  +  4�  +      B  , ,  6�  +  6�  �  7�  �  7�  +  6�  +      B  , ,  9I  +  9I  �  9�  �  9�  +  9I  +      B  , ,  ;�  �  ;�  �  <-  �  <-  �  ;�  �      B  , ,  �  +  �  �   �  �   �  +  �  +      B  , ,  �  �  �  �   �  �   �  �  �  �      B  , ,  �  �  �  -   �  -   �  �  �  �      B  , ,  �   �  �  c  r  c  r   �  �   �      B  , ,  !   �  !  c  !�  c  !�   �  !   �      B  , ,  #d   �  #d  c  $  c  $   �  #d   �      B  , ,  %�   �  %�  c  &\  c  &\   �  %�   �      B  , ,  (    �  (   c  (�  c  (�   �  (    �      B  , ,  *N   �  *N  c  *�  c  *�   �  *N   �      B  , ,  ,�   �  ,�  c  -F  c  -F   �  ,�   �      B  , ,  .�   �  .�  c  /�  c  /�   �  .�   �      B  , ,  18   �  18  c  1�  c  1�   �  18   �      B  , ,  3�   �  3�  c  40  c  40   �  3�   �      B  , ,  5�   �  5�  c  6~  c  6~   �  5�   �      B  , ,  8"   �  8"  c  8�  c  8�   �  8"   �      B  , ,  ;�   U  ;�   �  <-   �  <-   U  ;�   U      B  , ,  "=  �  "=  -  "�  -  "�  �  "=  �      B  , ,  $�  �  $�  -  %5  -  %5  �  $�  �      B  , ,  &�  �  &�  -  '�  -  '�  �  &�  �      B  , ,  )'  �  )'  -  )�  -  )�  �  )'  �      B  , ,  +u  �  +u  -  ,  -  ,  �  +u  �      B  , ,  -�  �  -�  -  .m  -  .m  �  -�  �      B  , ,  0  �  0  -  0�  -  0�  �  0  �      B  , ,  2_  �  2_  -  3	  -  3	  �  2_  �      B  , ,���  +���  ����_  ����_  +���  +      B  , ,���  '���  ����_  ����_  '���  '      B  , ,���  ����  ����_  ����_  ����  �      B  , ,���  ����  -���_  -���_  ����  �      B  , ,���  	����  
}���_  
}���_  	����  	�      B  , ,���  {���  %���_  %���_  {���  {      B  , ,���  /���  ����_  ����_  /���  /      B  , ,����  M����  ����}  ����}  M����  M      B  , ,���  ���  	)��Ʒ  	)��Ʒ  ���        B  , ,���[  ���[  	)���  	)���  ���[        B  , ,��ʩ  ��ʩ  	)���S  	)���S  ��ʩ        B  , ,����  ����  	)��͡  	)��͡  ����        B  , ,���E  ���E  	)����  	)����  ���E        B  , ,��ѓ  ��ѓ  	)���=  	)���=  ��ѓ        B  , ,����  ����  	)��ԋ  	)��ԋ  ����        B  , ,���/  ���/  	)����  	)����  ���/        B  , ,���}  ���}  	)���'  	)���'  ���}        B  , ,����  ����  	)���u  	)���u  ����        B  , ,���  ���  	)����  	)����  ���        B  , ,���g  ���g  	)���  	)���  ���g        B  , ,���  ���  	)���_  	)���_  ���        B  , ,���  ���  	)���  	)���  ���        B  , ,���Q  ���Q  	)����  	)����  ���Q        B  , ,���  ���  	)���I  	)���I  ���        B  , ,����  ����  	)���  	)���  ����        B  , ,���;  ���;  	)����  	)����  ���;        B  , ,���  ���  	)���3  	)���3  ���        B  , ,����  ����  	)���  	)���  ����        B  , ,���%  ���%  	)����  	)����  ���%        B  , ,���s  ���s  	)���  	)���  ���s        B  , ,����  ����  	)���k  	)���k  ����        B  , ,���  ���  	)����  	)����  ���        B  , ,���]  ���]  	)���  	)���  ���]        B  , ,����  �����  ����s  ����s  �����  �      B  , ,���  	����  
}���I  
}���I  	����  	�      B  , ,����  	�����  
}���  
}���  	�����  	�      B  , ,���;  	����;  
}����  
}����  	����;  	�      B  , ,���  	����  
}���3  
}���3  	����  	�      B  , ,����  	�����  
}���  
}���  	�����  	�      B  , ,���%  	����%  
}����  
}����  	����%  	�      B  , ,���s  	����s  
}���  
}���  	����s  	�      B  , ,����  	�����  
}���k  
}���k  	�����  	�      B  , ,���  	����  
}����  
}����  	����  	�      B  , ,���]  	����]  
}���  
}���  	����]  	�      B  , ,����  '����  ����  ����  '����  '      B  , ,���  {���  %���  %���  {���  {      B  , ,���Q  {���Q  %����  %����  {���Q  {      B  , ,���  {���  %���I  %���I  {���  {      B  , ,����  {����  %���  %���  {����  {      B  , ,���;  {���;  %����  %����  {���;  {      B  , ,���;  '���;  �����  �����  '���;  '      B  , ,���  {���  %���3  %���3  {���  {      B  , ,����  {����  %���  %���  {����  {      B  , ,���%  {���%  %����  %����  {���%  {      B  , ,���s  {���s  %���  %���  {���s  {      B  , ,����  {����  %���k  %���k  {����  {      B  , ,���  {���  %����  %����  {���  {      B  , ,���]  {���]  %���  %���  {���]  {      B  , ,���  '���  ����3  ����3  '���  '      B  , ,����  '����  ����  ����  '����  '      B  , ,���%  '���%  �����  �����  '���%  '      B  , ,���s  '���s  ����  ����  '���s  '      B  , ,����  '����  ����k  ����k  '����  '      B  , ,���  '���  �����  �����  '���  '      B  , ,���]  '���]  ����  ����  '���]  '      B  , ,���i  ����i  ����  ����  ����i  �      B  , ,���  ����  ����g  ����g  ����  �      B  , ,���  ����  ����  ����  ����  �      B  , ,���e  ����e  ����  ����  ����e  �      B  , ,���  ����  ����c  ����c  ����  �      B  , ,���  ����  ����  ����  ����  �      B  , ,���a  ����a  ����  ����  ����a  �      B  , ,����  �����  ����_  ����_  �����  �      B  , ,���	  ����	  �����  �����  ����	  �      B  , ,���]  ����]  ����  ����  ����]  �      B  , ,���  '���  ����  ����  '���  '      B  , ,����  �����  ����[  ����[  �����  �      B  , ,���  ����  �����  �����  ����  �      B  , ,���Y  ����Y  ����  ����  ����Y  �      B  , ,����  �����  ����W  ����W  �����  �      B  , ,���  ����  �����  �����  ����  �      B  , ,���Q  '���Q  �����  �����  '���Q  '      B  , ,���  '���  ����I  ����I  '���  '      B  , ,���  	����  
}���  
}���  	����  	�      B  , ,���Q  	����Q  
}����  
}����  	����Q  	�      B  , ,���  ����  �����  �����  ����  �      B  , ,���q  ����q  ����  ����  ����q  �      B  , ,����  �����  ����o  ����o  �����  �      B  , ,���  ����  �����  �����  ����  �      B  , ,���m  ����m  ����  ����  ����m  �      B  , ,����  �����  ����k  ����k  �����  �      B  , ,���  ����  ����  ����  ����  �      B  , ,��ѓ  {��ѓ  %���=  %���=  {��ѓ  {      B  , ,����  {����  %��ԋ  %��ԋ  {����  {      B  , ,����  	�����  
K���}  
K���}  	�����  	�      B  , ,���  	����  
}��Ʒ  
}��Ʒ  	����  	�      B  , ,���[  	����[  
}���  
}���  	����[  	�      B  , ,��ʩ  	���ʩ  
}���S  
}���S  	���ʩ  	�      B  , ,����  	�����  
}��͡  
}��͡  	�����  	�      B  , ,��ȍ  ���ȍ  ����7  ����7  ���ȍ  �      B  , ,����  �����  ���ʋ  ���ʋ  �����  �      B  , ,���5  ����5  �����  �����  ����5  �      B  , ,��̉  ���̉  ����3  ����3  ���̉  �      B  , ,����  �����  ���·  ���·  �����  �      B  , ,���1  ����1  �����  �����  ����1  �      B  , ,��Ѕ  ���Ѕ  ����/  ����/  ���Ѕ  �      B  , ,����  �����  ���҃  ���҃  �����  �      B  , ,���-  ����-  �����  �����  ����-  �      B  , ,���E  	����E  
}����  
}����  	����E  	�      B  , ,��ѓ  	���ѓ  
}���=  
}���=  	���ѓ  	�      B  , ,����  	�����  
}��ԋ  
}��ԋ  	�����  	�      B  , ,���/  	����/  
}����  
}����  	����/  	�      B  , ,���}  	����}  
}���'  
}���'  	����}  	�      B  , ,���}  '���}  ����'  ����'  '���}  '      B  , ,����  	�����  
}���u  
}���u  	�����  	�      B  , ,���  	����  
}����  
}����  	����  	�      B  , ,���g  	����g  
}���  
}���  	����g  	�      B  , ,����  '����  ����u  ����u  '����  '      B  , ,���  '���  �����  �����  '���  '      B  , ,���g  '���g  ����  ����  '���g  '      B  , ,��ʩ  '��ʩ  ����S  ����S  '��ʩ  '      B  , ,����  '����  ���͡  ���͡  '����  '      B  , ,���E  '���E  �����  �����  '���E  '      B  , ,��ѓ  '��ѓ  ����=  ����=  '��ѓ  '      B  , ,����  '����  ���ԋ  ���ԋ  '����  '      B  , ,���/  '���/  �����  �����  '���/  '      B  , ,���[  '���[  ����  ����  '���[  '      B  , ,����  �����  ����}  ����}  �����  �      B  , ,����  �����  ���Ə  ���Ə  �����  �      B  , ,����  �����  G���}  G���}  �����  �      B  , ,���/  {���/  %����  %����  {���/  {      B  , ,���}  {���}  %���'  %���'  {���}  {      B  , ,����  {����  %���u  %���u  {����  {      B  , ,���  {���  %����  %����  {���  {      B  , ,��ԁ  ���ԁ  ����+  ����+  ���ԁ  �      B  , ,����  �����  ����  ����  �����  �      B  , ,���)  ����)  �����  �����  ����)  �      B  , ,���}  ����}  ����'  ����'  ����}  �      B  , ,����  �����  ����{  ����{  �����  �      B  , ,���%  ����%  �����  �����  ����%  �      B  , ,���y  ����y  ����#  ����#  ����y  �      B  , ,����  �����  ����w  ����w  �����  �      B  , ,���!  ����!  �����  �����  ����!  �      B  , ,���u  ����u  ����  ����  ����u  �      B  , ,���g  {���g  %���  %���  {���g  {      B  , ,���9  ����9  �����  �����  ����9  �      B  , ,����  I����  ����}  ����}  I����  I      B  , ,���  {���  %��Ʒ  %��Ʒ  {���  {      B  , ,���[  {���[  %���  %���  {���[  {      B  , ,��ʩ  {��ʩ  %���S  %���S  {��ʩ  {      B  , ,����  {����  %��͡  %��͡  {����  {      B  , ,���E  {���E  %����  %����  {���E  {      B  , ,����  
�����  ����}  ����}  
�����  
�      B  , ,���  '���  ���Ʒ  ���Ʒ  '���  '      B  , ,����  +����  ���͡  ���͡  +����  +      B  , ,���E  +���E  �����  �����  +���E  +      B  , ,��ѓ  +��ѓ  ����=  ����=  +��ѓ  +      B  , ,����  +����  ���ԋ  ���ԋ  +����  +      B  , ,���/  +���/  �����  �����  +���/  +      B  , ,���}  +���}  ����'  ����'  +���}  +      B  , ,����  +����  ����u  ����u  +����  +      B  , ,���  +���  �����  �����  +���  +      B  , ,���g  +���g  ����  ����  +���g  +      B  , ,����  �����  ����}  ����}  �����  �      B  , ,���  +���  ���Ʒ  ���Ʒ  +���  +      B  , ,����  �����  O���}  O���}  �����  �      B  , ,���  ����  ���Ʒ  ���Ʒ  ����  �      B  , ,���[  ����[  ����  ����  ����[  �      B  , ,��ʩ  ���ʩ  ����S  ����S  ���ʩ  �      B  , ,����  �����  ���͡  ���͡  �����  �      B  , ,���E  ����E  �����  �����  ����E  �      B  , ,����  �����  S���}  S���}  �����  �      B  , ,��ѓ  ���ѓ  ����=  ����=  ���ѓ  �      B  , ,����   U����   ����}   ����}   U����   U      B  , ,���4   ����4  c����  c����   ����4   �      B  , ,��ɂ   ���ɂ  c���,  c���,   ���ɂ   �      B  , ,����   �����  c���z  c���z   �����   �      B  , ,���   ����  c����  c����   ����   �      B  , ,���l   ����l  c���  c���   ����l   �      B  , ,��Һ   ���Һ  c���d  c���d   ���Һ   �      B  , ,���   ����  c��ղ  c��ղ   ����   �      B  , ,���V   ����V  c���   c���    ����V   �      B  , ,��٤   ���٤  c���N  c���N   ���٤   �      B  , ,����   �����  c��ܜ  c��ܜ   �����   �      B  , ,���@   ����@  c����  c����   ����@   �      B  , ,����   �����  c���8  c���8   �����   �      B  , ,����  �����  ���ԋ  ���ԋ  �����  �      B  , ,���/  ����/  �����  �����  ����/  �      B  , ,���}  ����}  ����'  ����'  ����}  �      B  , ,����  �����  ����u  ����u  �����  �      B  , ,���  ����  �����  �����  ����  �      B  , ,���g  ����g  ����  ����  ����g  �      B  , ,���[  +���[  ����  ����  +���[  +      B  , ,��ʩ  +��ʩ  ����S  ����S  +��ʩ  +      B  , ,����  Q����  ����}  ����}  Q����  Q      B  , ,���  ����  -��Ʒ  -��Ʒ  ����  �      B  , ,����  �����  ����}  ����}  �����  �      B  , ,���  /���  ���Ʒ  ���Ʒ  /���  /      B  , ,���[  /���[  ����  ����  /���[  /      B  , ,��ʩ  /��ʩ  ����S  ����S  /��ʩ  /      B  , ,����  /����  ���͡  ���͡  /����  /      B  , ,���E  /���E  �����  �����  /���E  /      B  , ,��ѓ  /��ѓ  ����=  ����=  /��ѓ  /      B  , ,����  /����  ���ԋ  ���ԋ  /����  /      B  , ,���/  /���/  �����  �����  /���/  /      B  , ,���}  /���}  ����'  ����'  /���}  /      B  , ,����  /����  ����u  ����u  /����  /      B  , ,���  /���  �����  �����  /���  /      B  , ,���g  /���g  ����  ����  /���g  /      B  , ,���[  ����[  -���  -���  ����[  �      B  , ,��ʩ  ���ʩ  -���S  -���S  ���ʩ  �      B  , ,����  �����  -��͡  -��͡  �����  �      B  , ,���E  ����E  -����  -����  ����E  �      B  , ,��ѓ  ���ѓ  -���=  -���=  ���ѓ  �      B  , ,����  �����  -��ԋ  -��ԋ  �����  �      B  , ,���/  ����/  -����  -����  ����/  �      B  , ,���}  ����}  -���'  -���'  ����}  �      B  , ,����  �����  -���u  -���u  �����  �      B  , ,���  ����  -����  -����  ����  �      B  , ,���g  ����g  -���  -���  ����g  �      B  , ,����  �����  -���k  -���k  �����  �      B  , ,���  ����  -����  -����  ����  �      B  , ,���]  ����]  -���  -���  ����]  �      B  , ,���  ����  ����3  ����3  ����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,���%  ����%  �����  �����  ����%  �      B  , ,���s  ����s  ����  ����  ����s  �      B  , ,����  �����  ����k  ����k  �����  �      B  , ,���  /���  ����  ����  /���  /      B  , ,���Q  /���Q  �����  �����  /���Q  /      B  , ,���  /���  ����I  ����I  /���  /      B  , ,����  /����  ����  ����  /����  /      B  , ,���;  /���;  �����  �����  /���;  /      B  , ,���  /���  ����3  ����3  /���  /      B  , ,����   �����  c���  c���   �����   �      B  , ,���*   ����*  c����  c����   ����*   �      B  , ,���x   ����x  c���"  c���"   ����x   �      B  , ,����   �����  c���p  c���p   �����   �      B  , ,���   ����  c���  c���   ����   �      B  , ,���b   ����b  c���  c���   ����b   �      B  , ,���   ����  c���Z  c���Z   ����   �      B  , ,����   �����  c���  c���   �����   �      B  , ,���L   ����L  c����  c����   ����L   �      B  , ,����   �����  c���D  c���D   �����   �      B  , ,����   �����  c����  c����   �����   �      B  , ,���6   ����6  c����  c����   ����6   �      B  , ,����   �����  c���.  c���.   �����   �      B  , ,����  /����  ����  ����  /����  /      B  , ,���%  /���%  �����  �����  /���%  /      B  , ,���s  /���s  ����  ����  /���s  /      B  , ,����  /����  ����k  ����k  /����  /      B  , ,���  /���  �����  �����  /���  /      B  , ,���]  /���]  ����  ����  /���]  /      B  , ,���  ����  �����  �����  ����  �      B  , ,���]  ����]  ����  ����  ����]  �      B  , ,���  +���  ����3  ����3  +���  +      B  , ,����  +����  ����  ����  +����  +      B  , ,���%  +���%  �����  �����  +���%  +      B  , ,���s  +���s  ����  ����  +���s  +      B  , ,����  +����  ����k  ����k  +����  +      B  , ,���  +���  �����  �����  +���  +      B  , ,���]  +���]  ����  ����  +���]  +      B  , ,���  +���  ����  ����  +���  +      B  , ,���Q  +���Q  �����  �����  +���Q  +      B  , ,���  +���  ����I  ����I  +���  +      B  , ,����  +����  ����  ����  +����  +      B  , ,���;  +���;  �����  �����  +���;  +      B  , ,���  ����  ����  ����  ����  �      B  , ,���Q  ����Q  �����  �����  ����Q  �      B  , ,���  ����  ����I  ����I  ����  �      B  , ,����  �����  ����  ����  �����  �      B  , ,���;  ����;  �����  �����  ����;  �      B  , ,���  ����  -���  -���  ����  �      B  , ,���Q  ����Q  -����  -����  ����Q  �      B  , ,���  ����  -���I  -���I  ����  �      B  , ,����  �����  -���  -���  �����  �      B  , ,���;  ����;  -����  -����  ����;  �      B  , ,���  ����  -���3  -���3  ����  �      B  , ,����  �����  -���  -���  �����  �      B  , ,���%  ����%  -����  -����  ����%  �      B  , ,���s  ����s  -���  -���  ����s  �      B  , ,������'����������_�������_���'������'      B  , ,�������������}���_���}���_�����������      B  , ,������������)���_���)���_���������      B  , ,������+����������_�������_���+������+      B  , ,�������	�����������}�������}���	�������	      B  , ,����������������Ʒ������Ʒ�����������      B  , ,���[�������[���������������������[����      B  , ,��ʩ������ʩ�������S�������S������ʩ����      B  , ,������������������͡������͡������������      B  , ,���E�������E�����������������������E����      B  , ,��ѓ������ѓ�������=�������=������ѓ����      B  , ,������������������ԋ������ԋ������������      B  , ,���/�������/�����������������������/����      B  , ,���}�������}�������'�������'�������}����      B  , ,�������������������u�������u������������      B  , ,�������������������������������������      B  , ,���g�������g���������������������g����      B  , ,�����������������_�������_�����������      B  , ,�����������������������������������      B  , ,���Q�������Q�����������������������Q����      B  , ,�����������������I�������I�����������      B  , ,��������������������������������������      B  , ,���;�������;�����������������������;����      B  , ,�����������������3�������3�����������      B  , ,��������������������������������������      B  , ,���%�������%�����������������������%����      B  , ,���s�������s���������������������s����      B  , ,�������������������k�������k������������      B  , ,�������������������������������������      B  , ,���]�������]���������������������]����      B  , ,�������������-���_���-���_�����������      B  , ,������/����������_�������_���/������/      B  , ,����������������_������_�����������      B  , ,�������g����������s������s���g�������g      B  , ,���%�������%���}�������}�����������%����      B  , ,���s�������s���}������}����������s����      B  , ,���������������}���k���}���k������������      B  , ,�������������}�������}���������������      B  , ,���]�������]���}������}����������]����      B  , ,���x�������x���G���"���G���"�������x����      B  , ,������������)������)������������      B  , ,���Q������Q���)�������)����������Q���      B  , ,������������)���I���)���I���������      B  , ,��������������)������)�������������      B  , ,���;������;���)�������)����������;���      B  , ,������������)���3���)���3���������      B  , ,��������������)������)�������������      B  , ,���%������%���)�������)����������%���      B  , ,���s������s���)������)���������s���      B  , ,��������������)���k���)���k����������      B  , ,������������)�������)�������������      B  , ,���]������]���)������)���������]���      B  , ,���������������G���p���G���p������������      B  , ,������+��������������������+������+      B  , ,���Q���+���Q�������������������+���Q���+      B  , ,������+����������I�������I���+������+      B  , ,�������+���������������������+�������+      B  , ,���;���+���;�������������������+���;���+      B  , ,������+����������3�������3���+������+      B  , ,�������+���������������������+�������+      B  , ,���%���+���%�������������������+���%���+      B  , ,���s���+���s�����������������+���s���+      B  , ,�������+�����������k�������k���+�������+      B  , ,������+����������������������+������+      B  , ,���]���+���]�����������������+���]���+      B  , ,�������������G������G��������������      B  , ,���b�������b���G������G����������b����      B  , ,�������������G���Z���G���Z�����������      B  , ,���������������G������G���������������      B  , ,���L�������L���G�������G�����������L����      B  , ,���������������G���D���G���D������������      B  , ,���������������G�������G����������������      B  , ,���6�������6���G�������G�����������6����      B  , ,���������������G���.���G���.������������      B  , ,���������������G������G���������������      B  , ,������'��������������������'������'      B  , ,���Q���'���Q�������������������'���Q���'      B  , ,������'����������I�������I���'������'      B  , ,�������'���������������������'�������'      B  , ,���;���'���;�������������������'���;���'      B  , ,������'����������3�������3���'������'      B  , ,�������'���������������������'�������'      B  , ,���%���'���%�������������������'���%���'      B  , ,���s���'���s�����������������'���s���'      B  , ,�������'�����������k�������k���'�������'      B  , ,������'����������������������'������'      B  , ,���]���'���]�����������������'���]���'      B  , ,���*�������*���G�������G�����������*����      B  , ,�������������}������}��������������      B  , ,���Q�������Q���}�������}�����������Q����      B  , ,�������������}���I���}���I�����������      B  , ,���������������}������}���������������      B  , ,���;�������;���}�������}�����������;����      B  , ,�������������}���3���}���3�����������      B  , ,���������������}������}���������������      B  , ,���[�������[���}������}����������[����      B  , ,��ʩ������ʩ���}���S���}���S������ʩ����      B  , ,���������������}��͡���}��͡������������      B  , ,���E�������E���}�������}�����������E����      B  , ,��ɂ������ɂ���G���,���G���,������ɂ����      B  , ,�������]����������}������}���]�������]      B  , ,������+���������Ʒ������Ʒ���+������+      B  , ,���[���+���[�����������������+���[���+      B  , ,��ʩ���+��ʩ�������S�������S���+��ʩ���+      B  , ,�������+����������͡������͡���+�������+      B  , ,���E���+���E�������������������+���E���+      B  , ,��ѓ���+��ѓ�������=�������=���+��ѓ���+      B  , ,�������+����������ԋ������ԋ���+�������+      B  , ,���/���+���/�������������������+���/���+      B  , ,���}���+���}�������'�������'���+���}���+      B  , ,�������+�����������u�������u���+�������+      B  , ,������+����������������������+������+      B  , ,���g���+���g�����������������+���g���+      B  , ,��ѓ������ѓ���}���=���}���=������ѓ����      B  , ,���������������}��ԋ���}��ԋ������������      B  , ,���/�������/���}�������}�����������/����      B  , ,���}�������}���}���'���}���'�������}����      B  , ,���������������}���u���}���u������������      B  , ,�������������}�������}���������������      B  , ,���g�������g���}������}����������g����      B  , ,�������'����������ԋ������ԋ���'�������'      B  , ,���/���'���/�������������������'���/���'      B  , ,���}���'���}�������'�������'���'���}���'      B  , ,�������'�����������u�������u���'�������'      B  , ,������'����������������������'������'      B  , ,���g���'���g�����������������'���g���'      B  , ,���������������G���z���G���z������������      B  , ,���@�������@���G�������G�����������@����      B  , ,���������������G���8���G���8������������      B  , ,���V�������V���G��� ���G��� �������V����      B  , ,��٤������٤���G���N���G���N������٤����      B  , ,���������������G��ܜ���G��ܜ������������      B  , ,���������������W���}���W���}������������      B  , ,�������Y����������}������}���Y�������Y      B  , ,���4�������4���G�������G�����������4����      B  , ,���������������[���}���[���}������������      B  , ,������������)��Ʒ���)��Ʒ���������      B  , ,���[������[���)������)���������[���      B  , ,��ʩ�����ʩ���)���S���)���S�����ʩ���      B  , ,��������������)��͡���)��͡����������      B  , ,���E������E���)�������)����������E���      B  , ,��ѓ�����ѓ���)���=���)���=�����ѓ���      B  , ,��������������)��ԋ���)��ԋ����������      B  , ,���/������/���)�������)����������/���      B  , ,���}������}���)���'���)���'������}���      B  , ,��������������)���u���)���u����������      B  , ,������������)�������)�������������      B  , ,���g������g���)������)���������g���      B  , ,������'���������Ʒ������Ʒ���'������'      B  , ,���[���'���[�����������������'���[���'      B  , ,��ʩ���'��ʩ�������S�������S���'��ʩ���'      B  , ,�������'����������͡������͡���'�������'      B  , ,���E���'���E�������������������'���E���'      B  , ,�������������G�������G���������������      B  , ,��ѓ���'��ѓ�������=�������=���'��ѓ���'      B  , ,���l�������l���G������G����������l����      B  , ,������������������}�������}����������      B  , ,��Һ������Һ���G���d���G���d������Һ����      B  , ,������������������}�������}����������      B  , ,�������������G��ղ���G��ղ�����������      B  , ,�������������}��Ʒ���}��Ʒ�����������      B  , ,���������������-��ԋ���-��ԋ������������      B  , ,���/�������/���-�������-�����������/����      B  , ,���}�������}���-���'���-���'�������}����      B  , ,���������������-���u���-���u������������      B  , ,�������������-�������-���������������      B  , ,���g�������g���-������-����������g����      B  , ,���������������_���}���_���}������������      B  , ,�������������-��Ʒ���-��Ʒ�����������      B  , ,�������a����������}������}���a�������a      B  , ,������/���������Ʒ������Ʒ���/������/      B  , ,���[���/���[�����������������/���[���/      B  , ,��ʩ���/��ʩ�������S�������S���/��ʩ���/      B  , ,�������/����������͡������͡���/�������/      B  , ,���E���/���E�������������������/���E���/      B  , ,��ѓ���/��ѓ�������=�������=���/��ѓ���/      B  , ,�������/����������ԋ������ԋ���/�������/      B  , ,���/���/���/�������������������/���/���/      B  , ,���}���/���}�������'�������'���/���}���/      B  , ,�������/�����������u�������u���/�������/      B  , ,������/����������������������/������/      B  , ,���g���/���g�����������������/���g���/      B  , ,���[�������[���-������-����������[����      B  , ,��ʩ������ʩ���-���S���-���S������ʩ����      B  , ,�����������������}������}����������      B  , ,���������������Ʒ�����Ʒ�����������      B  , ,���[�������[�������������������[����      B  , ,��ʩ������ʩ������S������S������ʩ����      B  , ,�����������������͡�����͡������������      B  , ,���E�������E���������������������E����      B  , ,��ѓ������ѓ������=������=������ѓ����      B  , ,�����������������ԋ�����ԋ������������      B  , ,���/�������/���������������������/����      B  , ,���}�������}������'������'�������}����      B  , ,������������������u������u������������      B  , ,�����������������������������������      B  , ,���g�������g�������������������g����      B  , ,���������������-��͡���-��͡������������      B  , ,���E�������E���-�������-�����������E����      B  , ,��������������c���}���c���}����������      B  , ,�������e����������}������}���e�������e      B  , ,�������g���������Ə�����Ə���g�������g      B  , ,���9���g���9�����������������g���9���g      B  , ,��ȍ���g��ȍ������7������7���g��ȍ���g      B  , ,�������g���������ʋ�����ʋ���g�������g      B  , ,���5���g���5�����������������g���5���g      B  , ,��̉���g��̉������3������3���g��̉���g      B  , ,�������g���������·�����·���g�������g      B  , ,���1���g���1�����������������g���1���g      B  , ,��Ѕ���g��Ѕ������/������/���g��Ѕ���g      B  , ,�������g���������҃�����҃���g�������g      B  , ,���-���g���-�����������������g���-���g      B  , ,��ԁ���g��ԁ������+������+���g��ԁ���g      B  , ,�������g�������������������g�������g      B  , ,���)���g���)�����������������g���)���g      B  , ,���}���g���}������'������'���g���}���g      B  , ,�������g����������{������{���g�������g      B  , ,���%���g���%�����������������g���%���g      B  , ,���y���g���y������#������#���g���y���g      B  , ,�������g����������w������w���g�������g      B  , ,���!���g���!�����������������g���!���g      B  , ,���u���g���u���������������g���u���g      B  , ,��ѓ������ѓ���-���=���-���=������ѓ����      B  , ,���Q�������Q���������������������Q����      B  , ,����������������I������I�����������      B  , ,������������������������������������      B  , ,���;�������;���������������������;����      B  , ,����������������3������3�����������      B  , ,������������������������������������      B  , ,���%�������%���������������������%����      B  , ,���s�������s�������������������s����      B  , ,������������������k������k������������      B  , ,�����������������������������������      B  , ,���]�������]�������������������]����      B  , ,�������/���������������������/�������/      B  , ,���;���/���;�������������������/���;���/      B  , ,������/����������3�������3���/������/      B  , ,�������/���������������������/�������/      B  , ,���%���/���%�������������������/���%���/      B  , ,���s���/���s�����������������/���s���/      B  , ,�������/�����������k�������k���/�������/      B  , ,������/����������������������/������/      B  , ,���]���/���]�����������������/���]���/      B  , ,���������������-������-���������������      B  , ,���;�������;���-�������-�����������;����      B  , ,�������������-���3���-���3�����������      B  , ,���������������-������-���������������      B  , ,���%�������%���-�������-�����������%����      B  , ,���s�������s���-������-����������s����      B  , ,���������������-���k���-���k������������      B  , ,�������������-�������-���������������      B  , ,���]�������]���-������-����������]����      B  , ,�������������-������-��������������      B  , ,���Q�������Q���-�������-�����������Q����      B  , ,�������������-���I���-���I�����������      B  , ,������/��������������������/������/      B  , ,���Q���/���Q�������������������/���Q���/      B  , ,������/����������I�������I���/������/      B  , ,���������������������������������      B  , ,������g��������������������g������g      B  , ,���q���g���q���������������g���q���g      B  , ,�������g����������o������o���g�������g      B  , ,������g��������������������g������g      B  , ,���m���g���m���������������g���m���g      B  , ,�������g����������k������k���g�������g      B  , ,������g������������������g������g      B  , ,���i���g���i���������������g���i���g      B  , ,������g���������g������g���g������g      B  , ,������g������������������g������g      B  , ,���e���g���e���������������g���e���g      B  , ,������g���������c������c���g������g      B  , ,������g������������������g������g      B  , ,���a���g���a���������������g���a���g      B  , ,�������g����������_������_���g�������g      B  , ,���	���g���	�����������������g���	���g      B  , ,���]���g���]���������������g���]���g      B  , ,�������g����������[������[���g�������g      B  , ,������g��������������������g������g      B  , ,���Y���g���Y���������������g���Y���g      B  , ,�������g����������W������W���g�������g      B  , ,������g��������������������g������g      B  , ,  �����  �����  �����  �����  �����      B  , ,  G����  G����  �����  �����  G����      B  , ,  �����  �����  ?����  ?����  �����      B  , ,  �����  �����  	�����  	�����  �����      B  , ,  1����  1����  �����  �����  1����      B  , ,  ����  ����  )����  )����  ����      B  , ,  �����  �����  w����  w����  �����      B  , ,  ����  ����  �����  �����  ����      B  , ,  i����  i����  ����  ����  i����      B  , ,  �����  �����  a����  a����  �����      B  , ,  ����  ����  �����  �����  ����      B  , ,  S����  S����  �����  �����  S����      B  , ,  �����  �����  K����  K����  �����      B  , ,  �����  �����   �����   �����  �����      B  , ,  "=����  "=����  "�����  "�����  "=����      B  , ,  $�����  $�����  %5����  %5����  $�����      B  , ,  &�����  &�����  '�����  '�����  &�����      B  , ,  )'����  )'����  )�����  )�����  )'����      B  , ,  +u����  +u����  ,����  ,����  +u����      B  , ,  -�����  -�����  .m����  .m����  -�����      B  , ,  0����  0����  0�����  0�����  0����      B  , ,  2_����  2_����  3	����  3	����  2_����      B  , ,  4�����  4�����  5W����  5W����  4�����      B  , ,  6�����  6�����  7�����  7�����  6�����      B  , ,  9I����  9I����  9�����  9�����  9I����      B  , ,  ;����	  ;�����  <-����  <-���	  ;����	      B  , ,  ����'  �����  K����  K���'  ����'      B  , ,  �����  ����-  K���-  K����  �����      B  , ,  ����  ����)  K���)  K���  ����      B  , ,  ����/  �����  K����  K���/  ����/      B  , ,  �����  ����  K���  K����  �����      B  , ,  ����+  �����  K����  K���+  ����+      B  , ,  �����  ����}  K���}  K����  �����      B  , ,  ����g  ����  7���  7���g  ����g      B  , ,  +u���'  +u����  ,����  ,���'  +u���'      B  , ,  -����'  -�����  .m����  .m���'  -����'      B  , ,  0���'  0����  0�����  0����'  0���'      B  , ,  2_���'  2_����  3	����  3	���'  2_���'      B  , ,  4����'  4�����  5W����  5W���'  4����'      B  , ,  6����'  6�����  7�����  7����'  6����'      B  , ,  9I���'  9I����  9�����  9����'  9I���'      B  , ,  ;����Y  ;����  <-���  <-���Y  ;����Y      B  , ,  ;����  ;�����  <-����  <-���  ;����      B  , ,  9I����  9I���}  9����}  9�����  9I����      B  , ,  ����  ����)   ����)   ����  ����      B  , ,  "=���  "=���)  "����)  "����  "=���      B  , ,  $����  $����)  %5���)  %5���  $����      B  , ,  &����  &����)  '����)  '����  &����      B  , ,  )'���  )'���)  )����)  )����  )'���      B  , ,  +u���  +u���)  ,���)  ,���  +u���      B  , ,  -����  -����)  .m���)  .m���  -����      B  , ,  0���  0���)  0����)  0����  0���      B  , ,  2_���  2_���)  3	���)  3	���  2_���      B  , ,  4����  4����)  5W���)  5W���  4����      B  , ,  6����  6����)  7����)  7����  6����      B  , ,  9I���  9I���)  9����)  9����  9I���      B  , ,  ;�����  ;����[  <-���[  <-����  ;�����      B  , ,  ����'  �����   �����   ����'  ����'      B  , ,  �����  ����G  r���G  r����  �����      B  , ,  !����  !���G  !����G  !�����  !����      B  , ,  #d����  #d���G  $���G  $����  #d����      B  , ,  %�����  %����G  &\���G  &\����  %�����      B  , ,  ( ����  ( ���G  (����G  (�����  ( ����      B  , ,  *N����  *N���G  *����G  *�����  *N����      B  , ,  ,�����  ,����G  -F���G  -F����  ,�����      B  , ,  .�����  .����G  /����G  /�����  .�����      B  , ,  18����  18���G  1����G  1�����  18����      B  , ,  3�����  3����G  40���G  40����  3�����      B  , ,  5�����  5����G  6~���G  6~����  5�����      B  , ,  8"����  8"���G  8����G  8�����  8"����      B  , ,  ;����  ;�����  <-����  <-���  ;����      B  , ,  ;�����  ;����W  <-���W  <-����  ;�����      B  , ,  "=���'  "=����  "�����  "����'  "=���'      B  , ,  $����'  $�����  %5����  %5���'  $����'      B  , ,  ����+  �����   �����   ����+  ����+      B  , ,  "=���+  "=����  "�����  "����+  "=���+      B  , ,  $����+  $�����  %5����  %5���+  $����+      B  , ,  &����+  &�����  '�����  '����+  &����+      B  , ,  )'���+  )'����  )�����  )����+  )'���+      B  , ,  +u���+  +u����  ,����  ,���+  +u���+      B  , ,  -����+  -�����  .m����  .m���+  -����+      B  , ,  0���+  0����  0�����  0����+  0���+      B  , ,  2_���+  2_����  3	����  3	���+  2_���+      B  , ,  4����+  4�����  5W����  5W���+  4����+      B  , ,  6����+  6�����  7�����  7����+  6����+      B  , ,  9I���+  9I����  9�����  9����+  9I���+      B  , ,  ;����]  ;����  <-���  <-���]  ;����]      B  , ,  &����'  &�����  '�����  '����'  &����'      B  , ,  �����  ����}   ����}   �����  �����      B  , ,  "=����  "=���}  "����}  "�����  "=����      B  , ,  $�����  $����}  %5���}  %5����  $�����      B  , ,  &�����  &����}  '����}  '�����  &�����      B  , ,  )'����  )'���}  )����}  )�����  )'����      B  , ,  +u����  +u���}  ,���}  ,����  +u����      B  , ,  -�����  -����}  .m���}  .m����  -�����      B  , ,  0����  0���}  0����}  0�����  0����      B  , ,  2_����  2_���}  3	���}  3	����  2_����      B  , ,  4�����  4����}  5W���}  5W����  4�����      B  , ,  6�����  6����}  7����}  7�����  6�����      B  , ,  )'���'  )'����  )�����  )����'  )'���'      B  , ,  i���  i���)  ���)  ���  i���      B  , ,  ����  ����)  a���)  a���  ����      B  , ,  ���  ���)  ����)  ����  ���      B  , ,  S���  S���)  ����)  ����  S���      B  , ,  ����'  �����  	�����  	����'  ����'      B  , ,  1���'  1����  �����  ����'  1���'      B  , ,  ���'  ����  )����  )���'  ���'      B  , ,   �����   ����G  |���G  |����   �����      B  , ,  ����'  �����  w����  w���'  ����'      B  , ,  �����  ����}  ����}  �����  �����      B  , ,  ����+  �����  �����  ����+  ����+      B  , ,  G���+  G����  �����  ����+  G���+      B  , ,  ����+  �����  ?����  ?���+  ����+      B  , ,  ���'  ����  �����  ����'  ���'      B  , ,  ����+  �����  	�����  	����+  ����+      B  , ,  1���+  1����  �����  ����+  1���+      B  , ,  ���+  ����  )����  )���+  ���+      B  , ,  ����+  �����  w����  w���+  ����+      B  , ,  ���+  ����  �����  ����+  ���+      B  , ,  i���+  i����  ����  ���+  i���+      B  , ,  ����+  �����  a����  a���+  ����+      B  , ,  ���+  ����  �����  ����+  ���+      B  , ,  S���+  S����  �����  ����+  S���+      B  , ,  i���'  i����  ����  ���'  i���'      B  , ,  ����'  �����  a����  a���'  ����'      B  , ,  ���'  ����  �����  ����'  ���'      B  , ,  S���'  S����  �����  ����'  S���'      B  , ,  ����'  �����  �����  ����'  ����'      B  , ,  G���'  G����  �����  ����'  G���'      B  , ,   ����   ���G  ����G  �����   ����      B  , ,  ����  ����)  ����)  ����  ����      B  , ,  G���  G���)  ����)  ����  G���      B  , ,  n����  n���G  ���G  ����  n����      B  , ,  �����  ����G  f���G  f����  �����      B  , ,  

����  

���G  
����G  
�����  

����      B  , ,  ����'  �����  ?����  ?���'  ����'      B  , ,  X����  X���G  ���G  ����  X����      B  , ,  G����  G���}  ����}  �����  G����      B  , ,  �����  ����}  ?���}  ?����  �����      B  , ,  �����  ����}  	����}  	�����  �����      B  , ,  1����  1���}  ����}  �����  1����      B  , ,  ����  ���}  )���}  )����  ����      B  , ,  �����  ����}  w���}  w����  �����      B  , ,  ����  ���}  ����}  �����  ����      B  , ,  i����  i���}  ���}  ����  i����      B  , ,  �����  ����}  a���}  a����  �����      B  , ,  ����  ���}  ����}  �����  ����      B  , ,  S����  S���}  ����}  �����  S����      B  , ,  �����  ����G  P���G  P����  �����      B  , ,  �����  ����G  ����G  �����  �����      B  , ,  B����  B���G  ����G  �����  B����      B  , ,  �����  ����G  :���G  :����  �����      B  , ,  �����  ����G  ����G  �����  �����      B  , ,  ,����  ,���G  ����G  �����  ,����      B  , ,  z����  z���G  $���G  $����  z����      B  , ,  ����  ����)  ?���)  ?���  ����      B  , ,  ����  ����)  	����)  	����  ����      B  , ,  1���  1���)  ����)  ����  1���      B  , ,  ���  ���)  )���)  )���  ���      B  , ,  ����  ����)  w���)  w���  ����      B  , ,  ���  ���)  ����)  ����  ���      B  , ,  1���/  1����  �����  ����/  1���/      B  , ,  ���/  ����  )����  )���/  ���/      B  , ,  ����/  �����  w����  w���/  ����/      B  , ,  ���/  ����  �����  ����/  ���/      B  , ,  i���/  i����  ����  ���/  i���/      B  , ,  ����/  �����  a����  a���/  ����/      B  , ,  ���/  ����  �����  ����/  ���/      B  , ,  S���/  S����  �����  ����/  S���/      B  , ,  1����  1���-  ����-  �����  1����      B  , ,  ����  ���-  )���-  )����  ����      B  , ,  �����  ����-  w���-  w����  �����      B  , ,  ����  ���-  ����-  �����  ����      B  , ,  �����  ����  ����  �����  �����      B  , ,  G����  G���  ����  �����  G����      B  , ,  �����  ����  ?���  ?����  �����      B  , ,  �����  ����  	����  	�����  �����      B  , ,  1����  1���  ����  �����  1����      B  , ,  ����  ���  )���  )����  ����      B  , ,  �����  ����  w���  w����  �����      B  , ,  ����  ���  ����  �����  ����      B  , ,  i����  i���  ���  ����  i����      B  , ,  �����  ����  a���  a����  �����      B  , ,  ����  ���  ����  �����  ����      B  , ,  S����  S���  ����  �����  S����      B  , ,  i����  i���-  ���-  ����  i����      B  , ,  �����  ����-  a���-  a����  �����      B  , ,  ����  ���-  ����-  �����  ����      B  , ,  S����  S���-  ����-  �����  S����      B  , ,  �����  ����-  ����-  �����  �����      B  , ,  G����  G���-  ����-  �����  G����      B  , ,  �����  ����-  ?���-  ?����  �����      B  , ,  �����  ����-  	����-  	�����  �����      B  , ,  ����/  �����  �����  ����/  ����/      B  , ,  G���/  G����  �����  ����/  G���/      B  , ,  ����/  �����  ?����  ?���/  ����/      B  , ,   U���g   U���   ����   ����g   U���g      B  , ,  ����g  ����  S���  S���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  Q���g  Q���  ����  ����g  Q���g      B  , ,  ����g  ����  O���  O���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  M���g  M���  ����  ����g  M���g      B  , ,  	����g  	����  
K���  
K���g  	����g      B  , ,  
����g  
����  ����  ����g  
����g      B  , ,  I���g  I���  ����  ����g  I���g      B  , ,  ����g  ����  G���  G���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  E���g  E���  ����  ����g  E���g      B  , ,  ����g  ����  C���  C���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  A���g  A���  ����  ����g  A���g      B  , ,  ����g  ����  ?���  ?���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  =���g  =���  ����  ����g  =���g      B  , ,  ����g  ����  ;���  ;���g  ����g      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,  9���g  9���  ����  ����g  9���g      B  , ,  ����/  �����  	�����  	����/  ����/      B  , ,  $�����  $����  %5���  %5����  $�����      B  , ,  &�����  &����  '����  '�����  &�����      B  , ,  )'����  )'���  )����  )�����  )'����      B  , ,  +u����  +u���  ,���  ,����  +u����      B  , ,  -�����  -����  .m���  .m����  -�����      B  , ,  0����  0���  0����  0�����  0����      B  , ,  2_����  2_���  3	���  3	����  2_����      B  , ,  4�����  4����  5W���  5W����  4�����      B  , ,  6�����  6����  7����  7�����  6�����      B  , ,  9I����  9I���  9����  9�����  9I����      B  , ,  ;����  ;����  <-���  <-���  ;����      B  , ,  "=���/  "=����  "�����  "����/  "=���/      B  , ,  ;����  ;����c  <-���c  <-���  ;����      B  , ,  $����/  $�����  %5����  %5���/  $����/      B  , ,  ;����e  ;����  <-���  <-���e  ;����e      B  , ,  &����/  &�����  '�����  '����/  &����/      B  , ,  )'���/  )'����  )�����  )����/  )'���/      B  , ,  +u���/  +u����  ,����  ,���/  +u���/      B  , ,  -����/  -�����  .m����  .m���/  -����/      B  , ,  0���/  0����  0�����  0����/  0���/      B  , ,  2_���/  2_����  3	����  3	���/  2_���/      B  , ,  4����/  4�����  5W����  5W���/  4����/      B  , ,  6����/  6�����  7�����  7����/  6����/      B  , ,  9I���/  9I����  9�����  9����/  9I���/      B  , ,  ;����a  ;����  <-���  <-���a  ;����a      B  , ,  "=����  "=���-  "����-  "�����  "=����      B  , ,  $�����  $����-  %5���-  %5����  $�����      B  , ,  &�����  &����-  '����-  '�����  &�����      B  , ,  )'����  )'���-  )����-  )�����  )'����      B  , ,  +u����  +u���-  ,���-  ,����  +u����      B  , ,  -�����  -����-  .m���-  .m����  -�����      B  , ,  0����  0���-  0����-  0�����  0����      B  , ,  2_����  2_���-  3	���-  3	����  2_����      B  , ,  4�����  4����-  5W���-  5W����  4�����      B  , ,  6�����  6����-  7����-  7�����  6�����      B  , ,  9I����  9I���-  9����-  9�����  9I����      B  , ,  ;�����  ;����_  <-���_  <-����  ;�����      B  , ,  �����  ����-   ����-   �����  �����      B  , ,  ����/  �����   �����   ����/  ����/      B  , ,  �����  ����   ����   �����  �����      B  , ,  "=����  "=���  "����  "�����  "=����      B  , ,  ����g  ����  ����  ����g  ����g      B  , ,   5���g   5���   ����   ����g   5���g      B  , ,  !����g  !����  "3���  "3���g  !����g      B  , ,  "����g  "����  #����  #����g  "����g      B  , ,  $1���g  $1���  $����  $����g  $1���g      B  , ,  %����g  %����  &/���  &/���g  %����g      B  , ,  &����g  &����  '����  '����g  &����g      B  , ,  (-���g  (-���  (����  (����g  (-���g      B  , ,  )����g  )����  *+���  *+���g  )����g      B  , ,  *����g  *����  +���  +���g  *����g      B  , ,  ,)���g  ,)���  ,����  ,����g  ,)���g      B  , ,  -}���g  -}���  .'���  .'���g  -}���g      B  , ,  .����g  .����  /{���  /{���g  .����g      B  , ,  0%���g  0%���  0����  0����g  0%���g      B  , ,  1y���g  1y���  2#���  2#���g  1y���g      B  , ,  2����g  2����  3w���  3w���g  2����g      B  , ,  4!���g  4!���  4����  4����g  4!���g      B  , ,  5u���g  5u���  6���  6���g  5u���g      B  , ,  6����g  6����  7s���  7s���g  6����g      B  , ,  8���g  8���  8����  8����g  8���g      B  , ,  9q���g  9q���  :���  :���g  9q���g      _   ,�������9����  �  90  �  90���9�������9      C   ,����  �����  �  <-  �  <-  �����  �      C   ,�����������  ����}  ����}����������      C   ,����  :����     U     U  :����  :      C   ,����������������   U����   U������������      C   ,  ;����  ;�  �  <-  �  <-���  ;����      C   ,�������g�������  <-���  <-���g�������g      C   ,  �  :  �    	�    	�  :  �  :      C   ,  1  :  1    �    �  :  1  :      C   ,    :      )    )  :    :      C   ,  �  :  �    w    w  :  �  :      C   ,    :      �    �  :    :      C   ,  i  :  i          :  i  :      C   ,  �  :  �    a    a  :  �  :      C   ,    :      �    �  :    :      C   ,  S  :  S    �    �  :  S  :      C   ,  �  :  �    K    K  :  �  :      C   ,  �  :  �     �     �  :  �  :      C   ,  "=  :  "=    "�    "�  :  "=  :      C   ,  $�  :  $�    %5    %5  :  $�  :      C   ,  &�  :  &�    '�    '�  :  &�  :      C   ,  )'  :  )'    )�    )�  :  )'  :      C   ,  +u  :  +u    ,    ,  :  +u  :      C   ,  -�  :  -�    .m    .m  :  -�  :      C   ,  0  :  0    0�    0�  :  0  :      C   ,  2_  :  2_    3	    3	  :  2_  :      C   ,  4�  :  4�    5W    5W  :  4�  :      C   ,  6�  :  6�    7�    7�  :  6�  :      C   ,  9I  :  9I    9�    9�  :  9I  :      C   ,   �   �   �  c  �  c  �   �   �   �      C   ,  �   �  �  c    c     �  �   �      C   ,     �    c  h  c  h   �     �      C   ,  l   �  l  c  �  c  �   �  l   �      C   ,  	�   �  	�  c    c     �  	�   �      C   ,     �    c  R  c  R   �     �      C   ,  V   �  V  c  �  c  �   �  V   �      C   ,  �   �  �  c  �  c  �   �  �   �      C   ,  �   �  �  c  <  c  <   �  �   �      C   ,  @   �  @  c  �  c  �   �  @   �      C   ,  �   �  �  c  �  c  �   �  �   �      C   ,  �   �  �  c  &  c  &   �  �   �      C   ,  *   �  *  c  t  c  t   �  *   �      C   ,  x   �  x  c  �  c  �   �  x   �      C   ,   �   �   �  c  "  c  "   �   �   �      C   ,  #   �  #  c  $^  c  $^   �  #   �      C   ,  %b   �  %b  c  &�  c  &�   �  %b   �      C   ,  '�   �  '�  c  (�  c  (�   �  '�   �      C   ,  )�   �  )�  c  +H  c  +H   �  )�   �      C   ,  ,L   �  ,L  c  -�  c  -�   �  ,L   �      C   ,  .�   �  .�  c  /�  c  /�   �  .�   �      C   ,  0�   �  0�  c  22  c  22   �  0�   �      C   ,  36   �  36  c  4�  c  4�   �  36   �      C   ,  5�   �  5�  c  6�  c  6�   �  5�   �      C   ,  7�   �  7�  c  9  c  9   �  7�   �      C   ,  �  :  �    �    �  :  �  :      C   ,  G  :  G    �    �  :  G  :      C   ,  �  :  �    ?    ?  :  �  :      C   ,����   �����  c���  c���   �����   �      C   ,���   ����  c���f  c���f   ����   �      C   ,���j   ����j  c��Ӵ  c��Ӵ   ����j   �      C   ,��Ը   ���Ը  c���  c���   ���Ը   �      C   ,���   ����  c���P  c���P   ����   �      C   ,���T   ����T  c��ڞ  c��ڞ   ����T   �      C   ,��ۢ   ���ۢ  c����  c����   ���ۢ   �      C   ,����   �����  c���:  c���:   �����   �      C   ,���>   ����>  c���  c���   ����>   �      C   ,���   ����  c����  c����   ����   �      C   ,����   �����  c���$  c���$   �����   �      C   ,���(   ����(  c���r  c���r   ����(   �      C   ,���v   ����v  c����  c����   ����v   �      C   ,����   �����  c���  c���   �����   �      C   ,���   ����  c���\  c���\   ����   �      C   ,���`   ����`  c���  c���   ����`   �      C   ,���   ����  c����  c����   ����   �      C   ,����   �����  c���F  c���F   �����   �      C   ,���J   ����J  c����  c����   ����J   �      C   ,����   �����  c����  c����   �����   �      C   ,����   �����  c���0  c���0   �����   �      C   ,���4   ����4  c���~  c���~   ����4   �      C   ,���[  :���[  ���  ���  :���[  :      C   ,��ʩ  :��ʩ  ���S  ���S  :��ʩ  :      C   ,����  :����  ��͡  ��͡  :����  :      C   ,���E  :���E  ����  ����  :���E  :      C   ,��ѓ  :��ѓ  ���=  ���=  :��ѓ  :      C   ,����  :����  ��ԋ  ��ԋ  :����  :      C   ,���/  :���/  ����  ����  :���/  :      C   ,���}  :���}  ���'  ���'  :���}  :      C   ,����  :����  ���u  ���u  :����  :      C   ,���  :���  ����  ����  :���  :      C   ,���g  :���g  ���  ���  :���g  :      C   ,���  :���  ���_  ���_  :���  :      C   ,���  :���  ���  ���  :���  :      C   ,���Q  :���Q  ����  ����  :���Q  :      C   ,���  :���  ���I  ���I  :���  :      C   ,����  :����  ���  ���  :����  :      C   ,���;  :���;  ����  ����  :���;  :      C   ,���  :���  ���3  ���3  :���  :      C   ,����  :����  ���  ���  :����  :      C   ,���%  :���%  ����  ����  :���%  :      C   ,���s  :���s  ���  ���  :���s  :      C   ,����  :����  ���k  ���k  :����  :      C   ,���  :���  ����  ����  :���  :      C   ,���]  :���]  ���  ���  :���]  :      C   ,���  :���  ��Ʒ  ��Ʒ  :���  :      C   ,����   �����  c���.  c���.   �����   �      C   ,���2   ����2  c���|  c���|   ����2   �      C   ,��ˀ   ���ˀ  c����  c����   ���ˀ   �      C   ,���������������G������G���������������      C   ,�������������G���f���G���f�����������      C   ,���j�������j���G��Ӵ���G��Ӵ�������j����      C   ,��Ը������Ը���G������G���������Ը����      C   ,�������������G���P���G���P�����������      C   ,���T�������T���G��ڞ���G��ڞ�������T����      C   ,��ۢ������ۢ���G�������G����������ۢ����      C   ,���������������G���:���G���:������������      C   ,���>�������>���G������G����������>����      C   ,�������������G�������G���������������      C   ,���������������G���$���G���$������������      C   ,���(�������(���G���r���G���r�������(����      C   ,���v�������v���G�������G�����������v����      C   ,���������������G������G���������������      C   ,�������������G���\���G���\�����������      C   ,���`�������`���G������G����������`����      C   ,�������������G�������G���������������      C   ,���������������G���F���G���F������������      C   ,���J�������J���G�������G�����������J����      C   ,���������������G�������G����������������      C   ,���������������G���0���G���0������������      C   ,���4�������4���G���~���G���~�������4����      C   ,����������������Ʒ������Ʒ�����������      C   ,���[�������[���������������������[����      C   ,��ʩ������ʩ�������S�������S������ʩ����      C   ,������������������͡������͡������������      C   ,���E�������E�����������������������E����      C   ,��ѓ������ѓ�������=�������=������ѓ����      C   ,������������������ԋ������ԋ������������      C   ,���/�������/�����������������������/����      C   ,���}�������}�������'�������'�������}����      C   ,�������������������u�������u������������      C   ,�������������������������������������      C   ,���g�������g���������������������g����      C   ,�����������������_�������_�����������      C   ,�����������������������������������      C   ,���Q�������Q�����������������������Q����      C   ,�����������������I�������I�����������      C   ,��������������������������������������      C   ,���;�������;�����������������������;����      C   ,�����������������3�������3�����������      C   ,��������������������������������������      C   ,���%�������%�����������������������%����      C   ,���s�������s���������������������s����      C   ,�������������������k�������k������������      C   ,�������������������������������������      C   ,���]�������]���������������������]����      C   ,���������������G���.���G���.������������      C   ,���2�������2���G���|���G���|�������2����      C   ,��ˀ������ˀ���G�������G����������ˀ����      C   ,  l����  l���G  ����G  �����  l����      C   ,  	�����  	����G  ���G  ����  	�����      C   ,  ����  ���G  R���G  R����  ����      C   ,  V����  V���G  ����G  �����  V����      C   ,  �����  ����G  ����G  �����  �����      C   ,  �����  ����G  <���G  <����  �����      C   ,  @����  @���G  ����G  �����  @����      C   ,  �����  ����G  ����G  �����  �����      C   ,  �����  ����G  &���G  &����  �����      C   ,  *����  *���G  t���G  t����  *����      C   ,  x����  x���G  ����G  �����  x����      C   ,   �����   ����G  "���G  "����   �����      C   ,  #����  #���G  $^���G  $^����  #����      C   ,  %b����  %b���G  &����G  &�����  %b����      C   ,  '�����  '����G  (����G  (�����  '�����      C   ,  )�����  )����G  +H���G  +H����  )�����      C   ,  ,L����  ,L���G  -����G  -�����  ,L����      C   ,  .�����  .����G  /����G  /�����  .�����      C   ,  0�����  0����G  22���G  22����  0�����      C   ,  36����  36���G  4����G  4�����  36����      C   ,  5�����  5����G  6����G  6�����  5�����      C   ,  7�����  7����G  9���G  9����  7�����      C   ,   �����   ����G  ����G  �����   �����      C   ,  �����  �����  �����  �����  �����      C   ,  G����  G����  �����  �����  G����      C   ,  �����  �����  ?����  ?����  �����      C   ,  �����  �����  	�����  	�����  �����      C   ,  1����  1����  �����  �����  1����      C   ,  ����  ����  )����  )����  ����      C   ,  �����  �����  w����  w����  �����      C   ,  ����  ����  �����  �����  ����      C   ,  i����  i����  ����  ����  i����      C   ,  �����  �����  a����  a����  �����      C   ,  ����  ����  �����  �����  ����      C   ,  S����  S����  �����  �����  S����      C   ,  �����  �����  K����  K����  �����      C   ,  �����  �����   �����   �����  �����      C   ,  "=����  "=����  "�����  "�����  "=����      C   ,  $�����  $�����  %5����  %5����  $�����      C   ,  &�����  &�����  '�����  '�����  &�����      C   ,  )'����  )'����  )�����  )�����  )'����      C   ,  +u����  +u����  ,����  ,����  +u����      C   ,  -�����  -�����  .m����  .m����  -�����      C   ,  0����  0����  0�����  0�����  0����      C   ,  2_����  2_����  3	����  3	����  2_����      C   ,  4�����  4�����  5W����  5W����  4�����      C   ,  6�����  6�����  7�����  7�����  6�����      C   ,  9I����  9I����  9�����  9�����  9I����      C   ,  �����  ����G  ���G  ����  �����      C   ,  ����  ���G  h���G  h����  ����      C  , ,����  �����  k   U  k   U  �����  �      C  , ,����  Y����     U     U  Y����  Y      C  , ,����  	�����  
�   U  
�   U  	�����  	�      C  , ,����  �����  	3   U  	3   U  �����  �      C  , ,����  !����  �   U  �   U  !����  !      C  , ,����  �����  c   U  c   U  �����  �      C  , ,����  Q����  �   U  �   U  Q����  Q      C  , ,����  �����  �   U  �   U  �����  �      C  , ,�������m�������   U���   U���m�������m      C  , ,���������������   U����   U����������      C  , ,���������������G   U���G   U������������      C  , ,�������5��������   U����   U���5�������5      C  , ,���������������w   U���w   U������������      C  , ,�������e�������   U���   U���e�������e      C  , ,����������������   U����   U������������      C  , ,��������������?   U���?   U����������      C  , ,  z   �  z  c  $  c  $   �  z   �      C  , ,  &�  �  &�  k  '�  k  '�  �  &�  �      C  , ,  )'  �  )'  k  )�  k  )�  �  )'  �      C  , ,  +u  �  +u  k  ,  k  ,  �  +u  �      C  , ,  -�  �  -�  k  .m  k  .m  �  -�  �      C  , ,  0  �  0  k  0�  k  0�  �  0  �      C  , ,  2_  �  2_  k  3	  k  3	  �  2_  �      C  , ,  4�  �  4�  k  5W  k  5W  �  4�  �      C  , ,  6�  �  6�  k  7�  k  7�  �  6�  �      C  , ,  9I  �  9I  k  9�  k  9�  �  9I  �      C  , ,  �  Y  �    K    K  Y  �  Y      C  , ,  �  Y  �     �     �  Y  �  Y      C  , ,  "=  Y  "=    "�    "�  Y  "=  Y      C  , ,  $�  Y  $�    %5    %5  Y  $�  Y      C  , ,  &�  Y  &�    '�    '�  Y  &�  Y      C  , ,  )'  Y  )'    )�    )�  Y  )'  Y      C  , ,  +u  Y  +u    ,    ,  Y  +u  Y      C  , ,  -�  Y  -�    .m    .m  Y  -�  Y      C  , ,  0  Y  0    0�    0�  Y  0  Y      C  , ,  2_  Y  2_    3	    3	  Y  2_  Y      C  , ,  4�  Y  4�    5W    5W  Y  4�  Y      C  , ,  6�  Y  6�    7�    7�  Y  6�  Y      C  , ,  9I  Y  9I    9�    9�  Y  9I  Y      C  , ,  �  	�  �  
�  K  
�  K  	�  �  	�      C  , ,  �  	�  �  
�   �  
�   �  	�  �  	�      C  , ,  "=  	�  "=  
�  "�  
�  "�  	�  "=  	�      C  , ,  $�  	�  $�  
�  %5  
�  %5  	�  $�  	�      C  , ,  &�  	�  &�  
�  '�  
�  '�  	�  &�  	�      C  , ,  )'  	�  )'  
�  )�  
�  )�  	�  )'  	�      C  , ,  +u  	�  +u  
�  ,  
�  ,  	�  +u  	�      C  , ,  -�  	�  -�  
�  .m  
�  .m  	�  -�  	�      C  , ,  0  	�  0  
�  0�  
�  0�  	�  0  	�      C  , ,  2_  	�  2_  
�  3	  
�  3	  	�  2_  	�      C  , ,  4�  	�  4�  
�  5W  
�  5W  	�  4�  	�      C  , ,  6�  	�  6�  
�  7�  
�  7�  	�  6�  	�      C  , ,  9I  	�  9I  
�  9�  
�  9�  	�  9I  	�      C  , ,  �  �  �  	3  K  	3  K  �  �  �      C  , ,  �  �  �  	3   �  	3   �  �  �  �      C  , ,  "=  �  "=  	3  "�  	3  "�  �  "=  �      C  , ,  $�  �  $�  	3  %5  	3  %5  �  $�  �      C  , ,  &�  �  &�  	3  '�  	3  '�  �  &�  �      C  , ,  )'  �  )'  	3  )�  	3  )�  �  )'  �      C  , ,  +u  �  +u  	3  ,  	3  ,  �  +u  �      C  , ,  -�  �  -�  	3  .m  	3  .m  �  -�  �      C  , ,  0  �  0  	3  0�  	3  0�  �  0  �      C  , ,  2_  �  2_  	3  3	  	3  3	  �  2_  �      C  , ,  4�  �  4�  	3  5W  	3  5W  �  4�  �      C  , ,  6�  �  6�  	3  7�  	3  7�  �  6�  �      C  , ,  9I  �  9I  	3  9�  	3  9�  �  9I  �      C  , ,  �  !  �  �  K  �  K  !  �  !      C  , ,  �  !  �  �   �  �   �  !  �  !      C  , ,  "=  !  "=  �  "�  �  "�  !  "=  !      C  , ,  $�  !  $�  �  %5  �  %5  !  $�  !      C  , ,  &�  !  &�  �  '�  �  '�  !  &�  !      C  , ,  )'  !  )'  �  )�  �  )�  !  )'  !      C  , ,  +u  !  +u  �  ,  �  ,  !  +u  !      C  , ,  -�  !  -�  �  .m  �  .m  !  -�  !      C  , ,  0  !  0  �  0�  �  0�  !  0  !      C  , ,  2_  !  2_  �  3	  �  3	  !  2_  !      C  , ,  4�  !  4�  �  5W  �  5W  !  4�  !      C  , ,  6�  !  6�  �  7�  �  7�  !  6�  !      C  , ,  9I  !  9I  �  9�  �  9�  !  9I  !      C  , ,  $�  �  $�  k  %5  k  %5  �  $�  �      C  , ,  �  �  �  k  K  k  K  �  �  �      C  , ,  �  �  �  k   �  k   �  �  �  �      C  , ,  "=  �  "=  k  "�  k  "�  �  "=  �      C  , ,  �  �  �  	3  	�  	3  	�  �  �  �      C  , ,  1  �  1  	3  �  	3  �  �  1  �      C  , ,    �    	3  )  	3  )  �    �      C  , ,  �  �  �  	3  w  	3  w  �  �  �      C  , ,    �    	3  �  	3  �  �    �      C  , ,  i  �  i  	3    	3    �  i  �      C  , ,  �  �  �  	3  a  	3  a  �  �  �      C  , ,    �    	3  �  	3  �  �    �      C  , ,  S  �  S  	3  �  	3  �  �  S  �      C  , ,  G  �  G  k  �  k  �  �  G  �      C  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      C  , ,  G  	�  G  
�  �  
�  �  	�  G  	�      C  , ,  �  	�  �  
�  ?  
�  ?  	�  �  	�      C  , ,  �  	�  �  
�  	�  
�  	�  	�  �  	�      C  , ,  1  	�  1  
�  �  
�  �  	�  1  	�      C  , ,    	�    
�  )  
�  )  	�    	�      C  , ,  �  	�  �  
�  w  
�  w  	�  �  	�      C  , ,    	�    
�  �  
�  �  	�    	�      C  , ,  i  	�  i  
�    
�    	�  i  	�      C  , ,  �  	�  �  
�  a  
�  a  	�  �  	�      C  , ,    	�    
�  �  
�  �  	�    	�      C  , ,  S  	�  S  
�  �  
�  �  	�  S  	�      C  , ,  �  �  �  k  	�  k  	�  �  �  �      C  , ,  �  !  �  �  �  �  �  !  �  !      C  , ,  G  !  G  �  �  �  �  !  G  !      C  , ,  �  !  �  �  ?  �  ?  !  �  !      C  , ,  �  !  �  �  	�  �  	�  !  �  !      C  , ,  1  !  1  �  �  �  �  !  1  !      C  , ,    !    �  )  �  )  !    !      C  , ,  �  !  �  �  w  �  w  !  �  !      C  , ,    !    �  �  �  �  !    !      C  , ,  i  !  i  �    �    !  i  !      C  , ,  �  !  �  �  a  �  a  !  �  !      C  , ,    !    �  �  �  �  !    !      C  , ,  S  !  S  �  �  �  �  !  S  !      C  , ,  �  �  �  k  �  k  �  �  �  �      C  , ,  �  Y  �    �    �  Y  �  Y      C  , ,  G  Y  G    �    �  Y  G  Y      C  , ,  �  Y  �    ?    ?  Y  �  Y      C  , ,  �  Y  �    	�    	�  Y  �  Y      C  , ,  1  Y  1    �    �  Y  1  Y      C  , ,    Y      )    )  Y    Y      C  , ,  �  Y  �    w    w  Y  �  Y      C  , ,    Y      �    �  Y    Y      C  , ,  i  Y  i          Y  i  Y      C  , ,  �  Y  �    a    a  Y  �  Y      C  , ,    Y      �    �  Y    Y      C  , ,  S  Y  S    �    �  Y  S  Y      C  , ,  1  �  1  k  �  k  �  �  1  �      C  , ,    �    k  )  k  )  �    �      C  , ,  �  �  �  k  w  k  w  �  �  �      C  , ,  �  �  �  k  ?  k  ?  �  �  �      C  , ,    �    k  �  k  �  �    �      C  , ,  i  �  i  k    k    �  i  �      C  , ,  �  �  �  k  a  k  a  �  �  �      C  , ,    �    k  �  k  �  �    �      C  , ,  S  �  S  k  �  k  �  �  S  �      C  , ,  �  �  �  	3  �  	3  �  �  �  �      C  , ,  G  �  G  	3  �  	3  �  �  G  �      C  , ,  �  �  �  	3  ?  	3  ?  �  �  �      C  , ,  S  �  S  c  �  c  �  �  S  �      C  , ,  �  �  �  c  �  c  �  �  �  �      C  , ,  �  Q  �  �  �  �  �  Q  �  Q      C  , ,  G  Q  G  �  �  �  �  Q  G  Q      C  , ,  �  Q  �  �  ?  �  ?  Q  �  Q      C  , ,  �  Q  �  �  	�  �  	�  Q  �  Q      C  , ,  1  Q  1  �  �  �  �  Q  1  Q      C  , ,    Q    �  )  �  )  Q    Q      C  , ,  �  Q  �  �  w  �  w  Q  �  Q      C  , ,    Q    �  �  �  �  Q    Q      C  , ,  i  Q  i  �    �    Q  i  Q      C  , ,  �  Q  �  �  a  �  a  Q  �  Q      C  , ,    Q    �  �  �  �  Q    Q      C  , ,  S  Q  S  �  �  �  �  Q  S  Q      C  , ,  G  �  G  c  �  c  �  �  G  �      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,  G  �  G  �  �  �  �  �  G  �      C  , ,  �  �  �  �  ?  �  ?  �  �  �      C  , ,  �  �  �  �  	�  �  	�  �  �  �      C  , ,  1  �  1  �  �  �  �  �  1  �      C  , ,    �    �  )  �  )  �    �      C  , ,  �  �  �  �  w  �  w  �  �  �      C  , ,    �    �  �  �  �  �    �      C  , ,  i  �  i  �    �    �  i  �      C  , ,  �  �  �  �  a  �  a  �  �  �      C  , ,    �    �  �  �  �  �    �      C  , ,  S  �  S  �  �  �  �  �  S  �      C  , ,   �   �   �  c  |  c  |   �   �   �      C  , ,      �     c  �  c  �   �      �      C  , ,  n   �  n  c    c     �  n   �      C  , ,  �   �  �  c  f  c  f   �  �   �      C  , ,  

   �  

  c  
�  c  
�   �  

   �      C  , ,  X   �  X  c    c     �  X   �      C  , ,  �   �  �  c  P  c  P   �  �   �      C  , ,  �   �  �  c  �  c  �   �  �   �      C  , ,  B   �  B  c  �  c  �   �  B   �      C  , ,  �   �  �  c  :  c  :   �  �   �      C  , ,  �   �  �  c  �  c  �   �  �   �      C  , ,  ,   �  ,  c  �  c  �   �  ,   �      C  , ,  �  �  �  c  ?  c  ?  �  �  �      C  , ,  �  �  �  c  	�  c  	�  �  �  �      C  , ,  1  �  1  c  �  c  �  �  1  �      C  , ,    �    c  )  c  )  �    �      C  , ,  �  �  �  c  w  c  w  �  �  �      C  , ,    �    c  �  c  �  �    �      C  , ,  i  �  i  c    c    �  i  �      C  , ,  �  �  �  c  a  c  a  �  �  �      C  , ,    �    c  �  c  �  �    �      C  , ,  0  �  0  c  0�  c  0�  �  0  �      C  , ,  2_  �  2_  c  3	  c  3	  �  2_  �      C  , ,  4�  �  4�  c  5W  c  5W  �  4�  �      C  , ,  6�  �  6�  c  7�  c  7�  �  6�  �      C  , ,  9I  �  9I  c  9�  c  9�  �  9I  �      C  , ,  �  �  �  �  K  �  K  �  �  �      C  , ,  �  �  �  �   �  �   �  �  �  �      C  , ,  "=  �  "=  �  "�  �  "�  �  "=  �      C  , ,  $�  �  $�  �  %5  �  %5  �  $�  �      C  , ,  &�  �  &�  �  '�  �  '�  �  &�  �      C  , ,  )'  �  )'  �  )�  �  )�  �  )'  �      C  , ,  +u  �  +u  �  ,  �  ,  �  +u  �      C  , ,  -�  �  -�  �  .m  �  .m  �  -�  �      C  , ,  0  �  0  �  0�  �  0�  �  0  �      C  , ,  2_  �  2_  �  3	  �  3	  �  2_  �      C  , ,  4�  �  4�  �  5W  �  5W  �  4�  �      C  , ,  6�  �  6�  �  7�  �  7�  �  6�  �      C  , ,  9I  �  9I  �  9�  �  9�  �  9I  �      C  , ,  �  Q  �  �  K  �  K  Q  �  Q      C  , ,  �  Q  �  �   �  �   �  Q  �  Q      C  , ,  "=  Q  "=  �  "�  �  "�  Q  "=  Q      C  , ,  $�  Q  $�  �  %5  �  %5  Q  $�  Q      C  , ,  &�  Q  &�  �  '�  �  '�  Q  &�  Q      C  , ,  )'  Q  )'  �  )�  �  )�  Q  )'  Q      C  , ,  +u  Q  +u  �  ,  �  ,  Q  +u  Q      C  , ,  -�  Q  -�  �  .m  �  .m  Q  -�  Q      C  , ,  0  Q  0  �  0�  �  0�  Q  0  Q      C  , ,  2_  Q  2_  �  3	  �  3	  Q  2_  Q      C  , ,  4�  Q  4�  �  5W  �  5W  Q  4�  Q      C  , ,  6�  Q  6�  �  7�  �  7�  Q  6�  Q      C  , ,  9I  Q  9I  �  9�  �  9�  Q  9I  Q      C  , ,  �   �  �  c  r  c  r   �  �   �      C  , ,  !   �  !  c  !�  c  !�   �  !   �      C  , ,  #d   �  #d  c  $  c  $   �  #d   �      C  , ,  %�   �  %�  c  &\  c  &\   �  %�   �      C  , ,  (    �  (   c  (�  c  (�   �  (    �      C  , ,  *N   �  *N  c  *�  c  *�   �  *N   �      C  , ,  ,�   �  ,�  c  -F  c  -F   �  ,�   �      C  , ,  .�   �  .�  c  /�  c  /�   �  .�   �      C  , ,  18   �  18  c  1�  c  1�   �  18   �      C  , ,  3�   �  3�  c  40  c  40   �  3�   �      C  , ,  5�   �  5�  c  6~  c  6~   �  5�   �      C  , ,  8"   �  8"  c  8�  c  8�   �  8"   �      C  , ,  �  �  �  c  K  c  K  �  �  �      C  , ,  �  �  �  c   �  c   �  �  �  �      C  , ,  "=  �  "=  c  "�  c  "�  �  "=  �      C  , ,  $�  �  $�  c  %5  c  %5  �  $�  �      C  , ,  &�  �  &�  c  '�  c  '�  �  &�  �      C  , ,  )'  �  )'  c  )�  c  )�  �  )'  �      C  , ,  +u  �  +u  c  ,  c  ,  �  +u  �      C  , ,  -�  �  -�  c  .m  c  .m  �  -�  �      C  , ,����   �����  c���  c���   �����   �      C  , ,���  	����  
����I  
����I  	����  	�      C  , ,����  	�����  
����  
����  	�����  	�      C  , ,���;  	����;  
�����  
�����  	����;  	�      C  , ,���  	����  
����3  
����3  	����  	�      C  , ,����  	�����  
����  
����  	�����  	�      C  , ,���%  	����%  
�����  
�����  	����%  	�      C  , ,���s  	����s  
����  
����  	����s  	�      C  , ,����  	�����  
����k  
����k  	�����  	�      C  , ,���  	����  
�����  
�����  	����  	�      C  , ,���]  	����]  
����  
����  	����]  	�      C  , ,���  Y���  ���  ���  Y���  Y      C  , ,���Q  Y���Q  ����  ����  Y���Q  Y      C  , ,���  Y���  ���I  ���I  Y���  Y      C  , ,����  Y����  ���  ���  Y����  Y      C  , ,���;  Y���;  ����  ����  Y���;  Y      C  , ,���  Y���  ���3  ���3  Y���  Y      C  , ,����  Y����  ���  ���  Y����  Y      C  , ,���%  Y���%  ����  ����  Y���%  Y      C  , ,���s  Y���s  ���  ���  Y���s  Y      C  , ,����  Y����  ���k  ���k  Y����  Y      C  , ,���  Y���  ����  ����  Y���  Y      C  , ,���]  Y���]  ���  ���  Y���]  Y      C  , ,���  ����  	3���  	3���  ����  �      C  , ,���Q  ����Q  	3����  	3����  ����Q  �      C  , ,���  ����  	3���I  	3���I  ����  �      C  , ,����  �����  	3���  	3���  �����  �      C  , ,���;  ����;  	3����  	3����  ����;  �      C  , ,���  ����  	3���3  	3���3  ����  �      C  , ,����  �����  	3���  	3���  �����  �      C  , ,���%  ����%  	3����  	3����  ����%  �      C  , ,���s  ����s  	3���  	3���  ����s  �      C  , ,����  �����  	3���k  	3���k  �����  �      C  , ,���  ����  	3����  	3����  ����  �      C  , ,���]  ����]  	3���  	3���  ����]  �      C  , ,���  ����  k���  k���  ����  �      C  , ,���Q  ����Q  k����  k����  ����Q  �      C  , ,���  ����  k���I  k���I  ����  �      C  , ,����  �����  k���  k���  �����  �      C  , ,���;  ����;  k����  k����  ����;  �      C  , ,���  ����  k���3  k���3  ����  �      C  , ,����  �����  k���  k���  �����  �      C  , ,���%  ����%  k����  k����  ����%  �      C  , ,���s  ����s  k���  k���  ����s  �      C  , ,����  �����  k���k  k���k  �����  �      C  , ,���  ����  k����  k����  ����  �      C  , ,���]  ����]  k���  k���  ����]  �      C  , ,���Q  	����Q  
�����  
�����  	����Q  	�      C  , ,���  !���  ����  ����  !���  !      C  , ,���Q  !���Q  �����  �����  !���Q  !      C  , ,���  !���  ����I  ����I  !���  !      C  , ,����  !����  ����  ����  !����  !      C  , ,���;  !���;  �����  �����  !���;  !      C  , ,���  !���  ����3  ����3  !���  !      C  , ,����  !����  ����  ����  !����  !      C  , ,���%  !���%  �����  �����  !���%  !      C  , ,���s  !���s  ����  ����  !���s  !      C  , ,����  !����  ����k  ����k  !����  !      C  , ,���  !���  �����  �����  !���  !      C  , ,���]  !���]  ����  ����  !���]  !      C  , ,���  	����  
����  
����  	����  	�      C  , ,���  Y���  ���_  ���_  Y���  Y      C  , ,����  �����  k��͡  k��͡  �����  �      C  , ,���E  ����E  k����  k����  ����E  �      C  , ,��ѓ  ���ѓ  k���=  k���=  ���ѓ  �      C  , ,����  �����  k��ԋ  k��ԋ  �����  �      C  , ,���/  ����/  k����  k����  ����/  �      C  , ,���}  ����}  k���'  k���'  ����}  �      C  , ,����  �����  k���u  k���u  �����  �      C  , ,���  ����  k����  k����  ����  �      C  , ,���g  ����g  k���  k���  ����g  �      C  , ,���  ����  k���_  k���_  ����  �      C  , ,���[  ����[  k���  k���  ����[  �      C  , ,��ʩ  ���ʩ  k���S  k���S  ���ʩ  �      C  , ,���  ����  	3��Ʒ  	3��Ʒ  ����  �      C  , ,���[  ����[  	3���  	3���  ����[  �      C  , ,��ʩ  ���ʩ  	3���S  	3���S  ���ʩ  �      C  , ,����  �����  	3��͡  	3��͡  �����  �      C  , ,���E  ����E  	3����  	3����  ����E  �      C  , ,��ѓ  ���ѓ  	3���=  	3���=  ���ѓ  �      C  , ,����  �����  	3��ԋ  	3��ԋ  �����  �      C  , ,���/  ����/  	3����  	3����  ����/  �      C  , ,���}  ����}  	3���'  	3���'  ����}  �      C  , ,����  �����  	3���u  	3���u  �����  �      C  , ,���  ����  k��Ʒ  k��Ʒ  ����  �      C  , ,���  Y���  ��Ʒ  ��Ʒ  Y���  Y      C  , ,���  	����  
���Ʒ  
���Ʒ  	����  	�      C  , ,���[  	����[  
����  
����  	����[  	�      C  , ,���  !���  ���Ʒ  ���Ʒ  !���  !      C  , ,���[  !���[  ����  ����  !���[  !      C  , ,��ʩ  !��ʩ  ����S  ����S  !��ʩ  !      C  , ,����  !����  ���͡  ���͡  !����  !      C  , ,���  ����  	3����  	3����  ����  �      C  , ,���E  !���E  �����  �����  !���E  !      C  , ,��ѓ  !��ѓ  ����=  ����=  !��ѓ  !      C  , ,����  !����  ���ԋ  ���ԋ  !����  !      C  , ,���/  !���/  �����  �����  !���/  !      C  , ,���}  !���}  ����'  ����'  !���}  !      C  , ,����  !����  ����u  ����u  !����  !      C  , ,���  !���  �����  �����  !���  !      C  , ,���g  !���g  ����  ����  !���g  !      C  , ,���  !���  ����_  ����_  !���  !      C  , ,���g  ����g  	3���  	3���  ����g  �      C  , ,���  ����  	3���_  	3���_  ����  �      C  , ,���[  Y���[  ���  ���  Y���[  Y      C  , ,��ʩ  Y��ʩ  ���S  ���S  Y��ʩ  Y      C  , ,����  Y����  ��͡  ��͡  Y����  Y      C  , ,���E  Y���E  ����  ����  Y���E  Y      C  , ,��ѓ  Y��ѓ  ���=  ���=  Y��ѓ  Y      C  , ,����  Y����  ��ԋ  ��ԋ  Y����  Y      C  , ,���/  Y���/  ����  ����  Y���/  Y      C  , ,���}  Y���}  ���'  ���'  Y���}  Y      C  , ,����  Y����  ���u  ���u  Y����  Y      C  , ,���  Y���  ����  ����  Y���  Y      C  , ,��ʩ  	���ʩ  
����S  
����S  	���ʩ  	�      C  , ,����  	�����  
���͡  
���͡  	�����  	�      C  , ,���E  	����E  
�����  
�����  	����E  	�      C  , ,��ѓ  	���ѓ  
����=  
����=  	���ѓ  	�      C  , ,����  	�����  
���ԋ  
���ԋ  	�����  	�      C  , ,���/  	����/  
�����  
�����  	����/  	�      C  , ,���}  	����}  
����'  
����'  	����}  	�      C  , ,����  	�����  
����u  
����u  	�����  	�      C  , ,���  	����  
�����  
�����  	����  	�      C  , ,���g  	����g  
����  
����  	����g  	�      C  , ,���  	����  
����_  
����_  	����  	�      C  , ,���g  Y���g  ���  ���  Y���g  Y      C  , ,���}  Q���}  ����'  ����'  Q���}  Q      C  , ,����  Q����  ����u  ����u  Q����  Q      C  , ,���  Q���  �����  �����  Q���  Q      C  , ,���g  Q���g  ����  ����  Q���g  Q      C  , ,���  Q���  ����_  ����_  Q���  Q      C  , ,���4   ����4  c����  c����   ����4   �      C  , ,��ɂ   ���ɂ  c���,  c���,   ���ɂ   �      C  , ,����   �����  c���z  c���z   �����   �      C  , ,���   ����  c����  c����   ����   �      C  , ,���l   ����l  c���  c���   ����l   �      C  , ,��Һ   ���Һ  c���d  c���d   ���Һ   �      C  , ,���   ����  c��ղ  c��ղ   ����   �      C  , ,���V   ����V  c���   c���    ����V   �      C  , ,��٤   ���٤  c���N  c���N   ���٤   �      C  , ,����   �����  c��ܜ  c��ܜ   �����   �      C  , ,���@   ����@  c����  c����   ����@   �      C  , ,����   �����  c���8  c���8   �����   �      C  , ,���  ����  ���Ʒ  ���Ʒ  ����  �      C  , ,���[  ����[  ����  ����  ����[  �      C  , ,��ʩ  ���ʩ  ����S  ����S  ���ʩ  �      C  , ,����  �����  ���͡  ���͡  �����  �      C  , ,���E  ����E  �����  �����  ����E  �      C  , ,��ѓ  ���ѓ  ����=  ����=  ���ѓ  �      C  , ,����  �����  ���ԋ  ���ԋ  �����  �      C  , ,���/  ����/  �����  �����  ����/  �      C  , ,���}  ����}  ����'  ����'  ����}  �      C  , ,����  �����  ����u  ����u  �����  �      C  , ,���  ����  �����  �����  ����  �      C  , ,���g  ����g  ����  ����  ����g  �      C  , ,���  ����  ����_  ����_  ����  �      C  , ,���  ����  c��Ʒ  c��Ʒ  ����  �      C  , ,���[  ����[  c���  c���  ����[  �      C  , ,��ʩ  ���ʩ  c���S  c���S  ���ʩ  �      C  , ,����  �����  c��͡  c��͡  �����  �      C  , ,���E  ����E  c����  c����  ����E  �      C  , ,��ѓ  ���ѓ  c���=  c���=  ���ѓ  �      C  , ,����  �����  c��ԋ  c��ԋ  �����  �      C  , ,���/  ����/  c����  c����  ����/  �      C  , ,���}  ����}  c���'  c���'  ����}  �      C  , ,����  �����  c���u  c���u  �����  �      C  , ,���  ����  c����  c����  ����  �      C  , ,���g  ����g  c���  c���  ����g  �      C  , ,���  ����  c���_  c���_  ����  �      C  , ,���  Q���  ���Ʒ  ���Ʒ  Q���  Q      C  , ,���[  Q���[  ����  ����  Q���[  Q      C  , ,��ʩ  Q��ʩ  ����S  ����S  Q��ʩ  Q      C  , ,����  Q����  ���͡  ���͡  Q����  Q      C  , ,���E  Q���E  �����  �����  Q���E  Q      C  , ,��ѓ  Q��ѓ  ����=  ����=  Q��ѓ  Q      C  , ,����  Q����  ���ԋ  ���ԋ  Q����  Q      C  , ,���/  Q���/  �����  �����  Q���/  Q      C  , ,����  Q����  ����  ����  Q����  Q      C  , ,���;  Q���;  �����  �����  Q���;  Q      C  , ,���  Q���  ����3  ����3  Q���  Q      C  , ,���*   ����*  c����  c����   ����*   �      C  , ,���x   ����x  c���"  c���"   ����x   �      C  , ,����   �����  c���p  c���p   �����   �      C  , ,���   ����  c���  c���   ����   �      C  , ,���b   ����b  c���  c���   ����b   �      C  , ,���   ����  c���Z  c���Z   ����   �      C  , ,����   �����  c���  c���   �����   �      C  , ,���L   ����L  c����  c����   ����L   �      C  , ,����   �����  c���D  c���D   �����   �      C  , ,����   �����  c����  c����   �����   �      C  , ,���6   ����6  c����  c����   ����6   �      C  , ,����   �����  c���.  c���.   �����   �      C  , ,����  Q����  ����  ����  Q����  Q      C  , ,���%  Q���%  �����  �����  Q���%  Q      C  , ,���s  Q���s  ����  ����  Q���s  Q      C  , ,����  Q����  ����k  ����k  Q����  Q      C  , ,���  Q���  �����  �����  Q���  Q      C  , ,���]  Q���]  ����  ����  Q���]  Q      C  , ,����  �����  c���  c���  �����  �      C  , ,���;  ����;  c����  c����  ����;  �      C  , ,���  ����  c���3  c���3  ����  �      C  , ,����  �����  c���  c���  �����  �      C  , ,���%  ����%  c����  c����  ����%  �      C  , ,���s  ����s  c���  c���  ����s  �      C  , ,����  �����  c���k  c���k  �����  �      C  , ,���  ����  c����  c����  ����  �      C  , ,���]  ����]  c���  c���  ����]  �      C  , ,���  ����  c���  c���  ����  �      C  , ,���Q  ����Q  c����  c����  ����Q  �      C  , ,���  ����  c���I  c���I  ����  �      C  , ,���  Q���  ����  ����  Q���  Q      C  , ,���Q  Q���Q  �����  �����  Q���Q  Q      C  , ,���  Q���  ����I  ����I  Q���  Q      C  , ,���  ����  ����  ����  ����  �      C  , ,���Q  ����Q  �����  �����  ����Q  �      C  , ,���  ����  ����I  ����I  ����  �      C  , ,����  �����  ����  ����  �����  �      C  , ,���;  ����;  �����  �����  ����;  �      C  , ,���  ����  ����3  ����3  ����  �      C  , ,����  �����  ����  ����  �����  �      C  , ,���%  ����%  �����  �����  ����%  �      C  , ,���s  ����s  ����  ����  ����s  �      C  , ,����  �����  ����k  ����k  �����  �      C  , ,���  ����  �����  �����  ����  �      C  , ,���]  ����]  ����  ����  ����]  �      C  , ,���������������G������G���������������      C  , ,���*�������*���G�������G�����������*����      C  , ,���x�������x���G���"���G���"�������x����      C  , ,���������������G���p���G���p������������      C  , ,�������������G������G��������������      C  , ,���b�������b���G������G����������b����      C  , ,�������������G���Z���G���Z�����������      C  , ,���������������G������G���������������      C  , ,���L�������L���G�������G�����������L����      C  , ,���������������G���D���G���D������������      C  , ,���������������G�������G����������������      C  , ,���6�������6���G�������G�����������6����      C  , ,���������������G���.���G���.������������      C  , ,������m������������������m������m      C  , ,���Q���m���Q�����������������m���Q���m      C  , ,������m���������I������I���m������m      C  , ,�������m�������������������m�������m      C  , ,���;���m���;�����������������m���;���m      C  , ,������m���������3������3���m������m      C  , ,�������m�������������������m�������m      C  , ,���%���m���%�����������������m���%���m      C  , ,���s���m���s���������������m���s���m      C  , ,�������m����������k������k���m�������m      C  , ,������m��������������������m������m      C  , ,���]���m���]���������������m���]���m      C  , ,��������������������������������      C  , ,���Q������Q����������������������Q���      C  , ,����������������I�������I���������      C  , ,�����������������������������������      C  , ,���;������;����������������������;���      C  , ,����������������3�������3���������      C  , ,�����������������������������������      C  , ,���%������%����������������������%���      C  , ,���s������s��������������������s���      C  , ,������������������k�������k����������      C  , ,����������������������������������      C  , ,���]������]��������������������]���      C  , ,�������������G������G��������������      C  , ,���Q�������Q���G�������G�����������Q����      C  , ,�������������G���I���G���I�����������      C  , ,���������������G������G���������������      C  , ,���;�������;���G�������G�����������;����      C  , ,�������������G���3���G���3�����������      C  , ,���������������G������G���������������      C  , ,���%�������%���G�������G�����������%����      C  , ,���s�������s���G������G����������s����      C  , ,���������������G���k���G���k������������      C  , ,�������������G�������G���������������      C  , ,���]�������]���G������G����������]����      C  , ,�����������������ԋ������ԋ����������      C  , ,���/������/����������������������/���      C  , ,���}������}�������'�������'������}���      C  , ,������������������u�������u����������      C  , ,����������������������������������      C  , ,���g������g��������������������g���      C  , ,����������������_�������_���������      C  , ,���}���m���}������'������'���m���}���m      C  , ,�������m����������u������u���m�������m      C  , ,������m��������������������m������m      C  , ,���g���m���g���������������m���g���m      C  , ,������m���������_������_���m������m      C  , ,���������������G��ܜ���G��ܜ������������      C  , ,���@�������@���G�������G�����������@����      C  , ,���������������G���8���G���8������������      C  , ,��٤������٤���G���N���G���N������٤����      C  , ,������m��������Ʒ�����Ʒ���m������m      C  , ,���[���m���[���������������m���[���m      C  , ,��ʩ���m��ʩ������S������S���m��ʩ���m      C  , ,��ɂ������ɂ���G���,���G���,������ɂ����      C  , ,�������������G��Ʒ���G��Ʒ�����������      C  , ,���[�������[���G������G����������[����      C  , ,��ʩ������ʩ���G���S���G���S������ʩ����      C  , ,���������������G��͡���G��͡������������      C  , ,���E�������E���G�������G�����������E����      C  , ,��ѓ������ѓ���G���=���G���=������ѓ����      C  , ,���������������G��ԋ���G��ԋ������������      C  , ,���/�������/���G�������G�����������/����      C  , ,���}�������}���G���'���G���'�������}����      C  , ,���������������G���u���G���u������������      C  , ,�������������G�������G���������������      C  , ,���g�������g���G������G����������g����      C  , ,�������������G���_���G���_�����������      C  , ,�������m���������͡�����͡���m�������m      C  , ,���E���m���E�����������������m���E���m      C  , ,��ѓ���m��ѓ������=������=���m��ѓ���m      C  , ,�������m���������ԋ�����ԋ���m�������m      C  , ,���/���m���/�����������������m���/���m      C  , ,���4�������4���G�������G�����������4����      C  , ,���������������Ʒ������Ʒ���������      C  , ,���[������[��������������������[���      C  , ,��ʩ�����ʩ�������S�������S�����ʩ���      C  , ,�����������������͡������͡����������      C  , ,���E������E����������������������E���      C  , ,��ѓ�����ѓ�������=�������=�����ѓ���      C  , ,���������������G���z���G���z������������      C  , ,�������������G�������G���������������      C  , ,���l�������l���G������G����������l����      C  , ,��Һ������Һ���G���d���G���d������Һ����      C  , ,�������������G��ղ���G��ղ�����������      C  , ,���V�������V���G��� ���G��� �������V����      C  , ,��ѓ���5��ѓ�������=�������=���5��ѓ���5      C  , ,�������5����������ԋ������ԋ���5�������5      C  , ,���/���5���/�������������������5���/���5      C  , ,���}���5���}�������'�������'���5���}���5      C  , ,�������5�����������u�������u���5�������5      C  , ,������5����������������������5������5      C  , ,���g���5���g�����������������5���g���5      C  , ,������5����������_�������_���5������5      C  , ,������5���������Ʒ������Ʒ���5������5      C  , ,�������������w��Ʒ���w��Ʒ�����������      C  , ,���[�������[���w������w����������[����      C  , ,��ʩ������ʩ���w���S���w���S������ʩ����      C  , ,���������������w��͡���w��͡������������      C  , ,���E�������E���w�������w�����������E����      C  , ,��ѓ������ѓ���w���=���w���=������ѓ����      C  , ,���������������w��ԋ���w��ԋ������������      C  , ,���/�������/���w�������w�����������/����      C  , ,���}�������}���w���'���w���'�������}����      C  , ,���������������w���u���w���u������������      C  , ,�������������w�������w���������������      C  , ,���g�������g���w������w����������g����      C  , ,�������������w���_���w���_�����������      C  , ,���[���5���[�����������������5���[���5      C  , ,������e��������Ʒ�����Ʒ���e������e      C  , ,���[���e���[���������������e���[���e      C  , ,��ʩ���e��ʩ������S������S���e��ʩ���e      C  , ,�������e���������͡�����͡���e�������e      C  , ,���E���e���E�����������������e���E���e      C  , ,��ѓ���e��ѓ������=������=���e��ѓ���e      C  , ,�������e���������ԋ�����ԋ���e�������e      C  , ,���/���e���/�����������������e���/���e      C  , ,���}���e���}������'������'���e���}���e      C  , ,�������e����������u������u���e�������e      C  , ,������e��������������������e������e      C  , ,���g���e���g���������������e���g���e      C  , ,������e���������_������_���e������e      C  , ,��ʩ���5��ʩ�������S�������S���5��ʩ���5      C  , ,����������������Ʒ������Ʒ�����������      C  , ,���[�������[���������������������[����      C  , ,��ʩ������ʩ�������S�������S������ʩ����      C  , ,������������������͡������͡������������      C  , ,���E�������E�����������������������E����      C  , ,��ѓ������ѓ�������=�������=������ѓ����      C  , ,������������������ԋ������ԋ������������      C  , ,���/�������/�����������������������/����      C  , ,���}�������}�������'�������'�������}����      C  , ,�������������������u�������u������������      C  , ,�������������������������������������      C  , ,���g�������g���������������������g����      C  , ,�����������������_�������_�����������      C  , ,�������5����������͡������͡���5�������5      C  , ,������������?��Ʒ���?��Ʒ���������      C  , ,���[������[���?������?���������[���      C  , ,��ʩ�����ʩ���?���S���?���S�����ʩ���      C  , ,��������������?��͡���?��͡����������      C  , ,���E������E���?�������?����������E���      C  , ,��ѓ�����ѓ���?���=���?���=�����ѓ���      C  , ,��������������?��ԋ���?��ԋ����������      C  , ,���/������/���?�������?����������/���      C  , ,���}������}���?���'���?���'������}���      C  , ,��������������?���u���?���u����������      C  , ,������������?�������?�������������      C  , ,���g������g���?������?���������g���      C  , ,������������?���_���?���_���������      C  , ,���E���5���E�������������������5���E���5      C  , ,������e���������3������3���e������e      C  , ,�������e�������������������e�������e      C  , ,���%���e���%�����������������e���%���e      C  , ,���s���e���s���������������e���s���e      C  , ,�������e����������k������k���e�������e      C  , ,������e��������������������e������e      C  , ,���]���e���]���������������e���]���e      C  , ,�������������w���I���w���I�����������      C  , ,���������������w������w���������������      C  , ,���;�������;���w�������w�����������;����      C  , ,�������������w���3���w���3�����������      C  , ,���������������w������w���������������      C  , ,���%�������%���w�������w�����������%����      C  , ,���s�������s���w������w����������s����      C  , ,���������������w���k���w���k������������      C  , ,�������������w�������w���������������      C  , ,���]�������]���w������w����������]����      C  , ,������5����������I�������I���5������5      C  , ,�������5���������������������5�������5      C  , ,���;���5���;�������������������5���;���5      C  , ,������5����������3�������3���5������5      C  , ,�����������������������������������      C  , ,���Q�������Q�����������������������Q����      C  , ,�����������������I�������I�����������      C  , ,��������������������������������������      C  , ,���;�������;�����������������������;����      C  , ,�����������������3�������3�����������      C  , ,��������������������������������������      C  , ,���%�������%�����������������������%����      C  , ,���s�������s���������������������s����      C  , ,�������������������k�������k������������      C  , ,�������������������������������������      C  , ,���]�������]���������������������]����      C  , ,�������5���������������������5�������5      C  , ,���%���5���%�������������������5���%���5      C  , ,���s���5���s�����������������5���s���5      C  , ,�������5�����������k�������k���5�������5      C  , ,������5����������������������5������5      C  , ,���]���5���]�����������������5���]���5      C  , ,������5��������������������5������5      C  , ,���Q���5���Q�������������������5���Q���5      C  , ,�������������w������w��������������      C  , ,���Q�������Q���w�������w�����������Q����      C  , ,������e������������������e������e      C  , ,���Q���e���Q�����������������e���Q���e      C  , ,������e���������I������I���e������e      C  , ,�������e�������������������e�������e      C  , ,������������?������?������������      C  , ,���Q������Q���?�������?����������Q���      C  , ,������������?���I���?���I���������      C  , ,��������������?������?�������������      C  , ,���;������;���?�������?����������;���      C  , ,������������?���3���?���3���������      C  , ,��������������?������?�������������      C  , ,���%������%���?�������?����������%���      C  , ,���s������s���?������?���������s���      C  , ,��������������?���k���?���k����������      C  , ,������������?�������?�������������      C  , ,���]������]���?������?���������]���      C  , ,���;���e���;�����������������e���;���e      C  , ,  z����  z���G  $���G  $����  z����      C  , ,  ����  �����   �����   ����  ����      C  , ,  "=���  "=����  "�����  "����  "=���      C  , ,  $����  $�����  %5����  %5���  $����      C  , ,  &����  &�����  '�����  '����  &����      C  , ,  )'���  )'����  )�����  )����  )'���      C  , ,  +u���  +u����  ,����  ,���  +u���      C  , ,  -����  -�����  .m����  .m���  -����      C  , ,  0���  0����  0�����  0����  0���      C  , ,  2_���  2_����  3	����  3	���  2_���      C  , ,  4����  4�����  5W����  5W���  4����      C  , ,  6����  6�����  7�����  7����  6����      C  , ,  9I���  9I����  9�����  9����  9I���      C  , ,  ����m  ����  K���  K���m  ����m      C  , ,  ����m  ����   ����   ����m  ����m      C  , ,  "=���m  "=���  "����  "����m  "=���m      C  , ,  $����m  $����  %5���  %5���m  $����m      C  , ,  &����m  &����  '����  '����m  &����m      C  , ,  )'���m  )'���  )����  )����m  )'���m      C  , ,  +u���m  +u���  ,���  ,���m  +u���m      C  , ,  -����m  -����  .m���  .m���m  -����m      C  , ,  0���m  0���  0����  0����m  0���m      C  , ,  2_���m  2_���  3	���  3	���m  2_���m      C  , ,  4����m  4����  5W���  5W���m  4����m      C  , ,  6����m  6����  7����  7����m  6����m      C  , ,  9I���m  9I���  9����  9����m  9I���m      C  , ,  �����  ����G  K���G  K����  �����      C  , ,  �����  ����G   ����G   �����  �����      C  , ,  "=����  "=���G  "����G  "�����  "=����      C  , ,  $�����  $����G  %5���G  %5����  $�����      C  , ,  &�����  &����G  '����G  '�����  &�����      C  , ,  )'����  )'���G  )����G  )�����  )'����      C  , ,  +u����  +u���G  ,���G  ,����  +u����      C  , ,  -�����  -����G  .m���G  .m����  -�����      C  , ,  0����  0���G  0����G  0�����  0����      C  , ,  2_����  2_���G  3	���G  3	����  2_����      C  , ,  4�����  4����G  5W���G  5W����  4�����      C  , ,  6�����  6����G  7����G  7�����  6�����      C  , ,  9I����  9I���G  9����G  9�����  9I����      C  , ,  ����  �����  K����  K���  ����      C  , ,  �����  ����G  r���G  r����  �����      C  , ,  !����  !���G  !����G  !�����  !����      C  , ,  #d����  #d���G  $���G  $����  #d����      C  , ,  %�����  %����G  &\���G  &\����  %�����      C  , ,  ( ����  ( ���G  (����G  (�����  ( ����      C  , ,  *N����  *N���G  *����G  *�����  *N����      C  , ,  ,�����  ,����G  -F���G  -F����  ,�����      C  , ,  .�����  .����G  /����G  /�����  .�����      C  , ,  18����  18���G  1����G  1�����  18����      C  , ,  3�����  3����G  40���G  40����  3�����      C  , ,  5�����  5����G  6~���G  6~����  5�����      C  , ,  8"����  8"���G  8����G  8�����  8"����      C  , ,  �����  ����G  	����G  	�����  �����      C  , ,  1����  1���G  ����G  �����  1����      C  , ,  ����  ���G  )���G  )����  ����      C  , ,  �����  ����G  w���G  w����  �����      C  , ,  ����  ���G  ����G  �����  ����      C  , ,  i����  i���G  ���G  ����  i����      C  , ,  �����  ����G  a���G  a����  �����      C  , ,  ����  ���G  ����G  �����  ����      C  , ,  S����  S���G  ����G  �����  S����      C  , ,  1���m  1���  ����  ����m  1���m      C  , ,  ���m  ���  )���  )���m  ���m      C  , ,  ����m  ����  w���  w���m  ����m      C  , ,  ���m  ���  ����  ����m  ���m      C  , ,  i���m  i���  ���  ���m  i���m      C  , ,  ����m  ����  a���  a���m  ����m      C  , ,  ���m  ���  ����  ����m  ���m      C  , ,  S���m  S���  ����  ����m  S���m      C  , ,  ���  ����  )����  )���  ���      C  , ,  ����  �����  w����  w���  ����      C  , ,  ���  ����  �����  ����  ���      C  , ,  i���  i����  ����  ���  i���      C  , ,  ����  �����  a����  a���  ����      C  , ,  �����  ����G  f���G  f����  �����      C  , ,  

����  

���G  
����G  
�����  

����      C  , ,  X����  X���G  ���G  ����  X����      C  , ,  �����  ����G  P���G  P����  �����      C  , ,  �����  ����G  ����G  �����  �����      C  , ,  B����  B���G  ����G  �����  B����      C  , ,  �����  ����G  :���G  :����  �����      C  , ,  �����  ����G  ����G  �����  �����      C  , ,  ,����  ,���G  ����G  �����  ,����      C  , ,  ���  ����  �����  ����  ���      C  , ,  S���  S����  �����  ����  S���      C  , ,  ����  �����  ?����  ?���  ����      C  , ,  ����  �����  	�����  	����  ����      C  , ,  1���  1����  �����  ����  1���      C  , ,  G���m  G���  ����  ����m  G���m      C  , ,  ����m  ����  ?���  ?���m  ����m      C  , ,  ����m  ����  	����  	����m  ����m      C  , ,   ����   ���G  ����G  �����   ����      C  , ,  n����  n���G  ���G  ����  n����      C  , ,  �����  ����G  ����G  �����  �����      C  , ,  G����  G���G  ����G  �����  G����      C  , ,  �����  ����G  ?���G  ?����  �����      C  , ,   �����   ����G  |���G  |����   �����      C  , ,  ����m  ����  ����  ����m  ����m      C  , ,  ����  �����  �����  ����  ����      C  , ,  G���  G����  �����  ����  G���      C  , ,  i���5  i����  ����  ���5  i���5      C  , ,  ����5  �����  a����  a���5  ����5      C  , ,  ���5  ����  �����  ����5  ���5      C  , ,  S���5  S����  �����  ����5  S���5      C  , ,  ����e  ����  ����  ����e  ����e      C  , ,  G���e  G���  ����  ����e  G���e      C  , ,  ����e  ����  ?���  ?���e  ����e      C  , ,  ����e  ����  	����  	����e  ����e      C  , ,  1���e  1���  ����  ����e  1���e      C  , ,  ���e  ���  )���  )���e  ���e      C  , ,  �����  �����  �����  �����  �����      C  , ,  G����  G����  �����  �����  G����      C  , ,  �����  �����  ?����  ?����  �����      C  , ,  �����  �����  	�����  	�����  �����      C  , ,  1����  1����  �����  �����  1����      C  , ,  ����  ����  )����  )����  ����      C  , ,  �����  �����  w����  w����  �����      C  , ,  ����  ����  �����  �����  ����      C  , ,  i����  i����  ����  ����  i����      C  , ,  �����  �����  a����  a����  �����      C  , ,  ����  ����  �����  �����  ����      C  , ,  S����  S����  �����  �����  S����      C  , ,  ����e  ����  w���  w���e  ����e      C  , ,  ���e  ���  ����  ����e  ���e      C  , ,  i���e  i���  ���  ���e  i���e      C  , ,  ����e  ����  a���  a���e  ����e      C  , ,  ���e  ���  ����  ����e  ���e      C  , ,  S���e  S���  ����  ����e  S���e      C  , ,  1���5  1����  �����  ����5  1���5      C  , ,  ���5  ����  )����  )���5  ���5      C  , ,  �����  ����w  ����w  �����  �����      C  , ,  G����  G���w  ����w  �����  G����      C  , ,  �����  ����w  ?���w  ?����  �����      C  , ,  �����  ����w  	����w  	�����  �����      C  , ,  1����  1���w  ����w  �����  1����      C  , ,  ����  ���w  )���w  )����  ����      C  , ,  �����  ����w  w���w  w����  �����      C  , ,  ����  ���w  ����w  �����  ����      C  , ,  i����  i���w  ���w  ����  i����      C  , ,  �����  ����w  a���w  a����  �����      C  , ,  ����  ���w  ����w  �����  ����      C  , ,  S����  S���w  ����w  �����  S����      C  , ,  ����5  �����  w����  w���5  ����5      C  , ,  ���5  ����  �����  ����5  ���5      C  , ,  ����5  �����  �����  ����5  ����5      C  , ,  G���5  G����  �����  ����5  G���5      C  , ,  ����5  �����  ?����  ?���5  ����5      C  , ,  ����5  �����  	�����  	����5  ����5      C  , ,  ����  ����?  ����?  ����  ����      C  , ,  G���  G���?  ����?  ����  G���      C  , ,  ����  ����?  ?���?  ?���  ����      C  , ,  ����  ����?  	����?  	����  ����      C  , ,  1���  1���?  ����?  ����  1���      C  , ,  ���  ���?  )���?  )���  ���      C  , ,  ����  ����?  w���?  w���  ����      C  , ,  ���  ���?  ����?  ����  ���      C  , ,  i���  i���?  ���?  ���  i���      C  , ,  ����  ����?  a���?  a���  ����      C  , ,  ���  ���?  ����?  ����  ���      C  , ,  S���  S���?  ����?  ����  S���      C  , ,  6����e  6����  7����  7����e  6����e      C  , ,  �����  �����  K����  K����  �����      C  , ,  �����  �����   �����   �����  �����      C  , ,  "=����  "=����  "�����  "�����  "=����      C  , ,  $�����  $�����  %5����  %5����  $�����      C  , ,  &�����  &�����  '�����  '�����  &�����      C  , ,  )'����  )'����  )�����  )�����  )'����      C  , ,  +u����  +u����  ,����  ,����  +u����      C  , ,  -�����  -�����  .m����  .m����  -�����      C  , ,  0����  0����  0�����  0�����  0����      C  , ,  2_����  2_����  3	����  3	����  2_����      C  , ,  4�����  4�����  5W����  5W����  4�����      C  , ,  6�����  6�����  7�����  7�����  6�����      C  , ,  9I����  9I����  9�����  9�����  9I����      C  , ,  9I���e  9I���  9����  9����e  9I���e      C  , ,  6����5  6�����  7�����  7����5  6����5      C  , ,  �����  ����w  K���w  K����  �����      C  , ,  �����  ����w   ����w   �����  �����      C  , ,  "=����  "=���w  "����w  "�����  "=����      C  , ,  $�����  $����w  %5���w  %5����  $�����      C  , ,  &�����  &����w  '����w  '�����  &�����      C  , ,  )'����  )'���w  )����w  )�����  )'����      C  , ,  +u����  +u���w  ,���w  ,����  +u����      C  , ,  -�����  -����w  .m���w  .m����  -�����      C  , ,  0����  0���w  0����w  0�����  0����      C  , ,  2_����  2_���w  3	���w  3	����  2_����      C  , ,  4�����  4����w  5W���w  5W����  4�����      C  , ,  6�����  6����w  7����w  7�����  6�����      C  , ,  9I����  9I���w  9����w  9�����  9I����      C  , ,  9I���5  9I����  9�����  9����5  9I���5      C  , ,  ����5  �����  K����  K���5  ����5      C  , ,  ����5  �����   �����   ����5  ����5      C  , ,  "=���5  "=����  "�����  "����5  "=���5      C  , ,  $����5  $�����  %5����  %5���5  $����5      C  , ,  &����5  &�����  '�����  '����5  &����5      C  , ,  )'���5  )'����  )�����  )����5  )'���5      C  , ,  +u���5  +u����  ,����  ,���5  +u���5      C  , ,  -����5  -�����  .m����  .m���5  -����5      C  , ,  0���5  0����  0�����  0����5  0���5      C  , ,  2_���5  2_����  3	����  3	���5  2_���5      C  , ,  4����5  4�����  5W����  5W���5  4����5      C  , ,  ����e  ����  K���  K���e  ����e      C  , ,  ����e  ����   ����   ����e  ����e      C  , ,  "=���e  "=���  "����  "����e  "=���e      C  , ,  $����e  $����  %5���  %5���e  $����e      C  , ,  &����e  &����  '����  '����e  &����e      C  , ,  )'���e  )'���  )����  )����e  )'���e      C  , ,  +u���e  +u���  ,���  ,���e  +u���e      C  , ,  -����e  -����  .m���  .m���e  -����e      C  , ,  0���e  0���  0����  0����e  0���e      C  , ,  2_���e  2_���  3	���  3	���e  2_���e      C  , ,  4����e  4����  5W���  5W���e  4����e      C  , ,  ����  ����?  K���?  K���  ����      C  , ,  ����  ����?   ����?   ����  ����      C  , ,  "=���  "=���?  "����?  "����  "=���      C  , ,  $����  $����?  %5���?  %5���  $����      C  , ,  &����  &����?  '����?  '����  &����      C  , ,  )'���  )'���?  )����?  )����  )'���      C  , ,  +u���  +u���?  ,���?  ,���  +u���      C  , ,  -����  -����?  .m���?  .m���  -����      C  , ,  0���  0���?  0����?  0����  0���      C  , ,  2_���  2_���?  3	���?  3	���  2_���      C  , ,  4����  4����?  5W���?  5W���  4����      C  , ,  6����  6����?  7����?  7����  6����      C  , ,  9I���  9I���?  9����?  9����  9I���      D   ,����  N����     s     s  N����  N      D   ,����������������   s����   s������������      D   ,  )  N  )          N  )  N      D   ,  w  N  w    ]    ]  N  w  N      D   ,  �  N  �    	�    	�  N  �  N      D   ,    N      �    �  N    N      D   ,  a  N  a    G    G  N  a  N      D   ,  �  N  �    �    �  N  �  N      D   ,  �  N  �    �    �  N  �  N      D   ,  K  N  K    1    1  N  K  N      D   ,  �  N  �          N  �  N      D   ,  �  N  �    �    �  N  �  N      D   ,  5  N  5          N  5  N      D   ,  �  N  �    i    i  N  �  N      D   ,  �  N  �     �     �  N  �  N      D   ,  "  N  "    #    #  N  "  N      D   ,  $m  N  $m    %S    %S  N  $m  N      D   ,  &�  N  &�    '�    '�  N  &�  N      D   ,  )	  N  )	    )�    )�  N  )	  N      D   ,  +W  N  +W    ,=    ,=  N  +W  N      D   ,  -�  N  -�    .�    .�  N  -�  N      D   ,  /�  N  /�    0�    0�  N  /�  N      D   ,  2A  N  2A    3'    3'  N  2A  N      D   ,  4�  N  4�    5u    5u  N  4�  N      D   ,  6�  N  6�    7�    7�  N  6�  N      D   ,  9+  N  9+    :    :  N  9+  N      D   ,   �   �   �  �  �  �  �   �   �   �      D   ,  �   �  �  �    �     �  �   �      D   ,  2   �  2  �  T  �  T   �  2   �      D   ,  �   �  �  �  �  �  �   �  �   �      D   ,  	�   �  	�  �  
�  �  
�   �  	�   �      D   ,     �    �  >  �  >   �     �      D   ,  j   �  j  �  �  �  �   �  j   �      D   ,  �   �  �  �  �  �  �   �  �   �      D   ,     �    �  (  �  (   �     �      D   ,  T   �  T  �  v  �  v   �  T   �      D   ,  �   �  �  �  �  �  �   �  �   �      D   ,  �   �  �  �    �     �  �   �      D   ,  >   �  >  �  `  �  `   �  >   �      D   ,  �   �  �  �  �  �  �   �  �   �      D   ,   �   �   �  �  !�  �  !�   �   �   �      D   ,  #(   �  #(  �  $J  �  $J   �  #(   �      D   ,  %v   �  %v  �  &�  �  &�   �  %v   �      D   ,  '�   �  '�  �  (�  �  (�   �  '�   �      D   ,  *   �  *  �  +4  �  +4   �  *   �      D   ,  ,`   �  ,`  �  -�  �  -�   �  ,`   �      D   ,  .�   �  .�  �  /�  �  /�   �  .�   �      D   ,  0�   �  0�  �  2  �  2   �  0�   �      D   ,  3J   �  3J  �  4l  �  4l   �  3J   �      D   ,  5�   �  5�  �  6�  �  6�   �  5�   �      D   ,  7�   �  7�  �  9  �  9   �  7�   �      D   ,  �  N  �    �    �  N  �  N      D   ,���F   ����F  ����h  ����h   ����F   �      D   ,��˔   ���˔  ���̶  ���̶   ���˔   �      D   ,����   �����  ����  ����   �����   �      D   ,���0   ����0  ����R  ����R   ����0   �      D   ,���~   ����~  ���Ӡ  ���Ӡ   ����~   �      D   ,����   �����  �����  �����   �����   �      D   ,���   ����  ����<  ����<   ����   �      D   ,���h   ����h  ���ڊ  ���ڊ   ����h   �      D   ,��۶   ���۶  �����  �����   ���۶   �      D   ,���   ����  ����&  ����&   ����   �      D   ,���R   ����R  ����t  ����t   ����R   �      D   ,���   ����  �����  �����   ����   �      D   ,����   �����  ����  ����   �����   �      D   ,���<   ����<  ����^  ����^   ����<   �      D   ,���   ����  ����  ����   ����   �      D   ,����   �����  �����  �����   �����   �      D   ,���&   ����&  ����H  ����H   ����&   �      D   ,���t   ����t  ����  ����   ����t   �      D   ,����   �����  �����  �����   �����   �      D   ,���   ����  ����2  ����2   ����   �      D   ,���^   ����^  �����  �����   ����^   �      D   ,����   �����  �����  �����   �����   �      D   ,����   �����  ����  ����   �����   �      D   ,���H   ����H  ����j  ����j   ����H   �      D   ,���=  N���=  ���#  ���#  N���=  N      D   ,��ʋ  N��ʋ  ���q  ���q  N��ʋ  N      D   ,����  N����  ��Ϳ  ��Ϳ  N����  N      D   ,���'  N���'  ���  ���  N���'  N      D   ,���u  N���u  ���[  ���[  N���u  N      D   ,����  N����  ��ԩ  ��ԩ  N����  N      D   ,���  N���  ����  ����  N���  N      D   ,���_  N���_  ���E  ���E  N���_  N      D   ,��ڭ  N��ڭ  ��ۓ  ��ۓ  N��ڭ  N      D   ,����  N����  ����  ����  N����  N      D   ,���I  N���I  ���/  ���/  N���I  N      D   ,���  N���  ���}  ���}  N���  N      D   ,����  N����  ����  ����  N����  N      D   ,���3  N���3  ���  ���  N���3  N      D   ,���  N���  ���g  ���g  N���  N      D   ,����  N����  ���  ���  N����  N      D   ,���  N���  ���  ���  N���  N      D   ,���k  N���k  ���Q  ���Q  N���k  N      D   ,���  N���  ���  ���  N���  N      D   ,���  N���  ����  ����  N���  N      D   ,���U  N���U  ���;  ���;  N���U  N      D   ,����  N����  ����  ����  N����  N      D   ,����  N����  ����  ����  N����  N      D   ,���?  N���?  ���%  ���%  N���?  N      D   ,����  N����  ����  ����  N����  N      D   ,����   �����  ����  ����   �����   �      D   ,���F������F���e���h���e���h������F���      D   ,��˔�����˔���e��̶���e��̶�����˔���      D   ,��������������e������e�������������      D   ,���0������0���e���R���e���R������0���      D   ,���~������~���e��Ӡ���e��Ӡ������~���      D   ,��������������e�������e��������������      D   ,������������e���<���e���<���������      D   ,���h������h���e��ڊ���e��ڊ������h���      D   ,��۶�����۶���e�������e���������۶���      D   ,������������e���&���e���&���������      D   ,���R������R���e���t���e���t������R���      D   ,������������e�������e�������������      D   ,��������������e������e�������������      D   ,���<������<���e���^���e���^������<���      D   ,������������e������e������������      D   ,��������������e�������e��������������      D   ,���&������&���e���H���e���H������&���      D   ,���t������t���e������e���������t���      D   ,��������������e�������e��������������      D   ,������������e���2���e���2���������      D   ,���^������^���e�������e����������^���      D   ,��������������e�������e��������������      D   ,��������������e������e�������������      D   ,���H������H���e���j���e���j������H���      D   ,����������������������������������������      D   ,���=�������=�������#�������#�������=����      D   ,��ʋ������ʋ�������q�������q������ʋ����      D   ,������������������Ϳ������Ϳ������������      D   ,���'�������'���������������������'����      D   ,���u�������u�������[�������[�������u����      D   ,������������������ԩ������ԩ������������      D   ,�������������������������������������      D   ,���_�������_�������E�������E�������_����      D   ,��ڭ������ڭ������ۓ������ۓ������ڭ����      D   ,����������������������������������������      D   ,���I�������I�������/�������/�������I����      D   ,�����������������}�������}�����������      D   ,����������������������������������������      D   ,���3�������3���������������������3����      D   ,�����������������g�������g�����������      D   ,��������������������������������������      D   ,�����������������������������������      D   ,���k�������k�������Q�������Q�������k����      D   ,�����������������������������������      D   ,�������������������������������������      D   ,���U�������U�������;�������;�������U����      D   ,����������������������������������������      D   ,����������������������������������������      D   ,���?�������?�������%�������%�������?����      D   ,��������������e������e�������������      D   ,  ����  ����e  ���e  ���  ����      D   ,  2���  2���e  T���e  T���  2���      D   ,  ����  ����e  ����e  ����  ����      D   ,  	����  	����e  
����e  
����  	����      D   ,  ���  ���e  >���e  >���  ���      D   ,  j���  j���e  ����e  ����  j���      D   ,  ����  ����e  ����e  ����  ����      D   ,  ���  ���e  (���e  (���  ���      D   ,  T���  T���e  v���e  v���  T���      D   ,  ����  ����e  ����e  ����  ����      D   ,  ����  ����e  ���e  ���  ����      D   ,  >���  >���e  `���e  `���  >���      D   ,  ����  ����e  ����e  ����  ����      D   ,   ����   ����e  !����e  !����   ����      D   ,  #(���  #(���e  $J���e  $J���  #(���      D   ,  %v���  %v���e  &����e  &����  %v���      D   ,  '����  '����e  (����e  (����  '����      D   ,  *���  *���e  +4���e  +4���  *���      D   ,  ,`���  ,`���e  -����e  -����  ,`���      D   ,  .����  .����e  /����e  /����  .����      D   ,  0����  0����e  2���e  2���  0����      D   ,  3J���  3J���e  4l���e  4l���  3J���      D   ,  5����  5����e  6����e  6����  5����      D   ,  7����  7����e  9���e  9���  7����      D   ,   ����   ����e  ����e  ����   ����      D   ,  �����  �����  �����  �����  �����      D   ,  )����  )����  ����  ����  )����      D   ,  w����  w����  ]����  ]����  w����      D   ,  �����  �����  	�����  	�����  �����      D   ,  ����  ����  �����  �����  ����      D   ,  a����  a����  G����  G����  a����      D   ,  �����  �����  �����  �����  �����      D   ,  �����  �����  �����  �����  �����      D   ,  K����  K����  1����  1����  K����      D   ,  �����  �����  ����  ����  �����      D   ,  �����  �����  �����  �����  �����      D   ,  5����  5����  ����  ����  5����      D   ,  �����  �����  i����  i����  �����      D   ,  �����  �����   �����   �����  �����      D   ,  "����  "����  #����  #����  "����      D   ,  $m����  $m����  %S����  %S����  $m����      D   ,  &�����  &�����  '�����  '�����  &�����      D   ,  )	����  )	����  )�����  )�����  )	����      D   ,  +W����  +W����  ,=����  ,=����  +W����      D   ,  -�����  -�����  .�����  .�����  -�����      D   ,  /�����  /�����  0�����  0�����  /�����      D   ,  2A����  2A����  3'����  3'����  2A����      D   ,  4�����  4�����  5u����  5u����  4�����      D   ,  6�����  6�����  7�����  7�����  6�����      D   ,  9+����  9+����  :����  :����  9+����      @   ,���������  M  <�  M  <����������     �     "�     " via_li_m1     C   ,      d       |    |   d      d      C  , ,   <   d   <     �     �   d   <   d      D   ,            r  |  r  |                �     "�     " "sky130_fd_pr__nfet_01v8_M4T2ST    �   ,���x������x  �  �  �  �������x���      A   ,���!���$���!  �  �  �  ����$���!���$      A  , ,���#  ����#  	B  �  	B  �  ����#  �      A  , ,���#���h���#  �����  ��������h���#���h      A  , ,  3���h  3  �  �  �  ����h  3���h      A  , ,���#�������#���h  ����h  ��������#����      ^   ,����  ����  	�  Z  	�  Z  ����        ^   ,������������  ���J  ���J������������      ^   ,  �����  �    Z    Z����  �����      ^   ,�������A��������  Z����  Z���A�������A      ]  , ,������������  Y  \  Y  \������������      B   ,���4  J���4  ����~  ����~  J���4  J      B   ,   �  J   �  �  �  �  �  J   �  J      B   ,���C�������C  J���o  J���o�������C����      B   ,   �����   �  J  �  J  �����   �����      B   ,���4���l���4�������~�������~���l���4���l      B   ,   ����l   �����  �����  ����l   ����l      B  , ,���  ����  	B����  	B����  ����  �      B  , ,���W  ����W  	B���  	B���  ����W  �      B  , ,����  �����  	B   U  	B   U  �����  �      B  , ,   �  �   �  	B  �  	B  �  �   �  �      B  , ,  S  �  S  	B  �  	B  �  �  S  �      B  , ,���#  O���#  �����  �����  O���#  O      B  , ,����  �����  D���.  D���.  �����  �      B  , ,   �  �   �  D  |  D  |  �   �  �      B  , ,  3  O  3  �  �  �  �  O  3  O      B  , ,���#  ����#  �����  �����  ����#  �      B  , ,  3  �  3  �  �  �  �  �  3  �      B  , ,���]  Q���]  ����  ����  Q���]  Q      B  , ,����  Q����  �   U  �   U  Q����  Q      B  , ,  �  Q  �  �  �  �  �  Q  �  Q      B  , ,���#  ����#  Q����  Q����  ����#  �      B  , ,  3  �  3  Q  �  Q  �  �  3  �      B  , ,���]  ����]  ����  ����  ����]  �      B  , ,����  �����  �   U  �   U  �����  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,���#  S���#  �����  �����  S���#  S      B  , ,  3  S  3  �  �  �  �  S  3  S      B  , ,���]  ����]  S���  S���  ����]  �      B  , ,����  �����  S   U  S   U  �����  �      B  , ,  �  �  �  S  �  S  �  �  �  �      B  , ,���#   ����#  �����  �����   ����#   �      B  , ,  3   �  3  �  �  �  �   �  3   �      B  , ,���]   U���]   ����   ����   U���]   U      B  , ,����   U����   �   U   �   U   U����   U      B  , ,  �   U  �   �  �   �  �   U  �   U      B  , ,���#�������#   U����   U�����������#����      B  , ,  3����  3   U  �   U  �����  3����      B  , ,���]������]��������������������]���      B  , ,���������������   U����   U����������      B  , ,  ����  �����  �����  ����  ����      B  , ,���#���W���#�����������������W���#���W      B  , ,  3���W  3���  ����  ����W  3���W      B  , ,���]�������]���W������W����������]����      B  , ,���������������W   U���W   U������������      B  , ,  �����  ����W  ����W  �����  �����      B  , ,���#������#����������������������#���      B  , ,  3���  3����  �����  ����  3���      B  , ,���]���Y���]���������������Y���]���Y      B  , ,�������Y�������   U���   U���Y�������Y      B  , ,  ����Y  ����  ����  ����Y  ����Y      B  , ,���#�������#���Y�������Y�����������#����      B  , ,  3����  3���Y  ����Y  �����  3����      B  , ,���]������]��������������������]���      B  , ,���������������   U����   U����������      B  , ,  ����  �����  �����  ����  ����      B  , ,���#���[���#�����������������[���#���[      B  , ,  3���[  3���  ����  ����[  3���[      B  , ,���#������#����������������������#���      B  , ,���������������f���.���f���.������������      B  , ,   �����   ����f  |���f  |����   �����      B  , ,  3���  3����  �����  ����  3���      B  , ,�������������h�������h���������������      B  , ,���W�������W���h������h����������W����      B  , ,���������������h   U���h   U������������      B  , ,   �����   ����h  ����h  �����   �����      B  , ,  S����  S���h  ����h  �����  S����      _   ,���   6���   �  �  �  �  6���   6      _   ,��� ���X��� ����  �����  ����X��� ���X      C   ,���#  ����#  	B  �  	B  �  ����#  �      C   ,���#���h���#  �����  ��������h���#���h      C   ,���4  ����4  D���~  D���~  ����4  �      C   ,   �  �   �  D  �  D  �  �   �  �      C   ,���]������]  ����  ����������]���      C   ,�����������  �   U  �   U����������      C   ,  ����  �  �  �  �  ����  ����      C   ,���4�������4���f���~���f���~�������4����      C   ,   �����   ����f  ����f  �����   �����      C   ,  3���h  3  �  �  �  ����h  3���h      C   ,���#�������#���h  ����h  ��������#����      C  , ,����  �����  D���.  D���.  �����  �      C  , ,   �  �   �  D  |  D  |  �   �  �      C  , ,���]  ����]  A���  A���  ����]  �      C  , ,����  �����  A   U  A   U  �����  �      C  , ,  �  �  �  A  �  A  �  �  �  �      C  , ,���]  /���]  ����  ����  /���]  /      C  , ,����  /����  �   U  �   U  /����  /      C  , ,  �  /  �  �  �  �  �  /  �  /      C  , ,���]  ����]  q���  q���  ����]  �      C  , ,����  �����  q   U  q   U  �����  �      C  , ,  �  �  �  q  �  q  �  �  �  �      C  , ,���]   _���]  	���  	���   _���]   _      C  , ,����   _����  	   U  	   U   _����   _      C  , ,  �   _  �  	  �  	  �   _  �   _      C  , ,���]�������]���������������������]����      C  , ,����������������   U����   U������������      C  , ,  �����  �����  �����  �����  �����      C  , ,���]�������]���9������9����������]����      C  , ,���������������9   U���9   U������������      C  , ,  �����  ����9  ����9  �����  �����      C  , ,���]���'���]�����������������'���]���'      C  , ,�������'��������   U����   U���'�������'      C  , ,  ����'  �����  �����  ����'  ����'      C  , ,���]�������]���i������i����������]����      C  , ,���������������i   U���i   U������������      C  , ,  �����  ����i  ����i  �����  �����      C  , ,���������������f���.���f���.������������      C  , ,   �����   ����f  |���f  |����   �����      D   ,���H  |���H  b���j  b���j  |���H  |      D   ,   �  |   �  b  �  b  �  |   �  |      D   ,���?���$���?  ����%  ����%���$���?���$      D   ,�������$����  �   s  �   s���$�������$      D   ,  ����$  �  �  �  �  ����$  ����$      D   ,���H�������H�������j�������j�������H����      D   ,   �����   �����  �����  �����   �����     �     "�     " opamp_v1 
  "sky130_fd_pr__nfet_01v8_M4T2ST   ���o�     via_li_m1   T    \���}e  ���}e  \���}e     via_li_m1   T    \���  ���  \���     via_li_m1   T    \���{�  ���{�  \���{�   
  "sky130_fd_pr__pfet_01v8_YCMRKB   �����   
  &sky130_fd_pr__cap_mim_m3_1_BLS9H9  �  B�        ����;   
  "sky130_fd_pr__nfet_01v8_8HUREQ   �h��ex   
  "sky130_fd_pr__nfet_01v8_8HUREQ   �b��ex   
  &sky130_fd_pr__cap_mim_m3_1_BLS9H9  �  B�        �����;   
  &sky130_fd_pr__cap_mim_m3_1_BLS9H9  �  B�        ^����;   
  "sky130_fd_pr__nfet_01v8_8JUMX6  a���_�   
  "sky130_fd_pr__pfet_01v8_YCMRKB   �����$   
  "sky130_fd_pr__pfet_01v8_YCMRKB   �����.   
  "sky130_fd_pr__pfet_01v8_YCMRKB   ��  	8   
  &sky130_fd_pr__cap_mim_m3_1_BLS9H9  �  B�        ^�����   
  &sky130_fd_pr__cap_mim_m3_1_BLS9H9  �  B�        �����   
  &sky130_fd_pr__cap_mim_m3_1_BLS9H9  �  B�        ������     via_li_m1   T    \�  3  �  3  \�  3     via_li_m1   T    \�  {  �  {  \�  {     via_li_m1   T    \�  �  �  �  \�  �   
  "sky130_fd_pr__pfet_01v8_YC9MKB   ��  .�   
  "sky130_fd_pr__pfet_01v8_YC9MKB   ��  .�   
  "sky130_fd_pr__pfet_01v8_YC9MKB   j�  .�     "sky130_fd_pr__pfet_01v8_YT7TV5     H  &p �  &p H  &p      E   , �  (� �  4D �  4D �  (� �  (�      E   ,  (i  $�  (i  ( �H  ( �H  $�  (i  $�      E   , �  � �  #� �  #� �  � �  �      E   ,  ]�����  ]���ޮ  ^���ޮ  ^�����  ]�����      E   ,  `����  `����  a+����  a+����  `����      E   ,  ba����  ba��ޮ  ce��ޮ  ce����  ba����      E   ,  d�����  d�����  e�����  e�����  d�����      E   ,  f�����  f���ޮ  h��ޮ  h����  f�����      E   ,  iK����  iK����  jc����  jc����  iK����      E   ,  k�����  k���ޮ  l���ޮ  l�����  k�����      E   ,  m�����  m�����  n�����  n�����  m�����      E   ,  p5����  p5��ޮ  q9��ޮ  q9����  p5����      E   ,  r�����  r�����  s�����  s�����  r�����      E   ,  t�����  t���ޮ  u���ޮ  u�����  t�����      E   ,  w����  w����  x7����  x7����  w����      E   ,  ym����  ym��ޮ  zq��ޮ  zq����  ym����      E   ,  {�����  {�����  |�����  |�����  {�����      E   ,  ~	����  ~	��ޮ  ��ޮ  ����  ~	����      E   ,  �W����  �W����  �o����  �o����  �W����      E   ,  ������  ����ޮ  ����ޮ  ������  ������      E   ,  ������  ������  �����  �����  ������      E   ,  �A����  �A��ޮ  �E��ޮ  �E����  �A����      E   ,  ������  ������  ������  ������  ������      E   ,  ������  ����ޮ  ����ޮ  ������  ������      E   ,  �+����  �+����  �C����  �C����  �+����      E   ,  �y����  �y��ޮ  �}��ޮ  �}����  �y����      E   ,  ������  ������  ������  ������  ������      E   ,  �����  ���ޮ  ���ޮ  �����  �����      E   ,  �c����  �c����  �{����  �{����  �c����      E   ,  ������  ����ޮ  ����ޮ  ������  ������      E   ,  ������  ������  �����  �����  ������      E   ,  �M����  �M��ޮ  �Q��ޮ  �Q����  �M����      E   ,  ������  ������  ������  ������  ������      E   ,  ������  ����ޮ  ����ޮ  ������  ������      E   ,  �7����  �7����  �O����  �O����  �7����      E   ,  ������  ����ޮ  ����ޮ  ������  ������      E   ,  ������  ������  ������  ������  ������      E   ,  �!����  �!��ޮ  �%��ޮ  �%����  �!����      E   ,  �o����  �o����  ������  ������  �o����      E   ,  ������  ����ޮ  ����ޮ  ������  ������      E   ,  �����  �����  �#����  �#����  �����      E   ,  �Y����  �Y��ޮ  �]��ޮ  �]����  �Y����      E   ,  ������  ������  ������  ������  ������      E   ,  ������  ����ޮ  ����ޮ  ������  ������      E   ,  �C����  �C����  �[����  �[����  �C����      E   ,  ������  ����ޮ  ����ޮ  ������  ������      E   ,  ������  ������  ������  ������  ������      E   ,  �-����  �-��ޮ  �1��ޮ  �1����  �-����      E   ,  �{����  �{����  Ɠ����  Ɠ����  �{����      E   ,  ������  ����ޮ  ����ޮ  ������  ������      E   ,  �����  �����  �/����  �/����  �����      E   ,  �e����  �e��ޮ  �i��ޮ  �i����  �e����      E   ,  γ����  γ����  ������  ������  γ����      E   ,  �����  ���ޮ  ���ޮ  �����  �����      E   ,  ����]�  ����aO ͐��aO ͐��]�  ����]�      E   , m�  � m�  #� n�  #� n�  � m�  �      E   , m�  (� m�  4D n�  4D n�  (� m�  (�      E   , �U  (� �U  4D �m  4D �m  (� �U  (�      E   , ��  (� ��  4D ��  4D ��  (� ��  (�      E   , ��  (� ��  4D �	  4D �	  (� ��  (�      E   , �I  (� �I  4D �M  4D �M  (� �I  (�      E   , ��  (� ��  4D ��  4D ��  (� ��  (�      E   , ��  (� ��  4D ��  4D ��  (� ��  (�      E   , �)  (� �)  4D �A  4D �A  (� �)  (�      E   , ��  (� ��  4D ��  4D ��  (� ��  (�      E   , ��  (� ��  4D ��  4D ��  (� ��  (�      E   , �  (� �  4D �!  4D �!  (� �  (�      E   , �a  (� �a  4D �y  4D �y  (� �a  (�      E   , ǹ  (� ǹ  4D Ƚ  4D Ƚ  (� ǹ  (�      E   , ��  (� ��  4D �  4D �  (� ��  (�      E   , �U  (� �U  4D �Y  4D �Y  (� �U  (�      E   , Ι  (� Ι  4D ϱ  4D ϱ  (� Ι  (�      E   , ��  (� ��  4D ��  4D ��  (� ��  (�      E   , p>  � p>  #� qV  #� qV  � p>  �      E   , r�  � r�  #� s�  #� s�  � r�  �      E   , t�  � t�  #� u�  #� u�  � t�  �      E   , w2  � w2  #� x6  #� x6  � w2  �      E   , yv  � yv  #� z�  #� z�  � yv  �      E   , {�  � {�  #� |�  #� |�  � {�  �      E   , ~  � ~  #� *  #� *  � ~  �      E   , �  � �  #� �	  #� �	  � �  �      E   , �I  � �I  #� �a  #� �a  � �I  �      E   , ��  � ��  #� ��  #� ��  � ��  �      E   , ��  � ��  #� ��  #� ��  � ��  �      E   , �=  � �=  #� �A  #� �A  � �=  �      E   , ��  � ��  #� ��  #� ��  � ��  �      E   , ��  � ��  #� ��  #� ��  � ��  �      E   , �  � �  #� �5  #� �5  � �  �      E   , �u  � �u  #� �y  #� �y  � �u  �      E   , ��  � ��  #� ��  #� ��  � ��  �      E   , �  � �  #� �  #� �  � �  �      E   , �U  � �U  #� �m  #� �m  � �U  �      E   , ��  � ��  #� ��  #� ��  � ��  �      E   , ��  � ��  #� �	  #� �	  � ��  �      E   , �I  � �I  #� �M  #� �M  � �I  �      E   , ��  � ��  #� ��  #� ��  � ��  �      E   , ��  � ��  #� ��  #� ��  � ��  �      E   , �)  � �)  #� �A  #� �A  � �)  �      E   , ��  � ��  #� ��  #� ��  � ��  �      E   , ��  � ��  #� ��  #� ��  � ��  �      E   , �  � �  #� �!  #� �!  � �  �      E   , �a  � �a  #� �y  #� �y  � �a  �      E   , ǹ  � ǹ  #� Ƚ  #� Ƚ  � ǹ  �      E   , ��  � ��  #� �  #� �  � ��  �      E   , �U  � �U  #� �Y  #� �Y  � �U  �      E   , Ι  � Ι  #� ϱ  #� ϱ  � Ι  �      E   , �  (� �  4D �  4D �  (� �  (�      E   , p>  (� p>  4D qV  4D qV  (� p>  (�      E   , r�  (� r�  4D s�  4D s�  (� r�  (�      E   , t�  (� t�  4D u�  4D u�  (� t�  (�      E   , w2  (� w2  4D x6  4D x6  (� w2  (�      E   , yv  (� yv  4D z�  4D z�  (� yv  (�      E   , {�  (� {�  4D |�  4D |�  (� {�  (�      E   , ~  (� ~  4D *  4D *  (� ~  (�      E   , �  (� �  4D �	  4D �	  (� �  (�      E   , �I  (� �I  4D �a  4D �a  (� �I  (�      E   , ��  (� ��  4D ��  4D ��  (� ��  (�      E   , ��  (� ��  4D ��  4D ��  (� ��  (�      E   , �=  (� �=  4D �A  4D �A  (� �=  (�      E   , ��  (� ��  4D ��  4D ��  (� ��  (�      E   , ��  (� ��  4D ��  4D ��  (� ��  (�      E   , �  (� �  4D �5  4D �5  (� �  (�      E   , �u  (� �u  4D �y  4D �y  (� �u  (�      E   ,   �   #� 3  #� 3  �   �      E   , s  � s  #� w  #� w  � s  �      E   , �  � �  #�  �  #�  �  � �  �      E   , "  � "  #� #  #� #  � "  �      E   , $S  � $S  #� %k  #� %k  � $S  �      E   , &�  � &�  #� '�  #� '�  � &�  �      E   , (�  � (�  #� *  #� *  � (�  �      E   , +G  � +G  #� ,K  #� ,K  � +G  �      E   , -�  � -�  #� .�  #� .�  � -�  �      E   , D~  � D~  #� E�  #� E�  � D~  �      E   , F�  � F�  #� G�  #� G�  � F�  �      E   , I  � I  #� J  #� J  � I  �      E   , K^  � K^  #� Lv  #� Lv  � K^  �      E   , M�  � M�  #� N�  #� N�  � M�  �      E   , O�  � O�  #� Q  #� Q  � O�  �      E   , RR  � RR  #� SV  #� SV  � RR  �      E   , T�  � T�  #� U�  #� U�  � T�  �      E   , V�  � V�  #� W�  #� W�  � V�  �      E   , Y2  � Y2  #� ZJ  #� ZJ  � Y2  �      E   , [�  � [�  #� \�  #� \�  � [�  �      E   , ]�  � ]�  #� ^�  #� ^�  � ]�  �      E   , `&  � `&  #� a*  #� a*  � `&  �      E   , �  (� �  4D 	�  4D 	�  (� �  (�      E   ,   (�   4D   4D   (�   (�      E   , G  (� G  4D _  4D _  (� G  (�      E   , �  (� �  4D �  4D �  (� �  (�      E   , �  (� �  4D �  4D �  (� �  (�      E   , ;  (� ;  4D ?  4D ?  (� ;  (�      E   ,   (�   4D �  4D �  (�   (�      E   , �  (� �  4D �  4D �  (� �  (�      E   ,   (�   4D 3  4D 3  (�   (�      E   , s  (� s  4D w  4D w  (� s  (�      E   , �  (� �  4D  �  4D  �  (� �  (�      E   , "  (� "  4D #  4D #  (� "  (�      E   , $S  (� $S  4D %k  4D %k  (� $S  (�      E   , &�  (� &�  4D '�  4D '�  (� &�  (�      E   , (�  (� (�  4D *  4D *  (� (�  (�      E   , +G  (� +G  4D ,K  4D ,K  (� +G  (�      E   , -�  (� -�  4D .�  4D .�  (� -�  (�      E   , D~  (� D~  4D E�  4D E�  (� D~  (�      E   , F�  (� F�  4D G�  4D G�  (� F�  (�      E   , I  (� I  4D J  4D J  (� I  (�      E   , K^  (� K^  4D Lv  4D Lv  (� K^  (�      E   , M�  (� M�  4D N�  4D N�  (� M�  (�      E   , O�  (� O�  4D Q  4D Q  (� O�  (�      E   , RR  (� RR  4D SV  4D SV  (� RR  (�      E   , T�  (� T�  4D U�  4D U�  (� T�  (�      E   , V�  (� V�  4D W�  4D W�  (� V�  (�      E   , Y2  (� Y2  4D ZJ  4D ZJ  (� Y2  (�      E   , [�  (� [�  4D \�  4D \�  (� [�  (�      E   , ]�  (� ]�  4D ^�  4D ^�  (� ]�  (�      E   , `&  (� `&  4D a*  4D a*  (� `&  (�      E   , bj  (� bj  4D c�  4D c�  (� bj  (�      E   , d�  (� d�  4D e�  4D e�  (� d�  (�      E   , g  (� g  4D h  4D h  (� g  (�      E   , i^  (� i^  4D jb  4D jb  (� i^  (�      E   , k�  (� k�  4D l�  4D l�  (� k�  (�      E   , bj  � bj  #� c�  #� c�  � bj  �      E   , d�  � d�  #� e�  #� e�  � d�  �      E   , g  � g  #� h  #� h  � g  �      E   , i^  � i^  #� jb  #� jb  � i^  �      E   , k�  � k�  #� l�  #� l�  � k�  �      E   ,   (�   4D '  4D '  (�   (�      E   , g  (� g  4D k  4D k  (� g  (�      E   ,   �   #� '  #� '  �   �      E   , g  � g  #� k  #� k  � g  �      E   , �  � �  #� 	�  #� 	�  � �  �      E   ,   �   #�   #�   �   �      E   , G  � G  #� _  #� _  � G  �      E   , �  � �  #� �  #� �  � �  �      E   , �  � �  #� �  #� �  � �  �      E   , ;  � ;  #� ?  #� ?  � ;  �      E   ,   �   #� �  #� �  �   �      E   , �  � �  #� �  #� �  � �  �      E   ,  P�  �  P�  
�  ��  
�  ��  �  P�  �      E   ,  P�����  P�  �  T  �  T����  P�����      E   ,  ]����  ]�  �  ^�  �  ^����  ]����      E   ,  ba���  ba  �  ce  �  ce���  ba���      E   ,  f����  f�  �  h  �  h���  f����      E   ,  k����  k�  �  l�  �  l����  k����      E   ,  p5���  p5  �  q9  �  q9���  p5���      E   ,  t����  t�  �  u�  �  u����  t����      E   ,  ym���  ym  �  zq  �  zq���  ym���      E   ,  ~	���  ~	  �    �  ���  ~	���      E   ,  �����  ��  �  ��  �  �����  �����      E   ,  �A���  �A  �  �E  �  �E���  �A���      E   ,  �����  ��  �  ��  �  �����  �����      E   ,  �y���  �y  �  �}  �  �}���  �y���      E   ,  ����  �  �  �  �  ����  ����      E   ,  �����  ��  �  ��  �  �����  �����      E   ,  �M���  �M  �  �Q  �  �Q���  �M���      E   ,  �����  ��  �  ��  �  �����  �����      E   ,  �����  ��  �  ��  �  �����  �����      E   ,  �!���  �!  �  �%  �  �%���  �!���      E   ,  �����  ��  �  ��  �  �����  �����      E   ,  �Y���  �Y  �  �]  �  �]���  �Y���      E   ,  �����  ��  �  ��  �  �����  �����      E   ,  �����  ��  �  ��  �  �����  �����      E   ,  �-���  �-  �  �1  �  �1���  �-���      E   ,  �����  ��  �  ��  �  �����  �����      E   ,  �e���  �e  �  �i  �  �i���  �e���      E   ,  ����  �  �  �  �  ����  ����      E   ,  P���ߏ  P�����  ������  ����ߏ  P���ߏ      E   ,  �  �  �  �  �  �  �  �  �  �      E   ,  �;  (�  �;  4D  �S  4D  �S  (�  �;  (�      E   ,  �����d  ��  �  ��  �  �����d  �����d      E   ,  ��  (�  ��  4D  ��  4D  ��  (�  ��  (�      E   ,  �[���d  �[  �  �s  �  �s���d  �[���d      E   ,  ��  (�  ��  4D  ��  4D  ��  (�  ��  (�      E   ,  �����d  ��  �  �  �  ����d  �����d      E   ,  �/  (�  �/  4D  �3  4D  �3  (�  �/  (�      E   ,  �����d  ��  �  ��  �  �����d  �����d      E   ,  �s  (�  �s  4D  �  4D  �  (�  �s  (�      E   ,  �/���d  �/  �  �G  �  �G���d  �/���d      E   ,  �O���d  �O  �  �g  �  �g���d  �O���d      E   ,  �����d  ��  �  ��  �  �����d  �����d      E   ,  ��  (�  ��  4D  ��  4D  ��  (�  ��  (�      E   ,  �g���d  �g  �  �  �  ����d  �g���d      E   ,  �����d  ��  �  �  �  ����d  �����d      E   ,  ����d  �  �  �  �  ����d  ����d      E   ,  �/  �  �/  #�  �3  #�  �3  �  �/  �      E   ,  Ο���d  Ο  �  Ϸ  �  Ϸ���d  Ο���d      E   ,  �����d  ��  �  ��  �  �����d  �����d      E   ,  �s  �  �s  #�  �  #�  �  �  �s  �      E   ,  �#���d  �#  �  �;  �  �;���d  �#���d      E   ,  �O  �  �O    �g    �g  �  �O  �      E   ,  ��  �  ��  �  ��  �  ��  �  ��  �      E   ,  ��  �  ��    �    �  �  ��  �      E   ,  �M  �  �M  �  �Q  �  �Q  �  �M  �      E   ,  ��  �  ��    ��    ��  �  ��  �      E   ,  ��  �  ��  �  ��  �  ��  �  ��  �      E   ,  �#  �  �#    �;    �;  �  �#  �      E   ,  ��  �  ��  �  ��  �  ��  �  ��  �      E   ,  ��  �  ��    ��    ��  �  ��  �      E   ,  �!  �  �!  �  �%  �  �%  �  �!  �      E   ,  �[  �  �[    �s    �s  �  �[  �      E   ,  ��  �  ��  �  ��  �  ��  �  ��  �      E   ,  ��  �  ��    �    �  �  ��  �      E   ,  �Y  �  �Y  �  �]  �  �]  �  �Y  �      E   ,  ��  �  ��    ��    ��  �  ��  �      E   ,  ��  �  ��  �  ��  �  ��  �  ��  �      E   ,  �/  �  �/    �G    �G  �  �/  �      E   ,  ��  �  ��  �  ��  �  ��  �  ��  �      E   ,  ��  �  ��    ��    ��  �  ��  �      E   ,  �-  �  �-  �  �1  �  �1  �  �-  �      E   ,  �g  �  �g    �    �  �  �g  �      E   ,  ��  �  ��  �  ��  �  ��  �  ��  �      E   ,  �  �  �    �    �  �  �  �      E   ,  �e  �  �e  �  �i  �  �i  �  �e  �      E   ,  Ο  �  Ο    Ϸ    Ϸ  �  Ο  �      E   ,  �  �  �  �  �  �  �  �  �  �      E   ,  ��  �  ��  #�  ��  #�  ��  �  ��  �      E   ,  �;  �  �;  #�  �S  #�  �S  �  �;  �      E   ,  ��  �  ��  #�  ��  #�  ��  �  ��  �      E   ,  ��  �  ��  #�  ��  #�  ��  �  ��  �      E   ,  �A  �  �A  �  �E  �  �E  �  �A  �      E   ,  �{  �  �{    ��    ��  �  �{  �      E   ,  ��  �  ��  �  ��  �  ��  �  ��  �      E   ,  �  �  �    �/    �/  �  �  �      E   ,  �y  �  �y  �  �}  �  �}  �  �y  �      E   ,  ��  �  ��    ��    ��  �  ��  �      E   ,  _�  �  _�    a    a  �  _�  �      E   ,  ����d  �  �  �/  �  �/���d  ����d      E   ,  m����d  m�  �  n�  �  n����d  m����d      E   ,  �����d  ��  �  ��  �  �����d  �����d      E   ,  ba  �  ba  �  ce  �  ce  �  ba  �      E   ,  ro���d  ro  �  s�  �  s����d  ro���d      E   ,  _����d  _�  �  a  �  a���d  _����d      E   ,  w���d  w  �  x#  �  x#���d  w���d      E   ,  P�  
�  P�  
�  ^�  
�  ^�  
�  P�  
�      E   ,  {����d  {�  �  |�  �  |����d  {����d      E   ,  d����d  d�  �  e�  �  e����d  d����d      E   ,  �C���d  �C  �  �[  �  �[���d  �C���d      E   ,  ]�  �  ]�  �  ^�  �  ^�  �  ]�  �      E   ,  �����d  ��  �  ��  �  �����d  �����d      E   ,  i7���d  i7  �  jO  �  jO���d  i7���d      E   ,  �{���d  �{  �  ��  �  �����d  �{���d      E   ,  d�  �  d�    e�    e�  �  d�  �      E   ,  f�  �  f�  �  h  �  h  �  f�  �      E   ,  i7  �  i7    jO    jO  �  i7  �      E   ,  k�  �  k�  �  l�  �  l�  �  k�  �      E   ,  m�  �  m�    n�    n�  �  m�  �      E   ,  p5  �  p5  �  q9  �  q9  �  p5  �      E   ,  ro  �  ro    s�    s�  �  ro  �      E   ,  t�  �  t�  �  u�  �  u�  �  t�  �      E   ,  w  �  w    x#    x#  �  w  �      E   ,  ym  �  ym  �  zq  �  zq  �  ym  �      E   ,  {�  �  {�    |�    |�  �  {�  �      E   ,  ~	  �  ~	  �    �    �  ~	  �      E   ,  �C  �  �C    �[    �[  �  �C  �      E   ,  ��  �  ��  �  ��  �  ��  �  ��  �      E   ,  ��  �  ��    ��    ��  �  ��  �      E   ,  m����Z  m���ޮ  n���ޮ  n����Z  m����Z      E   ,  �{���  �{���  �����  �����  �{���      E   ,  d����  d����  e����  e����  d����      E   ,  ro���Z  ro��ޮ  s���ޮ  s����Z  ro���Z      E   ,  m����  m����  n����  n����  m����      E   ,  ����  ����  �/���  �/���  ����      E   ,  w���Z  w��ޮ  x#��ޮ  x#���Z  w���Z      E   ,  {����  {����  |����  |����  {����      E   ,  _����  _����  a���  a���  _����      E   ,  {����Z  {���ޮ  |���ޮ  |����Z  {����Z      E   ,  P�����  P�����  ^�����  ^�����  P�����      E   ,  �����  �����  �����  �����  �����      E   ,  �C���Z  �C��ޮ  �[��ޮ  �[���Z  �C���Z      E   ,  ;8����  ;8����  T����  T����  ;8����      E   ,  _����Z  _���ޮ  a��ޮ  a���Z  _����Z      E   ,  �����Z  ����ޮ  ����ޮ  �����Z  �����Z      E   ,  �C���  �C���  �[���  �[���  �C���      E   ,  ro���  ro���  s����  s����  ro���      E   ,  �{���Z  �{��ޮ  ����ޮ  �����Z  �{���Z      E   ,  d����Z  d���ޮ  e���ޮ  e����Z  d����Z      E   ,  i7���  i7���  jO���  jO���  i7���      E   ,  ����Z  ���ޮ  �/��ޮ  �/���Z  ����Z      E   ,  �����  �����  �����  �����  �����      E   ,  i7���Z  i7��ޮ  jO��ޮ  jO���Z  i7���Z      E   ,  �����Z  ����ޮ  ����ޮ  �����Z  �����Z      E   ,  P�����  P�����  T����  T����  P�����      E   ,  w���  w���  x#���  x#���  w���      E   ,  �#���  �#���  �;���  �;���  �#���      E   ,  �[���Z  �[��ޮ  �s��ޮ  �s���Z  �[���Z      E   ,  �[���  �[���  �s���  �s���  �[���      E   ,  Ο���  Ο���  Ϸ���  Ϸ���  Ο���      E   ,  �����Z  ����ޮ  ���ޮ  ����Z  �����Z      E   ,  �/���  �/���  �G���  �G���  �/���      E   ,  �O���Z  �O��ޮ  �g��ޮ  �g���Z  �O���Z      E   ,  �����Z  ����ޮ  ����ޮ  �����Z  �����Z      E   ,  �����  �����  �����  �����  �����      E   ,  �O���  �O���  �g���  �g���  �O���      E   ,  �/���Z  �/��ޮ  �G��ޮ  �G���Z  �/���Z      E   ,  �����Z  ����ޮ  ���ޮ  ����Z  �����Z      E   ,  �����  �����  �����  �����  �����      E   ,  �����Z  ����ޮ  ����ޮ  �����Z  �����Z      E   ,  �����  �����  ����  ����  �����      E   ,  �����Z  ����ޮ  ����ޮ  �����Z  �����Z      E   ,  �g���Z  �g��ޮ  ���ޮ  ����Z  �g���Z      E   ,  �����  �����  �����  �����  �����      E   ,  �g���  �g���  ����  ����  �g���      E   ,  ����Z  ���ޮ  ���ޮ  ����Z  ����Z      E   ,  �#���Z  �#��ޮ  �;��ޮ  �;���Z  �#���Z      E   ,  �����  �����  ����  ����  �����      E   ,  Ο���Z  Ο��ޮ  Ϸ��ޮ  Ϸ���Z  Ο���Z      E   ,  �����  �����  �����  �����  �����      E   ,  �����Z  ����ޮ  ����ޮ  �����Z  �����Z      E   ,  ����  ����  ����  ����  ����      E   ,  P�����  P�����  ������  ������  P�����      E   ,  �����  �����  �����  �����  �����      E   ,  P����{  P�����  ������  �����{  P����{      E   ,  ]���{{  ]�����  ^�����  ^���{{  ]���{{      E   ,  `���F  `����  a+����  a+���F  `���F      E   ,  ba��{{  ba����  ce����  ce��{{  ba��{{      E   ,  d����F  d�����  e�����  e����F  d����F      E   ,  f���{{  f�����  h����  h��{{  f���{{      E   ,  iK���F  iK����  jc����  jc���F  iK���F      E   ,  k���{{  k�����  l�����  l���{{  k���{{      E   ,  m����F  m�����  n�����  n����F  m����F      E   ,  p5��{{  p5����  q9����  q9��{{  p5��{{      E   ,  r����F  r�����  s�����  s����F  r����F      E   ,  t���{{  t�����  u�����  u���{{  t���{{      E   ,  w���F  w����  x7����  x7���F  w���F      E   ,  ym��{{  ym����  zq����  zq��{{  ym��{{      E   ,  {����F  {�����  |�����  |����F  {����F      E   ,  ~	��{{  ~	����  ����  ��{{  ~	��{{      E   ,  �W���F  �W����  �o����  �o���F  �W���F      E   ,  ����{{  ������  ������  ����{{  ����{{      E   ,  �����F  ������  �����  ����F  �����F      E   ,  �A��{{  �A����  �E����  �E��{{  �A��{{      E   ,  �����F  ������  ������  �����F  �����F      E   ,  ����{{  ������  ������  ����{{  ����{{      E   ,  �+���F  �+����  �C����  �C���F  �+���F      E   ,  �y��{{  �y����  �}����  �}��{{  �y��{{      E   ,  �����F  ������  ������  �����F  �����F      E   ,  ���{{  �����  �����  ���{{  ���{{      E   ,  �c���F  �c����  �{����  �{���F  �c���F      E   ,  ����{{  ������  ������  ����{{  ����{{      E   ,  �����F  ������  �����  ����F  �����F      E   ,  �M��{{  �M����  �Q����  �Q��{{  �M��{{      E   ,  �����F  ������  ������  �����F  �����F      E   ,  ����{{  ������  ������  ����{{  ����{{      E   ,  �7���F  �7����  �O����  �O���F  �7���F      E   ,  ����{{  ������  ������  ����{{  ����{{      E   ,  �����F  ������  ������  �����F  �����F      E   ,  �!��{{  �!����  �%����  �%��{{  �!��{{      E   ,  �o���F  �o����  ������  �����F  �o���F      E   ,  ����{{  ������  ������  ����{{  ����{{      E   ,  ����F  �����  �#����  �#���F  ����F      E   ,  �Y��{{  �Y����  �]����  �]��{{  �Y��{{      E   ,  �����F  ������  ������  �����F  �����F      E   ,  ����{{  ������  ������  ����{{  ����{{      E   ,  �C���F  �C����  �[����  �[���F  �C���F      E   ,  ����{{  ������  ������  ����{{  ����{{      E   ,  �����F  ������  ������  �����F  �����F      E   ,  �-��{{  �-����  �1����  �1��{{  �-��{{      E   ,  �{���F  �{����  Ɠ����  Ɠ���F  �{���F      E   ,  ����{{  ������  ������  ����{{  ����{{      E   ,  ����F  �����  �/����  �/���F  ����F      E   ,  �e��{{  �e����  �i����  �i��{{  �e��{{      E   ,  γ���F  γ����  ������  �����F  γ���F      E   ,  ���{{  �����  �����  ���{{  ���{{      E   ,  ���g+  ���s  �7��s  �7��g+  ���g+      E   ,  s���c�  s���g+  �=��g+  �=��c�  s���c�      E   ,  ���W�  ���c�  �7��c�  �7��W�  ���W�      E   ,  �o����  �o����  ������  ������  �o����      E   ,  ������  ������  ������  ������  ������      E   ,  ����P  �����  �#����  �#���P  ����P      E   ,  �����  �����  �#����  �#����  �����      E   ,  �Y����  �Y����  �]����  �]����  �Y����      E   ,  �����P  ������  ������  �����P  �����P      E   ,  ������  ������  ������  ������  ������      E   ,  ������  ������  ������  ������  ������      E   ,  �C���P  �C����  �[����  �[���P  �C���P      E   ,  �C����  �C����  �[����  �[����  �C����      E   ,  ������  ������  ������  ������  ������      E   ,  �����P  ������  ������  �����P  �����P      E   ,  ������  ������  ������  ������  ������      E   ,  �-����  �-����  �1����  �1����  �-����      E   ,  �{���P  �{����  Ɠ����  Ɠ���P  �{���P      E   ,  �{����  �{����  Ɠ����  Ɠ����  �{����      E   ,  ������  ������  ������  ������  ������      E   ,  ����P  �����  �/����  �/���P  ����P      E   ,  �����  �����  �/����  �/����  �����      E   ,  �e����  �e����  �i����  �i����  �e����      E   ,  γ���P  γ����  ������  �����P  γ���P      E   ,  γ����  γ����  ������  ������  γ����      E   ,  �����  �����  �����  �����  �����      E   ,  �c���P  �c����  �{����  �{���P  �c���P      E   ,  �c����  �c����  �{����  �{����  �c����      E   ,  ������  ������  ������  ������  ������      E   ,  �����P  ������  �����  ����P  �����P      E   ,  ������  ������  �����  �����  ������      E   ,  �M����  �M����  �Q����  �Q����  �M����      E   ,  �����P  ������  ������  �����P  �����P      E   ,  ������  ������  ������  ������  ������      E   ,  ������  ������  ������  ������  ������      E   ,  �7���P  �7����  �O����  �O���P  �7���P      E   ,  �7����  �7����  �O����  �O����  �7����      E   ,  ������  ������  ������  ������  ������      E   ,  �����P  ������  ������  �����P  �����P      E   ,  ������  ������  ������  ������  ������      E   ,  �!����  �!����  �%����  �%����  �!����      E   ,  �o���P  �o����  ������  �����P  �o���P      E   ,  r����P  r�����  s�����  s����P  r����P      E   ,  r�����  r�����  s�����  s�����  r�����      E   ,  t�����  t�����  u�����  u�����  t�����      E   ,  w���P  w����  x7����  x7���P  w���P      E   ,  w����  w����  x7����  x7����  w����      E   ,  ym����  ym����  zq����  zq����  ym����      E   ,  {����P  {�����  |�����  |����P  {����P      E   ,  {�����  {�����  |�����  |�����  {�����      E   ,  ~	����  ~	����  ����  ����  ~	����      E   ,  �W���P  �W����  �o����  �o���P  �W���P      E   ,  �W����  �W����  �o����  �o����  �W����      E   ,  ������  ������  ������  ������  ������      E   ,  �����P  ������  �����  ����P  �����P      E   ,  ������  ������  �����  �����  ������      E   ,  �A����  �A����  �E����  �E����  �A����      E   ,  �����P  ������  ������  �����P  �����P      E   ,  ������  ������  ������  ������  ������      E   ,  ������  ������  ������  ������  ������      E   ,  �+���P  �+����  �C����  �C���P  �+���P      E   ,  �+����  �+����  �C����  �C����  �+����      E   ,  �y����  �y����  �}����  �}����  �y����      E   ,  �����P  ������  ������  �����P  �����P      E   ,  ������  ������  ������  ������  ������      E   ,  P�����  P�����  T����  T����  P�����      E   ,  P�����  P�����  b9����  b9����  P�����      E   ,  ;8����  ;8����  T����  T����  ;8����      E   ,  P�����  P�����  T����  T����  P�����      E   ,  ]�����  ]�����  ^�����  ^�����  ]�����      E   ,  `���P  `����  a+����  a+���P  `���P      E   ,  `����  `����  a+����  a+����  `����      E   ,  ba����  ba����  ce����  ce����  ba����      E   ,  d����P  d�����  e�����  e����P  d����P      E   ,  d�����  d�����  e�����  e�����  d�����      E   ,  f�����  f�����  h����  h����  f�����      E   ,  iK���P  iK����  jc����  jc���P  iK���P      E   ,  iK����  iK����  jc����  jc����  iK����      E   ,  k�����  k�����  l�����  l�����  k�����      E   ,  m����P  m�����  n�����  n����P  m����P      E   ,  m�����  m�����  n�����  n�����  m�����      E   ,  p5����  p5����  q9����  q9����  p5����      E   ,  P�����  P�����  ^�����  ^�����  P�����      E   ,  w3��g�  w3��s  x7��s  x7��g�  w3��g�      E   ,  yw��g+  yw��s  z���s  z���g+  yw��g+      E   ,  {���g�  {���s  |���s  |���g�  {���g�      E   ,  ~��g+  ~��s  +��s  +��g+  ~��g+      E   ,  �k��g�  �k��s  �o��s  �o��g�  �k��g�      E   ,  ����g+  ����s  ����s  ����g+  ����g+      E   ,  ���g�  ���s  ���s  ���g�  ���g�      E   ,  �K��g+  �K��s  �c��s  �c��g+  �K��g+      E   ,  ����g�  ����s  ����s  ����g�  ����g�      E   ,  ����g+  ����s  ����s  ����g+  ����g+      E   ,  �?��g�  �?��s  �C��s  �C��g�  �?��g�      E   ,  ����g+  ����s  ����s  ����g+  ����g+      E   ,  ����g�  ����s  ����s  ����g�  ����g�      E   ,  J���o�  J���{S  K���{S  K���o�  J���o�      E   ,  N���o�  N���{S  O���{S  O���o�  N���o�      E   ,  r���W�  r���c%  s���c%  s���W�  r���W�      E   ,  t���W�  t���c�  u���c�  u���W�  t���W�      E   ,  w3��W�  w3��c%  x7��c%  x7��W�  w3��W�      E   ,  yw��W�  yw��c�  z���c�  z���W�  yw��W�      E   ,  {���W�  {���c%  |���c%  |���W�  {���W�      E   ,  ~��W�  ~��c�  +��c�  +��W�  ~��W�      E   ,  �k��W�  �k��c%  �o��c%  �o��W�  �k��W�      E   ,  ����W�  ����c�  ����c�  ����W�  ����W�      E   ,  ���W�  ���c%  ���c%  ���W�  ���W�      E   ,  �K��W�  �K��c�  �c��c�  �c��W�  �K��W�      E   ,  ����W�  ����c%  ����c%  ����W�  ����W�      E   ,  ����W�  ����c�  ����c�  ����W�  ����W�      E   ,  �?��W�  �?��c%  �C��c%  �C��W�  �?��W�      E   ,  ����W�  ����c�  ����c�  ����W�  ����W�      E   ,  ����W�  ����c%  ����c%  ����W�  ����W�      E   ,  r���g�  r���s  s���s  s���g�  r���g�      E   ,  t���g+  t���s  u���s  u���g+  t���g+      E   ,  �9��g�  �9��s  �=��s  �=��g�  �9��g�      E   ,  �}��g�  �}��s  ����s  ����g�  �}��g�      E   ,  ����g�  ����s  ����s  ����g�  ����g�      E   ,  ���g�  ���s  �1��s  �1��g�  ���g�      E   ,  �q��g�  �q��s  �u��s  �u��g�  �q��g�      E   ,  ����g�  ����s  ����s  ����g�  ����g�      E   ,  ���g�  ���s  ���s  ���g�  ���g�      E   ,  �Q��g�  �Q��s  �i��s  �i��g�  �Q��g�      E   ,  ����g�  ����s  ����s  ����g�  ����g�      E   ,  ����g�  ����s  ���s  ���g�  ����g�      E   ,  �E��g�  �E��s  �I��s  �I��g�  �E��g�      E   ,  ����g�  ����s  ����s  ����g�  ����g�      E   ,  ����g�  ����s  ����s  ����g�  ����g�      E   ,  �%��g�  �%��s  �=��s  �=��g�  �%��g�      E   ,  ����g�  ����s  ����s  ����g�  ����g�      E   ,  ����W�  ����c%  ����c%  ����W�  ����W�      E   ,  ����W�  ����c%  ����c%  ����W�  ����W�      E   ,  �9��W�  �9��c%  �=��c%  �=��W�  �9��W�      E   ,  �}��W�  �}��c%  ����c%  ����W�  �}��W�      E   ,  ����W�  ����c%  ����c%  ����W�  ����W�      E   ,  ���W�  ���c%  �1��c%  �1��W�  ���W�      E   ,  �q��W�  �q��c%  �u��c%  �u��W�  �q��W�      E   ,  ����W�  ����c%  ����c%  ����W�  ����W�      E   ,  ���W�  ���c%  ���c%  ���W�  ���W�      E   ,  �Q��W�  �Q��c%  �i��c%  �i��W�  �Q��W�      E   ,  ����W�  ����c%  ����c%  ����W�  ����W�      E   ,  ����W�  ����c%  ���c%  ���W�  ����W�      E   ,  �E��W�  �E��c%  �I��c%  �I��W�  �E��W�      E   ,  ����W�  ����c%  ����c%  ����W�  ����W�      E   ,  ����W�  ����c%  ����c%  ����W�  ����W�      E   ,  �%��W�  �%��c%  �=��c%  �=��W�  �%��W�      E   ,  ����bg  ����s3  ����s3  ����bg  ����bg      E   ,  �{��bg  �{��s3  ����s3  ����bg  �{��bg      E   ,  �_��bg  �_��s3  �w��s3  �w��bg  �_��bg      E   ,  �C��bg  �C��s3  �[��s3  �[��bg  �C��bg      E   ,  '��bg  '��s3 ?��s3 ?��bg  '��bg      E   ,  ����g�  ����s  ����s  ����g�  ����g�      E   ,  ����L  ����\�  ����\�  ����L  ����L      E   ,  �{��L  �{��\�  ����\�  ����L  �{��L      E   ,  �_��L  �_��\�  �w��\�  �w��L  �_��L      E   ,  �C��L  �C��\�  �[��\�  �[��L  �C��L      E   ,  '��L  '��\� ?��\� ?��L  '��L      E   , m���bg m���s3 o��s3 o��bg m���bg      E   , m���L m���\� o��\� o��L m���L      E   , +��bg +��s3 C��s3 C��bg +��bg      E   , ��bg ��s3 '��s3 '��bg ��bg      E   , ���bg ���s3 !��s3 !��bg ���bg      E   , "���bg "���s3 #���s3 #���bg "���bg      E   , %���bg %���s3 &���s3 &���bg %���bg      E   , (���bg (���s3 )���s3 )���bg (���bg      E   , +���bg +���s3 ,���s3 ,���bg +���bg      E   , .g��bg .g��s3 /��s3 /��bg .g��bg      E   , 1K��bg 1K��s3 2c��s3 2c��bg 1K��bg      E   , 4/��bg 4/��s3 5G��s3 5G��bg 4/��bg      E   , 7��bg 7��s3 8+��s3 8+��bg 7��bg      E   , 9���bg 9���s3 ;��s3 ;��bg 9���bg      E   , <���bg <���s3 =���s3 =���bg <���bg      E   , ?���bg ?���s3 @���s3 @���bg ?���bg      E   , B���bg B���s3 C���s3 C���bg B���bg      E   , E���bg E���s3 F���s3 F���bg E���bg      E   , Hk��bg Hk��s3 I���s3 I���bg Hk��bg      E   , KO��bg KO��s3 Lg��s3 Lg��bg KO��bg      E   , N3��bg N3��s3 OK��s3 OK��bg N3��bg      E   , Q��bg Q��s3 R/��s3 R/��bg Q��bg      E   , S���bg S���s3 U��s3 U��bg S���bg      E   , V���bg V���s3 W���s3 W���bg V���bg      E   , Y���bg Y���s3 Z���s3 Z���bg Y���bg      E   , \���bg \���s3 ]���s3 ]���bg \���bg      E   , _���bg _���s3 `���s3 `���bg _���bg      E   , bo��bg bo��s3 c���s3 c���bg bo��bg      E   , eS��bg eS��s3 fk��s3 fk��bg eS��bg      E   , h7��bg h7��s3 iO��s3 iO��bg h7��bg      E   , k��bg k��s3 l3��s3 l3��bg k��bg      E   , c��bg c��s3 {��s3 {��bg c��bg      E   , ��bg ��s3 #��s3 #��bg ��bg      E   , ���bg ���s3 ��s3 ��bg ���bg      E   , ���bg ���s3 	���s3 	���bg ���bg      E   , ���bg ���s3 ���s3 ���bg ���bg      E   , ���bg ���s3 ���s3 ���bg ���bg      E   , ��bg ��s3 ���s3 ���bg ��bg      E   , ��L ��\� #��\� #��L ��L      E   , ���L ���\� ��\� ��L ���L      E   , ���L ���\� 	���\� 	���L ���L      E   , ���L ���\� ���\� ���L ���L      E   , ���L ���\� ���\� ���L ���L      E   , ��L ��\� ���\� ���L ��L      E   , c��L c��\� {��\� {��L c��L      E   , G��L G��\� _��\� _��L G��L      E   , +��L +��\� C��\� C��L +��L      E   , ��L ��\� '��\� '��L ��L      E   , ���L ���\� !��\� !��L ���L      E   , "���L "���\� #���\� #���L "���L      E   , %���L %���\� &���\� &���L %���L      E   , (���L (���\� )���\� )���L (���L      E   , +���L +���\� ,���\� ,���L +���L      E   , .g��L .g��\� /��\� /��L .g��L      E   , 1K��L 1K��\� 2c��\� 2c��L 1K��L      E   , 4/��L 4/��\� 5G��\� 5G��L 4/��L      E   , 7��L 7��\� 8+��\� 8+��L 7��L      E   , 9���L 9���\� ;��\� ;��L 9���L      E   , <���L <���\� =���\� =���L <���L      E   , ?���L ?���\� @���\� @���L ?���L      E   , B���L B���\� C���\� C���L B���L      E   , E���L E���\� F���\� F���L E���L      E   , Hk��L Hk��\� I���\� I���L Hk��L      E   , KO��L KO��\� Lg��\� Lg��L KO��L      E   , N3��L N3��\� OK��\� OK��L N3��L      E   , Q��L Q��\� R/��\� R/��L Q��L      E   , S���L S���\� U��\� U��L S���L      E   , V���L V���\� W���\� W���L V���L      E   , Y���L Y���\� Z���\� Z���L Y���L      E   , \���L \���\� ]���\� ]���L \���L      E   , _���L _���\� `���\� `���L _���L      E   , bo��L bo��\� c���\� c���L bo��L      E   , eS��L eS��\� fk��\� fk��L eS��L      E   , h7��L h7��\� iO��\� iO��L h7��L      E   , k��L k��\� l3��\� l3��L k��L      E   , G��bg G��s3 _��s3 _��bg G��bg      E   , ����bg ����s3 ����s3 ����bg ����bg      E   , ����bg ����s3 ����s3 ����bg ����bg      E   , �w��bg �w��s3 ����s3 ����bg �w��bg      E   , �[��bg �[��s3 �s��s3 �s��bg �[��bg      E   , �?��bg �?��s3 �W��s3 �W��bg �?��bg      E   , �#��bg �#��s3 �;��s3 �;��bg �#��bg      E   , ���bg ���s3 ���s3 ���bg ���bg      E   , ����bg ����s3 ���s3 ���bg ����bg      E   , ����bg ����s3 ����s3 ����bg ����bg      E   , ����bg ����s3 ����s3 ����bg ����bg      E   , ����bg ����s3 ����s3 ����bg ����bg      E   , �{��bg �{��s3 ����s3 ����bg �{��bg      E   , �_��bg �_��s3 �w��s3 �w��bg �_��bg      E   , �C��bg �C��s3 �[��s3 �[��bg �C��bg      E   , �'��bg �'��s3 �?��s3 �?��bg �'��bg      E   , ���bg ���s3 �#��s3 �#��bg ���bg      E   , ����bg ����s3 ���s3 ���bg ����bg      E   , ����bg ����s3 ����s3 ����bg ����bg      E   , ķ��bg ķ��s3 ����s3 ����bg ķ��bg      E   , Ǜ��bg Ǜ��s3 ȳ��s3 ȳ��bg Ǜ��bg      E   , ���bg ���s3 ˗��s3 ˗��bg ���bg      E   , �c��bg �c��s3 �{��s3 �{��bg �c��bg      E   , p���bg p���s3 q���s3 q���bg p���bg      E   , s���bg s���s3 t���s3 t���bg s���bg      E   , v���bg v���s3 w���s3 w���bg v���bg      E   , y���bg y���s3 z���s3 z���bg y���bg      E   , |s��bg |s��s3 }���s3 }���bg |s��bg      E   , W��bg W��s3 �o��s3 �o��bg W��bg      E   , �;��bg �;��s3 �S��s3 �S��bg �;��bg      E   , ���bg ���s3 �7��s3 �7��bg ���bg      E   , ���bg ���s3 ���s3 ���bg ���bg      E   , ����bg ����s3 ����s3 ����bg ����bg      E   , ����bg ����s3 ����s3 ����bg ����bg      E   , p���L p���\� q���\� q���L p���L      E   , s���L s���\� t���\� t���L s���L      E   , v���L v���\� w���\� w���L v���L      E   , y���L y���\� z���\� z���L y���L      E   , |s��L |s��\� }���\� }���L |s��L      E   , W��L W��\� �o��\� �o��L W��L      E   , �;��L �;��\� �S��\� �S��L �;��L      E   , ���L ���\� �7��\� �7��L ���L      E   , ���L ���\� ���\� ���L ���L      E   , ����L ����\� ����\� ����L ����L      E   , ����L ����\� ����\� ����L ����L      E   , ����L ����\� ����\� ����L ����L      E   , ����L ����\� ����\� ����L ����L      E   , �w��L �w��\� ����\� ����L �w��L      E   , �[��L �[��\� �s��\� �s��L �[��L      E   , �?��L �?��\� �W��\� �W��L �?��L      E   , �#��L �#��\� �;��\� �;��L �#��L      E   , ���L ���\� ���\� ���L ���L      E   , ����L ����\� ���\� ���L ����L      E   , ����L ����\� ����\� ����L ����L      E   , ����L ����\� ����\� ����L ����L      E   , ����L ����\� ����\� ����L ����L      E   , �{��L �{��\� ����\� ����L �{��L      E   , �_��L �_��\� �w��\� �w��L �_��L      E   , �C��L �C��\� �[��\� �[��L �C��L      E   , �'��L �'��\� �?��\� �?��L �'��L      E   , ���L ���\� �#��\� �#��L ���L      E   , ����L ����\� ���\� ���L ����L      E   , ����L ����\� ����\� ����L ����L      E   , ķ��L ķ��\� ����\� ����L ķ��L      E   , Ǜ��L Ǜ��\� ȳ��\� ȳ��L Ǜ��L      E   , ���L ���\� ˗��\� ˗��L ���L      E   , �c��L �c��\� �{��\� �{��L �c��L      E   , ����Y� ����j� ����j� ����Y� ����Y�      E   , �,��Y� �,��j� �D��j� �D��Y� �,��Y�      E   , ڦ��Y� ڦ��jZ ۾��jZ ۾��Y� ڦ��Y�      F   ,  _�����  _�����  �����  �����  _�����      F   , ��b� ��s ���s ���b� ��b�      F   , ��L ��\� ���\� ���L ��L      F   , yD  4 yD  4+ z�  4+ z�  4 yD  4      F   , }�  4 }�  4+ \  4+ \  4 }�  4      F   , �  4 �  4+ ��  4+ ��  4 �  4      F   , ��  4 ��  4+ �/  4+ �/  4 ��  4      F   , �O  4 �O  4+ ��  4+ ��  4 �O  4      F   , ��  4 ��  4+ �g  4+ �g  4 ��  4      F   , ��  4 ��  4+ �  4+ �  4 ��  4      F   , �#  4 �#  4+ ��  4+ ��  4 �#  4      F   , ��  4 ��  4+ �;  4+ �;  4 ��  4      F   , �[  4 �[  4+ ��  4+ ��  4 �[  4      F   , ��  4 ��  4+ �s  4+ �s  4 ��  4      F   , ��  4 ��  4+ �  4+ �  4 ��  4      F   , �/  4 �/  4+ ƫ  4+ ƫ  4 �/  4      F   , ��  4 ��  4+ �G  4+ �G  4 ��  4      F   , �g  4 �g  4+ ��  4+ ��  4 �g  4      F   , y0  )" y0  4 z�  4 z�  )" y0  )"      F   , }�  )" }�  4 p  4 p  )" }�  )"      F   , �  )" �  4 ��  4 ��  )" �  )"      F   , ��  )" ��  4 �C  4 �C  )" ��  )"      F   , �;  )" �;  4 ��  4 ��  )" �;  )"      F   , ��  )" ��  4 �{  4 �{  )" ��  )"      F   , �s  )" �s  4 �  4 �  )" �s  )"      F   , �  )" �  4 ��  4 ��  )" �  )"      F   , ��  )" ��  4 �O  4 �O  )" ��  )"      F   , �G  )" �G  4 ��  4 ��  )" �G  )"      F   , ��  )" ��  4 ��  4 ��  )" ��  )"      F   , �  )" �  4 �#  4 �#  )" �  )"      F   , �  )" �  4 ƿ  4 ƿ  )" �  )"      F   , ɷ  )" ɷ  4 �[  4 �[  )" ɷ  )"      F   , �S  )" �S  4 ��  4 ��  )" �S  )"      F   , yD  )	 yD  )" z�  )" z�  )	 yD  )	      F   , }�  )	 }�  )" \  )" \  )	 }�  )	      F   , �  )	 �  )" ��  )" ��  )	 �  )	      F   , ��  )	 ��  )" �/  )" �/  )	 ��  )	      F   , �O  )	 �O  )" ��  )" ��  )	 �O  )	      F   , ��  )	 ��  )" �g  )" �g  )	 ��  )	      F   , ��  )	 ��  )" �  )" �  )	 ��  )	      F   , �#  )	 �#  )" ��  )" ��  )	 �#  )	      F   , ��  )	 ��  )" �;  )" �;  )	 ��  )	      F   , �[  )	 �[  )" ��  )" ��  )	 �[  )	      F   , ��  )	 ��  )" �s  )" �s  )	 ��  )	      F   , ��  )	 ��  )" �  )" �  )	 ��  )	      F   , �/  )	 �/  )" ƫ  )" ƫ  )	 �/  )	      F   , ��  )	 ��  )" �G  )" �G  )	 ��  )	      F   , �g  )	 �g  )" ��  )" ��  )	 �g  )	      F   , yD  #� yD  #� z�  #� z�  #� yD  #�      F   , }�  #� }�  #� \  #� \  #� }�  #�      F   , �  #� �  #� ��  #� ��  #� �  #�      F   , ��  #� ��  #� �/  #� �/  #� ��  #�      F   , �O  #� �O  #� ��  #� ��  #� �O  #�      F   , ��  #� ��  #� �g  #� �g  #� ��  #�      F   , ��  #� ��  #� �  #� �  #� ��  #�      F   , �#  #� �#  #� ��  #� ��  #� �#  #�      F   , ��  #� ��  #� �;  #� �;  #� ��  #�      F   , �[  #� �[  #� ��  #� ��  #� �[  #�      F   , ��  #� ��  #� �s  #� �s  #� ��  #�      F   , ��  #� ��  #� �  #� �  #� ��  #�      F   , �/  #� �/  #� ƫ  #� ƫ  #� �/  #�      F   , ��  #� ��  #� �G  #� �G  #� ��  #�      F   , �g  #� �g  #� ��  #� ��  #� �g  #�      F   , y0  � y0  #� z�  #� z�  � y0  �      F   , }�  � }�  #� p  #� p  � }�  �      F   , �  � �  #� ��  #� ��  � �  �      F   , ��  � ��  #� �C  #� �C  � ��  �      F   , �;  � �;  #� ��  #� ��  � �;  �      F   , ��  � ��  #� �{  #� �{  � ��  �      F   , �s  � �s  #� �  #� �  � �s  �      F   , �  � �  #� ��  #� ��  � �  �      F   , ��  � ��  #� �O  #� �O  � ��  �      F   , �G  � �G  #� ��  #� ��  � �G  �      F   , ��  � ��  #� ��  #� ��  � ��  �      F   , �  � �  #� �#  #� �#  � �  �      F   , �  � �  #� ƿ  #� ƿ  � �  �      F   , ɷ  � ɷ  #� �[  #� �[  � ɷ  �      F   , �S  � �S  #� ��  #� ��  � �S  �      F   , yD  � yD  � z�  � z�  � yD  �      F   , }�  � }�  � \  � \  � }�  �      F   , �  � �  � ��  � ��  � �  �      F   , ��  � ��  � �/  � �/  � ��  �      F   , �O  � �O  � ��  � ��  � �O  �      F   , ��  � ��  � �g  � �g  � ��  �      F   , ��  � ��  � �  � �  � ��  �      F   , �#  � �#  � ��  � ��  � �#  �      F   , ��  � ��  � �;  � �;  � ��  �      F   , �[  � �[  � ��  � ��  � �[  �      F   , ��  � ��  � �s  � �s  � ��  �      F   , ��  � ��  � �  � �  � ��  �      F   , �/  � �/  � ƫ  � ƫ  � �/  �      F   , ��  � ��  � �G  � �G  � ��  �      F   , �g  � �g  � ��  � ��  � �g  �      F   , F�  #� F�  #� H  #� H  #� F�  #�      F   , F�  4 F�  4+ H  4+ H  4 F�  4      F   , F|  � F|  #� H   #� H   � F|  �      F   , F�  )	 F�  )" H  )" H  )	 F�  )	      F   , F�  � F�  � H  � H  � F�  �      F   , F|  )" F|  4 H   4 H   )" F|  )"      F   , Td  #� Td  #� U�  #� U�  #� Td  #�      F   , Y   #� Y   #� Z|  #� Z|  #� Y   #�      F   , ]�  #� ]�  #� _  #� _  #� ]�  #�      F   , b8  #� b8  #� c�  #� c�  #� b8  #�      F   , f�  #� f�  #� hP  #� hP  #� f�  #�      F   , kp  #� kp  #� l�  #� l�  #� kp  #�      F   , p  #� p  #� q�  #� q�  #� p  #�      F   , t�  #� t�  #� v$  #� v$  #� t�  #�      F   , t�  )" t�  4 v8  4 v8  )" t�  )"      F   , k\  )" k\  4 m   4 m   )" k\  )"      F   , K,  4 K,  4+ L�  4+ L�  4 K,  4      F   , O�  4 O�  4+ QD  4+ QD  4 O�  4      F   , Td  4 Td  4+ U�  4+ U�  4 Td  4      F   , Y   4 Y   4+ Z|  4+ Z|  4 Y   4      F   , ]�  4 ]�  4+ _  4+ _  4 ]�  4      F   , b8  4 b8  4+ c�  4+ c�  4 b8  4      F   , f�  4 f�  4+ hP  4+ hP  4 f�  4      F   , kp  4 kp  4+ l�  4+ l�  4 kp  4      F   , p  4 p  4+ q�  4+ q�  4 p  4      F   , t�  4 t�  4+ v$  4+ v$  4 t�  4      F   , o�  )" o�  4 q�  4 q�  )" o�  )"      F   , K  � K  #� L�  #� L�  � K  �      F   , O�  � O�  #� QX  #� QX  � O�  �      F   , TP  � TP  #� U�  #� U�  � TP  �      F   , X�  � X�  #� Z�  #� Z�  � X�  �      F   , ]�  � ]�  #� _,  #� _,  � ]�  �      F   , b$  � b$  #� c�  #� c�  � b$  �      F   , f�  � f�  #� hd  #� hd  � f�  �      F   , k\  � k\  #� m   #� m   � k\  �      F   , o�  � o�  #� q�  #� q�  � o�  �      F   , t�  � t�  #� v8  #� v8  � t�  �      F   , f�  )" f�  4 hd  4 hd  )" f�  )"      F   , K,  )	 K,  )" L�  )" L�  )	 K,  )	      F   , O�  )	 O�  )" QD  )" QD  )	 O�  )	      F   , Td  )	 Td  )" U�  )" U�  )	 Td  )	      F   , Y   )	 Y   )" Z|  )" Z|  )	 Y   )	      F   , ]�  )	 ]�  )" _  )" _  )	 ]�  )	      F   , b8  )	 b8  )" c�  )" c�  )	 b8  )	      F   , f�  )	 f�  )" hP  )" hP  )	 f�  )	      F   , K,  #� K,  #� L�  #� L�  #� K,  #�      F   , K,  � K,  � L�  � L�  � K,  �      F   , O�  � O�  � QD  � QD  � O�  �      F   , Td  � Td  � U�  � U�  � Td  �      F   , Y   � Y   � Z|  � Z|  � Y   �      F   , ]�  � ]�  � _  � _  � ]�  �      F   , b8  � b8  � c�  � c�  � b8  �      F   , f�  � f�  � hP  � hP  � f�  �      F   , kp  � kp  � l�  � l�  � kp  �      F   , p  � p  � q�  � q�  � p  �      F   , t�  � t�  � v$  � v$  � t�  �      F   , kp  )	 kp  )" l�  )" l�  )	 kp  )	      F   , p  )	 p  )" q�  )" q�  )	 p  )	      F   , t�  )	 t�  )" v$  )" v$  )	 t�  )	      F   , O�  #� O�  #� QD  #� QD  #� O�  #�      F   , K  )" K  4 L�  4 L�  )" K  )"      F   , O�  )" O�  4 QX  4 QX  )" O�  )"      F   , TP  )" TP  4 U�  4 U�  )" TP  )"      F   , X�  )" X�  4 Z�  4 Z�  )" X�  )"      F   , ]�  )" ]�  4 _,  4 _,  )" ]�  )"      F   , b$  )" b$  4 c�  4 c�  )" b$  )"      F   , (�  4 (�  4+ *9  4+ *9  4 (�  4      F   , M  � M  � �  � �  � M  �      F   , �  � �  � e  � e  � �  �      F   , �  � �  � !  � !  � �  �      F   , $!  � $!  � %�  � %�  � $!  �      F   , (�  � (�  � *9  � *9  � (�  �      F   , -Y  � -Y  � .�  � .�  � -Y  �      F   , -Y  4 -Y  4+ .�  4+ .�  4 -Y  4      F   , M  #� M  #� �  #� �  #� M  #�      F   , �  #� �  #� e  #� e  #� �  #�      F   , �  #� �  #� !  #� !  #� �  #�      F   , $!  4 $!  4+ %�  4+ %�  4 $!  4      F   , 9  � 9  #� �  #� �  � 9  �      F   , �  � �  #� y  #� y  � �  �      F   , 9  )" 9  4 �  4 �  )" 9  )"      F   , M  )	 M  )" �  )" �  )	 M  )	      F   , �  )	 �  )" e  )" e  )	 �  )	      F   , �  )	 �  )" !  )" !  )	 �  )	      F   , $!  )	 $!  )" %�  )" %�  )	 $!  )	      F   , (�  )	 (�  )" *9  )" *9  )	 (�  )	      F   , -Y  )	 -Y  )" .�  )" .�  )	 -Y  )	      F   , �  )" �  4 y  4 y  )" �  )"      F   , q  )" q  4 !  4 !  )" q  )"      F   , $  )" $  4 %�  4 %�  )" $  )"      F   , (�  )" (�  4 *M  4 *M  )" (�  )"      F   , -E  )" -E  4 .�  4 .�  )" -E  )"      F   , q  � q  #� !  #� !  � q  �      F   , $  � $  #� %�  #� %�  � $  �      F   , (�  � (�  #� *M  #� *M  � (�  �      F   , -E  � -E  #� .�  #� .�  � -E  �      F   , $!  #� $!  #� %�  #� %�  #� $!  #�      F   , (�  #� (�  #� *9  #� *9  #� (�  #�      F   , -Y  #� -Y  #� .�  #� .�  #� -Y  #�      F   , M  4 M  4+ �  4+ �  4 M  4      F   , �  4 �  4+ e  4+ e  4 �  4      F   , �  4 �  4+ !  4+ !  4 �  4      F   ,  �	  �  �	  �  ��  �  ��  �  �	  �      F   ,  ��  �  ��  �  �!  �  �!  �  ��  �      F   ,  �A  �  �A  �  �  �  �  �  �A  �      F   , �  � �  � Y  � Y  � �  �      F   , y  � y  � 	�  � 	�  � y  �      F   ,   �   � �  � �  �   �      F   , �  � �  � -  � -  � �  �      F   , e  � e  #� 
	  #� 
	  � e  �      F   ,   �   #� �  #� �  �   �      F   , �  � �  #� A  #� A  � �  �      F   ,  ��  )	  ��  )"  �!  )"  �!  )	  ��  )	      F   ,  �A  )	  �A  )"  �  )"  �  )	  �A  )	      F   , �  )	 �  )" Y  )" Y  )	 �  )	      F   , y  )	 y  )" 	�  )" 	�  )	 y  )	      F   ,   )	   )" �  )" �  )	   )	      F   , �  )	 �  )" -  )" -  )	 �  )	      F   ,  ��  4  ��  4+  �!  4+  �!  4  ��  4      F   ,  �A  4  �A  4+  �  4+  �  4  �A  4      F   , �  4 �  4+ Y  4+ Y  4 �  4      F   ,  ��  )"  ��  4  ��  4  ��  )"  ��  )"      F   ,  ��  )"  ��  4  �5  4  �5  )"  ��  )"      F   ,  �-  )"  �-  4  �  4  �  )"  �-  )"      F   , �  )" �  4 m  4 m  )" �  )"      F   , e  )" e  4 
	  4 
	  )" e  )"      F   ,   )"   4 �  4 �  )"   )"      F   , �  )" �  4 A  4 A  )" �  )"      F   , y  4 y  4+ 	�  4+ 	�  4 y  4      F   ,  �	  #�  �	  #�  ��  #�  ��  #�  �	  #�      F   ,  ��  #�  ��  #�  �!  #�  �!  #�  ��  #�      F   ,  �A  #�  �A  #�  �  #�  �  #�  �A  #�      F   , �  #� �  #� Y  #� Y  #� �  #�      F   , y  #� y  #� 	�  #� 	�  #� y  #�      F   ,   #�   #� �  #� �  #�   #�      F   , �  #� �  #� -  #� -  #� �  #�      F   ,   4   4+ �  4+ �  4   4      F   , �  4 �  4+ -  4+ -  4 �  4      F   ,  �	  4  �	  4+  ��  4+  ��  4  �	  4      F   ,  �	  )	  �	  )"  ��  )"  ��  )	  �	  )	      F   ,  ��  �  ��  #�  ��  #�  ��  �  ��  �      F   ,  _�  �  _�  �  ��  �  ��  �  _�  �      F   ,  ��  �  ��  �  ��  �  ��  �  ��  �      F   ,  �G  �  �G  �  ��  �  ��  �  �G  �      F   ,  ��  �  ��  �  �-  �  �-  �  ��  �      F   ,  �X  �  �X  �  Ɲ  �  Ɲ  �  �X  �      F   ,  _����}  _�  �  ��  �  �����}  _����}      F   ,  _�����  _�����  ������  ������  _�����      F   ,  ����ޕ  ����ޚ  ����ޚ  ����ޕ  ����ޕ      F   ,  �G��ޕ  �G��ޚ  ����ޚ  ����ޕ  �G��ޕ      F   ,  ����ޕ  ����ޚ  �-��ޚ  �-��ޕ  ����ޕ      F   ,  �X��ޕ  �X��ޚ  Ɲ��ޚ  Ɲ��ޕ  �X��ޕ      F   ,  _����s  _���ޕ  ����ޕ  �����s  _����s      F   ,  ��  �  ��  #�  �5  #�  �5  �  ��  �      F   ,  �-  �  �-  #�  �  #�  �  �  �-  �      F   , �  � �  #� m  #� m  � �  �      F   ,  _����i  _�����  �����  ����i  _����i      F   ,  _�����  _�����  �����  �����  _�����      F   ,  _����_  _�����  �����  ����_  _����_      F   ,  ������  ������  �����  �����  ������      F   ,  i-����  i-����  jr����  jr����  i-����      F   ,  {�����  {�����  |�����  |�����  {�����      F   ,  �>����  �>����  ������  ������  �>����      F   ,  ������  ������  �����  �����  ������      F   ,  �>����  �>����  ������  ������  �>����      F   ,  i-����  i-����  jr����  jr����  i-����      F   ,  {�����  {�����  |�����  |�����  {�����      F   ,  t���r�  t���s  v%��s  v%��r�  t���r�      F   ,  yE��r�  yE��s  z���s  z���r�  yE��r�      F   ,  }���r�  }���s  ]��s  ]��r�  }���r�      F   ,  �}��r�  �}��s  ����s  ����r�  �}��r�      F   ,  ���r�  ���s  ����s  ����r�  ���r�      F   ,  ����r�  ����s  �1��s  �1��r�  ����r�      F   ,  �Q��r�  �Q��s  ����s  ����r�  �Q��r�      F   ,  ����r�  ����s  �i��s  �i��r�  ����r�      F   ,  ����r�  ����s  �+��s  �+��r�  ����r�      F   ,  �K��r�  �K��s  ����s  ����r�  �K��r�      F   ,  ����r�  ����s  �c��s  �c��r�  ����r�      F   ,  ����r�  ����s  ����s  ����r�  ����r�      F   ,  ���r�  ���s  ����s  ����r�  ���r�      F   ,  NR��p  NR��p1  O���p1  O���p  NR��p      F   ,  t���g�  t���r�  v9��r�  v9��g�  t���g�      F   ,  y1��g�  y1��r�  z���r�  z���g�  y1��g�      F   ,  }���g�  }���r�  q��r�  q��g�  }���g�      F   ,  �i��g�  �i��r�  ���r�  ���g�  �i��g�      F   ,  ���g�  ���r�  ����r�  ����g�  ���g�      F   ,  ����g�  ����r�  �E��r�  �E��g�  ����g�      F   ,  �=��g�  �=��r�  ����r�  ����g�  �=��g�      F   ,  ����g�  ����r�  �}��r�  �}��g�  ����g�      F   ,  ����g�  ����r�  �?��r�  �?��g�  ����g�      F   ,  �7��g�  �7��r�  ����r�  ����g�  �7��g�      F   ,  ����g�  ����r�  �w��r�  �w��g�  ����g�      F   ,  �o��g�  �o��r�  ���r�  ���g�  �o��g�      F   ,  ���g�  ���r�  ����r�  ����g�  ���g�      F   ,  t���g�  t���g�  v%��g�  v%��g�  t���g�      F   ,  yE��g�  yE��g�  z���g�  z���g�  yE��g�      F   ,  }���g�  }���g�  ]��g�  ]��g�  }���g�      F   ,  �}��g�  �}��g�  ����g�  ����g�  �}��g�      F   ,  ���g�  ���g�  ����g�  ����g�  ���g�      F   ,  ����g�  ����g�  �1��g�  �1��g�  ����g�      F   ,  �Q��g�  �Q��g�  ����g�  ����g�  �Q��g�      F   ,  ����g�  ����g�  �i��g�  �i��g�  ����g�      F   ,  ����g�  ����g�  �+��g�  �+��g�  ����g�      F   ,  �K��g�  �K��g�  ����g�  ����g�  �K��g�      F   ,  ����g�  ����g�  �c��g�  �c��g�  ����g�      F   ,  ����g�  ����g�  ����g�  ����g�  ����g�      F   ,  ���g�  ���g�  ����g�  ����g�  ���g�      F   ,  t���b�  t���c  v%��c  v%��b�  t���b�      F   ,  yE��b�  yE��c  z���c  z���b�  yE��b�      F   ,  }���b�  }���c  ]��c  ]��b�  }���b�      F   ,  �}��b�  �}��c  ����c  ����b�  �}��b�      F   ,  ���b�  ���c  ����c  ����b�  ���b�      F   ,  ����b�  ����c  �1��c  �1��b�  ����b�      F   ,  �Q��b�  �Q��c  ����c  ����b�  �Q��b�      F   ,  ����b�  ����c  �i��c  �i��b�  ����b�      F   ,  ����b�  ����c  �+��c  �+��b�  ����b�      F   ,  �K��b�  �K��c  ����c  ����b�  �K��b�      F   ,  ����b�  ����c  �c��c  �c��b�  ����b�      F   ,  ����b�  ����c  ����c  ����b�  ����b�      F   ,  ���b�  ���c  ����c  ����b�  ���b�      F   ,  t���X  t���b�  v9��b�  v9��X  t���X      F   ,  y1��X  y1��b�  z���b�  z���X  y1��X      F   ,  }���X  }���b�  q��b�  q��X  }���X      F   ,  �i��X  �i��b�  ���b�  ���X  �i��X      F   ,  ���X  ���b�  ����b�  ����X  ���X      F   ,  ����X  ����b�  �E��b�  �E��X  ����X      F   ,  �=��X  �=��b�  ����b�  ����X  �=��X      F   ,  ����X  ����b�  �}��b�  �}��X  ����X      F   ,  ����X  ����b�  �?��b�  �?��X  ����X      F   ,  �7��X  �7��b�  ����b�  ����X  �7��X      F   ,  ����X  ����b�  �w��b�  �w��X  ����X      F   ,  �o��X  �o��b�  ���b�  ���X  �o��X      F   ,  ���X  ���b�  ����b�  ����X  ���X      F   ,  t���W�  t���X  v%��X  v%��W�  t���W�      F   ,  yE��W�  yE��X  z���X  z���W�  yE��W�      F   ,  }���W�  }���X  ]��X  ]��W�  }���W�      F   ,  �}��W�  �}��X  ����X  ����W�  �}��W�      F   ,  ���W�  ���X  ����X  ����W�  ���W�      F   ,  ����W�  ����X  �1��X  �1��W�  ����W�      F   ,  �Q��W�  �Q��X  ����X  ����W�  �Q��W�      F   ,  ����W�  ����X  �i��X  �i��W�  ����W�      F   ,  ����W�  ����X  �+��X  �+��W�  ����W�      F   ,  �K��W�  �K��X  ����X  ����W�  �K��W�      F   ,  ����W�  ����X  �c��X  �c��W�  ����W�      F   ,  ����W�  ����X  ����X  ����W�  ����W�      F   ,  ���W�  ���X  ����X  ����W�  ���W�      F   ,  NR��{!  NR��{:  O���{:  O���{!  NR��{!      F   ,  N>��p1  N>��{!  O���{!  O���p1  N>��p1      F   ,  ����r�  ����s  �o��s  �o��r�  ����r�      F   ,  ����g�  ����g�  �7��g�  �7��g�  ����g�      F   ,  �W��g�  �W��g�  ����g�  ����g�  �W��g�      F   ,  ����g�  ����g�  �o��g�  �o��g�  ����g�      F   ,  ����r�  ����s  �7��s  �7��r�  ����r�      F   ,  �W��r�  �W��s  ����s  ����r�  �W��r�      F   ,  ����g�  ����r�  �K��r�  �K��g�  ����g�      F   ,  �C��g�  �C��r�  ����r�  ����g�  �C��g�      F   ,  ����b�  ����c  �7��c  �7��b�  ����b�      F   ,  �W��b�  �W��c  ����c  ����b�  �W��b�      F   ,  ����b�  ����c  �o��c  �o��b�  ����b�      F   ,  ����g�  ����r�  ����r�  ����g�  ����g�      F   ,  ����X  ����b�  �K��b�  �K��X  ����X      F   ,  ����W�  ����X  �7��X  �7��W�  ����W�      F   ,  �W��W�  �W��X  ����X  ����W�  �W��W�      F   ,  ����W�  ����X  �o��X  �o��W�  ����W�      F   ,  �e��L  �e��s  ����s  ����L  �e��L      F   ,  �5��b�  �5��s  ����s  ����b�  �5��b�      F   ,  �5��L  �5��\�  ����\�  ����L  �5��L      F   ,  �-��L  �-��s  ����s  ����L  �-��L      F   ,  ����b�  ����s  ����s  ����b�  ����b�      F   ,  ����L  ����\�  ����\�  ����L  ����L      F   ,  ����L  ����s q��s q��L  ����L      F   , ���b� ���s i��s i��b� ���b�      F   , ���L ���\� i��\� i��L ���L      F   , ���L ���s 9��s 9��L ���L      F   , ���b� ���s 
1��s 
1��b� ���b�      F   , ���L ���\� 
1��\� 
1��L ���L      F   , ���L ���s ��s ��L ���L      F   , U��b� U��s ���s ���b� U��b�      F   , U��L U��\� ���\� ���L U��L      F   , M��L M��s ���s ���L M��L      F   ,  �C��X  �C��b�  ����b�  ����X  �C��X      F   ,  ����X  ����b�  ����b�  ����X  ����X      F   , ��L ��s ���s ���L ��L      F   , ���b� ���s ���s ���b� ���b�      F   , ���L ���\� ���\� ���L ���L      F   , ���L ���s Y��s Y��L ���L      F   , ���b� ���s !Q��s !Q��b� ���b�      F   , ���L ���\� !Q��\� !Q��L ���L      F   , "���L "���s $!��s $!��L "���L      F   , %u��b� %u��s '��s '��b� %u��b�      F   , %u��L %u��\� '��\� '��L %u��L      F   , (m��L (m��s )���s )���L (m��L      F   , +=��b� +=��s ,���s ,���b� +=��b�      F   , +=��L +=��\� ,���\� ,���L +=��L      F   , .5��L .5��s /���s /���L .5��L      F   , 1��b� 1��s 2���s 2���b� 1��b�      F   , 1��L 1��\� 2���\� 2���L 1��L      F   , 3���L 3���s 5y��s 5y��L 3���L      F   , 6���b� 6���s 8q��s 8q��b� 6���b�      F   , 6���L 6���\� 8q��\� 8q��L 6���L      F   , 9���L 9���s ;A��s ;A��L 9���L      F   , <���b� <���s >9��s >9��b� <���b�      F   , <���L <���\� >9��\� >9��L <���L      F   , ?���L ?���s A	��s A	��L ?���L      F   , B]��b� B]��s D��s D��b� B]��b�      F   , B]��L B]��\� D��\� D��L B]��L      F   , EU��L EU��s F���s F���L EU��L      F   , H%��b� H%��s I���s I���b� H%��b�      F   , H%��L H%��\� I���\� I���L H%��L      F   , K��L K��s L���s L���L K��L      F   , M���b� M���s O���s O���b� M���b�      F   , M���L M���\� O���\� O���L M���L      F   , P���L P���s Ra��s Ra��L P���L      F   , S���b� S���s UY��s UY��b� S���b�      F   , S���L S���\� UY��\� UY��L S���L      F   , V���L V���s X)��s X)��L V���L      F   , Y}��b� Y}��s [!��s [!��b� Y}��b�      F   , Y}��L Y}��\� [!��\� [!��L Y}��L      F   , \u��L \u��s ]���s ]���L \u��L      F   , _E��b� _E��s `���s `���b� _E��b�      F   , _E��L _E��\� `���\� `���L _E��L      F   , b=��L b=��s c���s c���L b=��L      F   , e��b� e��s f���s f���b� e��b�      F   , e��L e��\� f���\� f���L e��L      F   , h��L h��s i���s i���L h��L      F   , j���b� j���s ly��s ly��b� j���b�      F   , j���L j���\� ly��\� ly��L j���L      F   , m���L m���s oI��s oI��L m���L      F   , p���b� p���s rA��s rA��b� p���b�      F   , p���L p���\� rA��\� rA��L p���L      F   , s���L s���s u��s u��L s���L      F   , ve��b� ve��s x	��s x	��b� ve��b�      F   , ve��L ve��\� x	��\� x	��L ve��L      F   , y]��L y]��s z���s z���L y]��L      F   , |-��b� |-��s }���s }���b� |-��b�      F   , |-��L |-��\� }���\� }���L |-��L      F   , %��L %��s ����s ����L %��L      F   , ����b� ����s ����s ����b� ����b�      F   , ����L ����\� ����\� ����L ����L      F   , ����L ����s �i��s �i��L ����L      F   , ����b� ����s �a��s �a��b� ����b�      F   , ����L ����\� �a��\� �a��L ����L      F   , ����L ����s �1��s �1��L ����L      F   , ����b� ����s �)��s �)��b� ����b�      F   , ����L ����\� �)��\� �)��L ����L      F   , �}��L �}��s ����s ����L �}��L      F   , �M��b� �M��s ����s ����b� �M��b�      F   , �M��L �M��\� ����\� ����L �M��L      F   , �E��L �E��s ����s ����L �E��L      F   , ���b� ���s ����s ����b� ���b�      F   , ���L ���\� ����\� ����L ���L      F   , ���L ���s ����s ����L ���L      F   , ����b� ����s ����s ����b� ����b�      F   , ����L ����\� ����\� ����L ����L      F   , ����L ����s �Q��s �Q��L ����L      F   , ����b� ����s �I��s �I��b� ����b�      F   , ����L ����\� �I��\� �I��L ����L      F   , ����L ����s ���s ���L ����L      F   , �m��b� �m��s ���s ���b� �m��b�      F   , �m��L �m��\� ���\� ���L �m��L      F   , �e��L �e��s ����s ����L �e��L      F   , �5��b� �5��s ����s ����b� �5��b�      F   , �5��L �5��\� ����\� ����L �5��L      F   , �-��L �-��s ����s ����L �-��L      F   , ����b� ����s ����s ����b� ����b�      F   , ����L ����\� ����\� ����L ����L      F   , ����L ����s �q��s �q��L ����L      F   , ����b� ����s �i��s �i��b� ����b�      F   , ����L ����\� �i��\� �i��L ����L      F   , ����L ����s �9��s �9��L ����L      F   , ����b� ����s �1��s �1��b� ����b�      F   , ����L ����\� �1��\� �1��L ����L      F   , ą��L ą��s ���s ���L ą��L      F   , �U��b� �U��s ����s ����b� �U��b�      F   , �U��L �U��\� ����\� ����L �U��L      F   , �M��L �M��s ����s ����L �M��L      F   , ���b� ���s ����s ����b� ���b�      F   , ���L ���\� ����\� ����L ���L      F   , ����Y� ����j� �v��j� �v��Y� ����Y�      F   , �`��Y� �`��jA ���jA ���Y� �`��Y�      G   , -r  � -r  4 .�  4 .�  � -r  �      G   ,  s���r�  s����q  �����q  ����r�  s���r�      G   ,  ������  ������  ������  ������  ������      G   , ����T ����p ����p ����T ����T      G   , T}  # T}  4 U�  4 U�  # T}  #      G   , Y  # Y  4 Zc  4 Zc  # Y  #      G   , ]�  # ]�  4 ^�  4 ^�  # ]�  #      G   , bQ  # bQ  4 c�  4 c�  # bQ  #      G   , f�  # f�  4 h7  4 h7  # f�  #      G   , k�  # k�  4 l�  4 l�  # k�  #      G   , p%  # p%  4 qo  4 qo  # p%  #      G   , t�  # t�  4 v  4 v  # t�  #      G   , y]  # y]  4 z�  4 z�  # y]  #      G   , }�  # }�  4 C  4 C  # }�  #      G   , �0  # �0  4 �z  4 �z  # �0  #      G   , ��  # ��  4 �  4 �  # ��  #      G   , �h  # �h  4 ��  4 ��  # �h  #      G   , �  # �  4 �N  4 �N  # �  #      G   , ��  # ��  4 ��  4 ��  # ��  #      G   , �<  # �<  4 ��  4 ��  # �<  #      G   , ��  # ��  4 �"  4 �"  # ��  #      G   , �t  # �t  4 ��  4 ��  # �t  #      G   , �  # �  4 �Z  4 �Z  # �  #      G   , ��  # ��  4 ��  4 ��  # ��  #      G   , �H  # �H  4 ƒ  4 ƒ  # �H  #      G   , ��  # ��  4 �.  4 �.  # ��  #      G   , ΀  # ΀  4 ��  4 ��  # ΀  #      G   , �����p �����@ ����@ ����p �����p      G   , F�  # F�  4 G�  4 G�  # F�  #      G   , KE  # KE  4 L�  4 L�  # KE  #      G   , O�  # O�  4 Q+  4 Q+  # O�  #      G   , �  � �  4 	�  4 	�  � �  �      G   , .  � .  4 x  4 x  � .  �      G   , �  � �  4   4   � �  �      G   , f  � f  4 �  4 �  � f  �      G   ,   �   4 L  4 L  �   �      G   , �  � �  4  �  4  �  � �  �      G   , $:  � $:  4 %�  4 %�  � $:  �      G   , (�  � (�  4 *   4 *   � (�  �      G   ,  _�����  _�  �  �;  �  �;����  _�����      G   ,  �"  �  �"  4  �l  4  �l  �  �"  �      G   ,  s����q  s�����  ������  �����q  s����q      G   ,  ��  �  ��  4  �  4  �  �  ��  �      G   ,  �Z  �  �Z  4  �  4  �  �  �Z  �      G   , �  � �  4 @  4 @  � �  �      G   ,  Nk��p,  Nk��{&  O���{&  O���p,  Nk��p,      G   ,  ���r�  �����  �����  ���r�  ���r�      G   ,  s���X  s���r�  �P��r�  �P��X  s���X      G   ,  ����g�  ����r�  �V��r�  �V��g�  ����g�      G   ,  ����b�  ����g�  �V��g�  �V��b�  ����b�      G   ,  s���W�  s���X  v��X  v��W�  s���W�      G   ,  y^��W�  y^��X  z���X  z���W�  y^��W�      G   ,  }���W�  }���X  D��X  D��W�  }���W�      G   ,  ����W�  ����X  ����X  ����W�  ����W�      G   ,  �2��W�  �2��X  �|��X  �|��W�  �2��W�      G   ,  ����W�  ����X  ���X  ���W�  ����W�      G   ,  �j��W�  �j��X  ����X  ����W�  �j��W�      G   ,  ���W�  ���X  �P��X  �P��W�  ���W�      G   ,  ����X  ����b�  �V��b�  �V��X  ����X      G   ,  ����W�  ����X  ���X  ���W�  ����W�      G   ,  �d��W�  �d��X  ����X  ����W�  �d��W�      G   ,  � ��W�  � ��X  �J��X  �J��W�  � ��W�      G   ,  ����W�  ����X  ����X  ����W�  ����W�      G   ,  �8��W�  �8��X  ����X  ����W�  �8��W�      G   ,  ����W�  ����X  ���X  ���W�  ����W�      G   ,  �p��W�  �p��X  ����X  ����W�  �p��W�      G   ,  ���W�  ���X  �V��X  �V��W�  ���W�      G   ,  �I��L  �I���u  �����u  ����L  �I��L      G   ,  ���L  �����  ������  ����L  ���L      G   , ���L ����G U���G U��L ���L      G   , ���L ����u 
���u 
��L ���L      G   , i��L i���� ����� ���L i��L      G   , 1��L 1���G ����G ���L 1��L      G   , ���L ����u u���u u��L ���L      G   , ���L ����� !=���� !=��L ���L      G   , %���L %����G '���G '��L %���L      G   , +Q��L +Q���u ,����u ,���L +Q��L      G   , ������ �����T ����T ����� ������      G   , 1��L 1���u 2����u 2���L 1��L      G   , 6���L 6���� 8]��� 8]��L 6���L      G   , <���L <����a >%���a >%��L <���L      G   , Bq��L Bq���u C����u C���L Bq��L      G   , H9��L H9���� I����� I���L H9��L      G   , N��L N���G O}���G O}��L N��L      G   , S���L S����u UE���u UE��L S���L      G   , Y���L Y����� [���� [��L Y���L      G   , _Y��L _Y���G `����G `���L _Y��L      G   , e!��L e!���u f����u f���L e!��L      G   , j���L j����u le���u le��L j���L      G   , p���L p����� r-���� r-��L p���L      G   , vy��L vy���G w����G w���L vy��L      G   , |A��L |A���u }����u }���L |A��L      G   , �	��L �	��@ ����@ ����L �	��L      G   , ����L ������ �M���� �M��L ����L      G   , ����L �����u ����u ���L ����L      G   , �a��L �a���u �����u ����L �a��L      G   , �)��L �)���� ������ ����L �)��L      G   , ����L �����u �m���u �m��L ����L      G   , ����L �����u �5���u �5��L ����L      G   , ����L ������ ������ ����L ����L      G   , �I��L �I���G �����G ����L �I��L      G   , ���L ����u �����u ����L ���L      G   , ����L ������ �U���� �U��L ����L      G   , ����L �����G ����G ���L ����L      G   , �i��L �i���u �����u ����L �i��L      G   , �1��L �1���� έ���� έ��L �1��L      G   , ڍ��Y� ڍ��j ����j ����Y� ڍ��Y�      A   ,  ]����r  ]����*  ����*  ����r  ]����r      A   , r�  (� r�  4: sm  4: sm  (� r�  (�      A   , r�  � r�  #� sm  #� sm  � r�  �      A   , w_  (� w_  4: x	  4: x	  (� w_  (�      A   , y�  (� y�  4: zW  4: zW  (� y�  (�      A   , {�  (� {�  4: |�  4: |�  (� {�  (�      A   , ~I  (� ~I  4: ~�  4: ~�  (� ~I  (�      A   , �j  (� �j  4: �  4: �  (� �j  (�      A   , ��  (� ��  4: �b  4: �b  (� ��  (�      A   , �  (� �  4: ��  4: ��  (� �  (�      A   , �T  (� �T  4: ��  4: ��  (� �T  (�      A   , ��  (� ��  4: �L  4: �L  (� ��  (�      A   , ��  (� ��  4: ��  4: ��  (� ��  (�      A   , �>  (� �>  4: ��  4: ��  (� �>  (�      A   , ��  (� ��  4: �6  4: �6  (� ��  (�      A   , ��  (� ��  4: ��  4: ��  (� ��  (�      A   , �(  (� �(  4: ��  4: ��  (� �(  (�      A   , �v  (� �v  4: �   4: �   (� �v  (�      A   , ��  (� ��  4: �n  4: �n  (� ��  (�      A   , �  (� �  4: ��  4: ��  (� �  (�      A   , �`  (� �`  4: �
  4: �
  (� �`  (�      A   , ��  (� ��  4: �X  4: �X  (� ��  (�      A   , ��  (� ��  4: ��  4: ��  (� ��  (�      A   , �J  (� �J  4: ��  4: ��  (� �J  (�      A   , Ř  (� Ř  4: �B  4: �B  (� Ř  (�      A   , ��  (� ��  4: Ȑ  4: Ȑ  (� ��  (�      A   , �4  (� �4  4: ��  4: ��  (� �4  (�      A   , ̂  (� ̂  4: �,  4: �,  (� ̂  (�      A   , ��  (� ��  4: �z  4: �z  (� ��  (�      A   , u  (� u  4: u�  4: u�  (� u  (�      A   , u  � u  #� u�  #� u�  � u  �      A   , w_  � w_  #� x	  #� x	  � w_  �      A   , y�  � y�  #� zW  #� zW  � y�  �      A   , {�  � {�  #� |�  #� |�  � {�  �      A   , ~I  � ~I  #� ~�  #� ~�  � ~I  �      A   , �j  � �j  #� �  #� �  � �j  �      A   , ��  � ��  #� �b  #� �b  � ��  �      A   , �  � �  #� ��  #� ��  � �  �      A   , �T  � �T  #� ��  #� ��  � �T  �      A   , ��  � ��  #� �L  #� �L  � ��  �      A   , ��  � ��  #� ��  #� ��  � ��  �      A   , �>  � �>  #� ��  #� ��  � �>  �      A   , ��  � ��  #� �6  #� �6  � ��  �      A   , ��  � ��  #� ��  #� ��  � ��  �      A   , �(  � �(  #� ��  #� ��  � �(  �      A   , �v  � �v  #� �   #� �   � �v  �      A   , ��  � ��  #� �n  #� �n  � ��  �      A   , �  � �  #� ��  #� ��  � �  �      A   , �`  � �`  #� �
  #� �
  � �`  �      A   , ��  � ��  #� �X  #� �X  � ��  �      A   , ��  � ��  #� ��  #� ��  � ��  �      A   , �J  � �J  #� ��  #� ��  � �J  �      A   , Ř  � Ř  #� �B  #� �B  � Ř  �      A   , ��  � ��  #� Ȑ  #� Ȑ  � ��  �      A   , �4  � �4  #� ��  #� ��  � �4  �      A   , ̂  � ̂  #� �,  #� �,  � ̂  �      A   , ��  � ��  #� �z  #� �z  � ��  �      A   , R  � R  #� �  #� �  � R  �      A   , �  � �  #� J  #� J  � �  �      A   , �  � �  #�  �  #�  �  � �  �      A   , "<  � "<  #� "�  #� "�  � "<  �      A   , $�  � $�  #� %4  #� %4  � $�  �      A   , &�  � &�  #� '�  #� '�  � &�  �      A   , )&  � )&  #� )�  #� )�  � )&  �      A   , +t  � +t  #� ,  #� ,  � +t  �      A   , -�  � -�  #� .l  #� .l  � -�  �      A   , M�  � M�  #� N�  #� N�  � M�  �      A   , P1  � P1  #� P�  #� P�  � P1  �      A   , R  � R  #� S)  #� S)  � R  �      A   , T�  � T�  #� Uw  #� Uw  � T�  �      A   , W  � W  #� W�  #� W�  � W  �      A   , Yi  � Yi  #� Z  #� Z  � Yi  �      A   , [�  � [�  #� \a  #� \a  � [�  �      A   , ^  � ^  #� ^�  #� ^�  � ^  �      A   , `S  � `S  #� `�  #� `�  � `S  �      A   , b�  � b�  #� cK  #� cK  � b�  �      A   , d�  � d�  #� e�  #� e�  � d�  �      A   , g=  � g=  #� g�  #� g�  � g=  �      A   , i�  � i�  #� j5  #� j5  � i�  �      A   , k�  � k�  #� l�  #� l�  � k�  �      A   , n'  � n'  #� n�  #� n�  � n'  �      A   , pu  � pu  #� q  #� q  � pu  �      A   , �  (� �  4: J  4: J  (� �  (�      A   , �  (� �  4:  �  4:  �  (� �  (�      A   , "<  (� "<  4: "�  4: "�  (� "<  (�      A   , $�  (� $�  4: %4  4: %4  (� $�  (�      A   , &�  (� &�  4: '�  4: '�  (� &�  (�      A   , )&  (� )&  4: )�  4: )�  (� )&  (�      A   , +t  (� +t  4: ,  4: ,  (� +t  (�      A   , -�  (� -�  4: .l  4: .l  (� -�  (�      A   , M�  (� M�  4: N�  4: N�  (� M�  (�      A   , P1  (� P1  4: P�  4: P�  (� P1  (�      A   , R  (� R  4: S)  4: S)  (� R  (�      A   , T�  (� T�  4: Uw  4: Uw  (� T�  (�      A   , W  (� W  4: W�  4: W�  (� W  (�      A   , Yi  (� Yi  4: Z  4: Z  (� Yi  (�      A   , [�  (� [�  4: \a  4: \a  (� [�  (�      A   , ^  (� ^  4: ^�  4: ^�  (� ^  (�      A   , `S  (� `S  4: `�  4: `�  (� `S  (�      A   , b�  (� b�  4: cK  4: cK  (� b�  (�      A   , d�  (� d�  4: e�  4: e�  (� d�  (�      A   , g=  (� g=  4: g�  4: g�  (� g=  (�      A   , i�  (� i�  4: j5  4: j5  (� i�  (�      A   , k�  (� k�  4: l�  4: l�  (� k�  (�      A   , n'  (� n'  4: n�  4: n�  (� n'  (�      A   , pu  (� pu  4: q  4: q  (� pu  (�      A   ,   (�   4: �  4: �  (�   (�      A   , R  (� R  4: �  4: �  (� R  (�      A   , �  � �  #� `  #� `  � �  �      A   ,   �   #� �  #� �  �   �      A   , �  (� �  4: `  4: `  (� �  (�      A   ,  ��  �  ��  #�  T  #�  T  �  ��  �      A   , �  � �  #� �  #� �  � �  �      A   , F  � F  #� �  #� �  � F  �      A   , �  � �  #� >  #� >  � �  �      A   , �  � �  #� 	�  #� 	�  � �  �      A   , 0  � 0  #� �  #� �  � 0  �      A   , ~  � ~  #� (  #� (  � ~  �      A   , �  � �  #� v  #� v  � �  �      A   ,   �   #� �  #� �  �   �      A   , h  � h  #�   #�   � h  �      A   ,  �\  (�  �\  4:  �  4:  �  (�  �\  (�      A   ,  ��  (�  ��  4:  T  4:  T  (�  ��  (�      A   , �  (� �  4: �  4: �  (� �  (�      A   , F  (� F  4: �  4: �  (� F  (�      A   , �  (� �  4: >  4: >  (� �  (�      A   , �  (� �  4: 	�  4: 	�  (� �  (�      A   , 0  (� 0  4: �  4: �  (� 0  (�      A   , ~  (� ~  4: (  4: (  (� ~  (�      A   , �  (� �  4: v  4: v  (� �  (�      A   ,   (�   4: �  4: �  (�   (�      A   , h  (� h  4:   4:   (� h  (�      A   ,  ]�  �  ]�  >  �  >  �  �  ]�  �      A   ,  ]����2  ]�  �  �  �  ����2  ]����2      A   ,  ]����|  ]����4  ����4  ����|  ]����|      A   ,  ]����(  ]�����  �����  ����(  ]����(      A   ,  �\  �  �\  #�  �  #�  �  �  �\  �      A   ,  ]����  ]�����  �����  ����  ]����      A   ,  pb����  pb����  q����  q����  pb����      A   ,  r�����  r�����  sZ����  sZ����  r�����      A   ,  t�����  t�����  u�����  u�����  t�����      A   ,  wL����  wL����  w�����  w�����  wL����      A   ,  ������  ������  ������  ������  ������      A   ,  �8����  �8����  ������  ������  �8����      A   ,  ������  ������  �0����  �0����  ������      A   ,  ������  ������  �~����  �~����  ������      A   ,  �"����  �"����  ������  ������  �"����      A   ,  �p����  �p����  �����  �����  �p����      A   ,  ������  ������  �h����  �h����  ������      A   ,  �����  �����  ������  ������  �����      A   ,  �Z����  �Z����  �����  �����  �Z����      A   ,  Ũ����  Ũ����  �R����  �R����  Ũ����      A   ,  ������  ������  Ƞ����  Ƞ����  ������      A   ,  �D����  �D����  ������  ������  �D����      A   ,  pb���P  pb����  q����  q���P  pb���P      A   ,  r����P  r�����  sZ����  sZ���P  r����P      A   ,  t����P  t�����  u�����  u����P  t����P      A   ,  wL���P  wL����  w�����  w����P  wL���P      A   ,  �����P  ������  ������  �����P  �����P      A   ,  �8���P  �8����  ������  �����P  �8���P      A   ,  �����P  ������  �0����  �0���P  �����P      A   ,  �����P  ������  �~����  �~���P  �����P      A   ,  �"���P  �"����  ������  �����P  �"���P      A   ,  �p���P  �p����  �����  ����P  �p���P      A   ,  �����P  ������  �h����  �h���P  �����P      A   ,  ����P  �����  ������  �����P  ����P      A   ,  �Z���P  �Z����  �����  ����P  �Z���P      A   ,  Ũ���P  Ũ����  �R����  �R���P  Ũ���P      A   ,  �����P  ������  Ƞ����  Ƞ���P  �����P      A   ,  �D���P  �D����  ������  �����P  �D���P      A   ,  {���g�  {���s  |���s  |���g�  {���g�      A   ,  ~J��g�  ~J��s  ~���s  ~���g�  ~J��g�      A   ,  ����g�  ����s  �B��s  �B��g�  ����g�      A   ,  ����g�  ����s  ����s  ����g�  ����g�      A   ,  ����g�  ����s  �t��s  �t��g�  ����g�      A   ,  ���g�  ���s  ����s  ����g�  ���g�      A   ,  �f��g�  �f��s  ���s  ���g�  �f��g�      A   ,  ����g�  ����s  �^��s  �^��g�  ����g�      A   ,  ���g�  ���s  ����s  ����g�  ���g�      A   ,  �P��g�  �P��s  ����s  ����g�  �P��g�      A   ,  ����g�  ����s  �H��s  �H��g�  ����g�      A   ,  ����g�  ����s  ����s  ����g�  ����g�      A   ,  �:��g�  �:��s  ����s  ����g�  �:��g�      A   ,  ����g�  ����s  �2��s  �2��g�  ����g�      A   ,  ����g�  ����s  ����s  ����g�  ����g�      A   ,  �$��g�  �$��s  ����s  ����g�  �$��g�      A   ,  �r��g�  �r��s  ���s  ���g�  �r��g�      A   ,  ����g�  ����s  �j��s  �j��g�  ����g�      A   ,  ���g�  ���s  ����s  ����g�  ���g�      A   ,  �\��g�  �\��s  ���s  ���g�  �\��g�      A   ,  {���W�  {���c  |���c  |���W�  {���W�      A   ,  ~J��W�  ~J��c  ~���c  ~���W�  ~J��W�      A   ,  ����W�  ����c  �B��c  �B��W�  ����W�      A   ,  ����W�  ����c  ����c  ����W�  ����W�      A   ,  ����W�  ����c  �t��c  �t��W�  ����W�      A   ,  ���W�  ���c  ����c  ����W�  ���W�      A   ,  �f��W�  �f��c  ���c  ���W�  �f��W�      A   ,  ����W�  ����c  �^��c  �^��W�  ����W�      A   ,  ���W�  ���c  ����c  ����W�  ���W�      A   ,  �P��W�  �P��c  ����c  ����W�  �P��W�      A   ,  ����W�  ����c  �H��c  �H��W�  ����W�      A   ,  ����W�  ����c  ����c  ����W�  ����W�      A   ,  �:��W�  �:��c  ����c  ����W�  �:��W�      A   ,  ����W�  ����c  �2��c  �2��W�  ����W�      A   ,  ����W�  ����c  ����c  ����W�  ����W�      A   ,  �$��W�  �$��c  ����c  ����W�  �$��W�      A   ,  �r��W�  �r��c  ���c  ���W�  �r��W�      A   ,  ����W�  ����c  �j��c  �j��W�  ����W�      A   ,  ���W�  ���c  ����c  ����W�  ���W�      A   ,  �\��W�  �\��c  ���c  ���W�  �\��W�      A   , ���a� ���s ���s ���a� ���a�      A   , ���a� ���s |��s |��a� ���a�      A   , ���a� ���s `��s `��a� ���a�      A   , ���a� ���s D��s D��a� ���a�      A   , ~��a� ~��s (��s (��a� ~��a�      A   , b��a� b��s ��s ��a� b��a�      A   , F��a� F��s ���s ���a� F��a�      A   ,  *��a�  *��s  ���s  ���a�  *��a�      A   , #��a� #��s #���s #���a� #��a�      A   , %���a� %���s &���s &���a� %���a�      A   , (���a� (���s )���s )���a� (���a�      A   , +���a� +���s ,d��s ,d��a� +���a�      A   , .���a� .���s /H��s /H��a� .���a�      A   , 1���a� 1���s 2,��s 2,��a� 1���a�      A   , 4f��a� 4f��s 5��s 5��a� 4f��a�      A   , 7J��a� 7J��s 7���s 7���a� 7J��a�      A   , :.��a� :.��s :���s :���a� :.��a�      A   , =��a� =��s =���s =���a� =��a�      A   , ?���a� ?���s @���s @���a� ?���a�      A   , B���a� B���s C���s C���a� B���a�      A   , E���a� E���s Fh��s Fh��a� E���a�      A   , H���a� H���s IL��s IL��a� H���a�      A   , K���a� K���s L0��s L0��a� K���a�      A   , Nj��a� Nj��s O��s O��a� Nj��a�      A   , QN��a� QN��s Q���s Q���a� QN��a�      A   , T2��a� T2��s T���s T���a� T2��a�      A   , W��a� W��s W���s W���a� W��a�      A   , Y���a� Y���s Z���s Z���a� Y���a�      A   , \���a� \���s ]���s ]���a� \���a�      A   , _���a� _���s `l��s `l��a� _���a�      A   , b���a� b���s cP��s cP��a� b���a�      A   , e���a� e���s f4��s f4��a� e���a�      A   , hn��a� hn��s i��s i��a� hn��a�      A   , kR��a� kR��s k���s k���a� kR��a�      A   , n6��a� n6��s n���s n���a� n6��a�      A   , q��a� q��s q���s q���a� q��a�      A   , s���a� s���s t���s t���a� s���a�      A   , v���a� v���s w���s w���a� v���a�      A   , y���a� y���s zp��s zp��a� y���a�      A   , |���a� |���s }T��s }T��a� |���a�      A   , ���a� ���s �8��s �8��a� ���a�      A   , �r��a� �r��s ���s ���a� �r��a�      A   , �V��a� �V��s � ��s � ��a� �V��a�      A   , �:��a� �:��s ����s ����a� �:��a�      A   , ���a� ���s ����s ����a� ���a�      A   , ���a� ���s ����s ����a� ���a�      A   , ����a� ����s ����s ����a� ����a�      A   , ����a� ����s �t��s �t��a� ����a�      A   , ����a� ����s �X��s �X��a� ����a�      A   , ����a� ����s �<��s �<��a� ����a�      A   , �v��a� �v��s � ��s � ��a� �v��a�      A   , �Z��a� �Z��s ���s ���a� �Z��a�      A   , �>��a� �>��s ����s ����a� �>��a�      A   , �"��a� �"��s ����s ����a� �"��a�      A   , ���a� ���s ����s ����a� ���a�      A   , ����a� ����s ����s ����a� ����a�      A   , ����a� ����s �x��s �x��a� ����a�      A   , ����a� ����s �\��s �\��a� ����a�      A   , ����a� ����s �@��s �@��a� ����a�      A   , �z��a� �z��s �$��s �$��a� �z��a�      A   , �^��a� �^��s ���s ���a� �^��a�      A   , �B��a� �B��s ����s ����a� �B��a�      A   , �&��a� �&��s ����s ����a� �&��a�      A   , �
��a� �
��s ´��s ´��a� �
��a�      A   , �>��L# �>��]? ����]? ����L# �>��L#      A   , �"��L# �"��]? ����]? ����L# �"��L#      A   , ���L# ���]? ����]? ����L# ���L#      A   , ����L# ����]? ����]? ����L# ����L#      A   , ����L# ����]? �x��]? �x��L# ����L#      A   , ����L# ����]? �\��]? �\��L# ����L#      A   , ����L# ����]? �@��]? �@��L# ����L#      A   , �z��L# �z��]? �$��]? �$��L# �z��L#      A  , ,  ]   �  ]   �  Ҫ  �  Ҫ  �  ]   �      A  , ,  [�  '  [�  �  �  �  �  '  [�  '      A  , ,  [����I  [�  '  \b  '  \b���I  [����I      A  , ,  �h���I  �h  '  �  '  ����I  �h���I      A  , ,  [�����  [����I  ����I  �����  [�����      A  , ,  ] ����  ] ����  Ҫ����  Ҫ����  ] ����      A  , ,  ] ���/  ] ����  Ҫ����  Ҫ���/  ] ���/      A  , ,  [����  [�����  �����  ����  [����      A  , ,  [����?  [����  \b���  \b���?  [����?      A  , ,  �h���?  �h���  ����  ����?  �h���?      A  , ,  [���ϕ  [����?  ����?  ���ϕ  [���ϕ      A  , ,  ] ����  ] ��·  Ҫ��·  Ҫ����  ] ����      A  , ,  ] ���%  ] ����  Ҫ����  Ҫ���%  ] ���%      A  , ,  [����  [���ʽ  ���ʽ  ����  [����      A  , ,  [����5  [����  \b���  \b���5  [����5      A  , ,  �h���5  �h���  ����  ����5  �h���5      A  , ,  [�����  [����5  ����5  �����  [�����      A  , ,  ] ����  ] ���}  Ҫ���}  Ҫ����  ] ����      A  , ,  ] ���  ] ����  Ҫ����  Ҫ���  ] ���      A  , ,  ] ��}�  ] ��~s  Ҫ��~s  Ҫ��}�  ] ��}�      A  , ,  ] ��|  ] ��|�  Ҫ��|�  Ҫ��|  ] ��|      ^   ,  ��  (}  ��  4� .�  4� .�  (}  ��  (}      ^   , Mf  (} Mf  4� p  4� p  (} Mf  (}      ^   , ��  (} ��  4� ��  4� ��  (} ��  (}      ^   ,  ��  )  ��  $c .�  $c .�  )  ��  )      ^   , Mf  ) Mf  $c p  $c p  ) Mf  )      ^   , ��  ) ��  $c ��  $c ��  ) ��  )      ^   ,  ]9  	  ]9  �  ґ  �  ґ  	  ]9  	      ^   ,  ]9����  ]9  g  ґ  g  ґ����  ]9����      ^   ,  ]9����  ]9���  ґ���  ґ����  ]9����      ^   ,  ]9��ҫ  ]9���]  ґ���]  ґ��ҫ  ]9��ҫ      ^   ,  ]9����  ]9��ǧ  ґ��ǧ  ґ����  ]9����      ^   ,  ]9����  ]9���S  ґ���S  ґ����  ]9����      ^   ,  o����'  o����a  xs���a  xs���'  o����'      ^   ,  �m���'  �m���a  �k���a  �k���'  �m���'      ^   ,  o�����  o����  xs���  xs����  o�����      ^   ,  �m����  �m���  �k���  �k����  �m����      ]  , ,  \�  p  \�    �'    �'  p  \�  p      ]  , ,  [;  �  [;  p  ԏ  p  ԏ  �  [;  �      ]  , ,  [;����  [;  �  \�  �  \�����  [;����      ]  , ,  ������  ��  �  ԏ  �  ԏ����  ������      ]  , ,  [;���   [;����  ԏ����  ԏ���   [;���       ]  , ,  \�����  \����   �'���   �'����  \�����      ]  , ,  [;���  [;����  ԏ����  ԏ���  [;���      ]  , ,  [;��м  [;���  \����  \���м  [;��м      ]  , ,  ����м  �����  ԏ���  ԏ��м  ����м      ]  , ,  [;����  [;��м  ԏ��м  ԏ����  [;����      ]  , ,  \���̶  \�����  �'����  �'��̶  \���̶      ]  , ,  [;��ɖ  [;��̶  ԏ��̶  ԏ��ɖ  [;��ɖ      ]  , ,  [;����  [;��ɖ  \���ɖ  \�����  [;����      ]  , ,  ������  ����ɖ  ԏ��ɖ  ԏ����  ������      ]  , ,  [;����  [;����  ԏ����  ԏ����  [;����      ]  , ,  \�����  \�����  �'����  �'����  \�����      ]  , ,  [;���0  [;����  ԏ����  ԏ���0  [;���0      ]  , ,  [;��}�  [;��  ԏ��  ԏ��}�  [;��}�      ]  , ,  \���{�  \���}�  �'��}�  �'��{�  \���{�      ]  , ,  {��gX  {��s�  ���s�  ���gX  {��gX      ]  , ,  �M��gX  �M��s�  ����s�  ����gX  �M��gX      ]  , ,  {��W^  {��c�  ���c�  ���W^  {��W^      ]  , ,  �M��W^  �M��c�  ����c�  ����W^  �M��W^      ]  , , q��a| q��s� �1��s� �1��a| q��a|      ]  , , ����K� ����]� ����]� ����K� ����K�      B   ,  ^�����  ^�����  `����  `����  ^�����      B   ,  a&����  a&����  bR����  bR����  a&����      B   ,  ct����  ct����  d�����  d�����  ct����      B   ,  e�����  e�����  f�����  f�����  e�����      B   ,  h����  h����  i<����  i<����  h����      B   ,  j^����  j^����  k�����  k�����  j^����      B   ,  l�����  l�����  m�����  m�����  l�����      B   ,  n�����  n�����  p&����  p&����  n�����      B   ,  qH����  qH����  rt����  rt����  qH����      B   ,  s�����  s�����  t�����  t�����  s�����      B   ,  u�����  u�����  w����  w����  u�����      B   ,  x2����  x2����  y^����  y^����  x2����      B   ,  z�����  z�����  {�����  {�����  z�����      B   ,  |�����  |�����  }�����  }�����  |�����      B   ,  ����  ����  �H����  �H����  ����      B   ,  �j����  �j����  ������  ������  �j����      B   ,  ������  ������  ������  ������  ������      B   ,  �����  �����  �2����  �2����  �����      B   ,  �T����  �T����  ������  ������  �T����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  �����  �����  ������      B   ,  �>����  �>����  �j����  �j����  �>����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  �����  �����  ������      B   ,  �(����  �(����  �T����  �T����  �(����      B   ,  �v����  �v����  ������  ������  �v����      B   ,  ������  ������  ������  ������  ������      B   ,  �����  �����  �>����  �>����  �����      B   ,  �`����  �`����  ������  ������  �`����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  �(����  �(����  ������      B   ,  �J����  �J����  �v����  �v����  �J����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  �����  �����  ������      B   ,  �4����  �4����  �`����  �`����  �4����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  ������  ������  ������      B   ,  �����  �����  �J����  �J����  �����      B   ,  �l����  �l����  ������  ������  �l����      B   ,  ������  ������  ������  ������  ������      B   ,  �����  �����  �4����  �4����  �����      B   ,  �V����  �V����  ������  ������  �V����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  �����  �����  ������      B   ,  �@����  �@����  �l����  �l����  �@����      B   ,  Ǝ����  Ǝ����  Ǻ����  Ǻ����  Ǝ����      B   ,  ������  ������  �����  �����  ������      B   ,  �*����  �*����  �V����  �V����  �*����      B   ,  �x����  �x����  Τ����  Τ����  �x����      B   ,  ������  ������  ������  ������  ������      B   , ���]� ���aO B��aO B��]� ���]�      B   , ��  &� ��  (# ��  (# ��  &� ��  &�      B   , ��  &� ��  (# �  (# �  &� ��  &�      B   , �!  &� �!  (# �k  (# �k  &� �!  &�      B   , �o  &� �o  (# ǹ  (# ǹ  &� �o  &�      B   , Ƚ  &� Ƚ  (# �  (# �  &� Ƚ  &�      B   , �  &� �  (# �U  (# �U  &� �  &�      B   , �Y  &� �Y  (# Σ  (# Σ  &� �Y  &�      B   , s�  $� s�  & t�  & t�  $� s�  $�      B   , u�  $� u�  & w2  & w2  $� u�  $�      B   , x6  $� x6  & y�  & y�  $� x6  $�      B   , z�  $� z�  & {�  & {�  $� z�  $�      B   , |�  $� |�  & ~  & ~  $� |�  $�      B   , �k  $� �k  & ��  & ��  $� �k  $�      B   , ��  $� ��  & ��  & ��  $� ��  $�      B   , ��  $� ��  & �=  & �=  $� ��  $�      B   , �A  $� �A  & ��  & ��  $� �A  $�      B   , ��  $� ��  & ��  & ��  $� ��  $�      B   , ��  $� ��  & �'  & �'  $� ��  $�      B   , �+  $� �+  & �u  & �u  $� �+  $�      B   , �y  $� �y  & ��  & ��  $� �y  $�      B   , ��  $� ��  & �  & �  $� ��  $�      B   , �  $� �  & �_  & �_  $� �  $�      B   , �c  $� �c  & ��  & ��  $� �c  $�      B   , ��  $� ��  & ��  & ��  $� ��  $�      B   , ��  $� ��  & �I  & �I  $� ��  $�      B   , �M  $� �M  & ��  & ��  $� �M  $�      B   , ��  $� ��  & ��  & ��  $� ��  $�      B   , ��  $� ��  & �3  & �3  $� ��  $�      B   , �7  $� �7  & ��  & ��  $� �7  $�      B   , ��  $� ��  & ��  & ��  $� ��  $�      B   , ��  $� ��  & �  & �  $� ��  $�      B   , �!  $� �!  & �k  & �k  $� �!  $�      B   , �o  $� �o  & ǹ  & ǹ  $� �o  $�      B   , Ƚ  $� Ƚ  & �  & �  $� Ƚ  $�      B   , �  $� �  & �U  & �U  $� �  $�      B   , �Y  $� �Y  & Σ  & Σ  $� �Y  $�      B   , s�  &� s�  (# t�  (# t�  &� s�  &�      B   , u�  &� u�  (# w2  (# w2  &� u�  &�      B   , x6  &� x6  (# y�  (# y�  &� x6  &�      B   , z�  &� z�  (# {�  (# {�  &� z�  &�      B   , |�  &� |�  (# ~  (# ~  &� |�  &�      B   , �k  &� �k  '� ��  '� ��  &� �k  &�      B   , ��  &� ��  (# ��  (# ��  &� ��  &�      B   , ��  &� ��  (# �=  (# �=  &� ��  &�      B   , �A  &� �A  (# ��  (# ��  &� �A  &�      B   , ��  &� ��  (# ��  (# ��  &� ��  &�      B   , ��  &� ��  (# �'  (# �'  &� ��  &�      B   , �+  &� �+  (# �u  (# �u  &� �+  &�      B   , �y  &� �y  (# ��  (# ��  &� �y  &�      B   , ��  &� ��  (# �  (# �  &� ��  &�      B   , �  &� �  (# �_  (# �_  &� �  &�      B   , �c  &� �c  (# ��  (# ��  &� �c  &�      B   , ��  &� ��  (# ��  (# ��  &� ��  &�      B   , ��  &� ��  (# �I  (# �I  &� ��  &�      B   , �M  &� �M  (# ��  (# ��  &� �M  &�      B   , ��  &� ��  (# ��  (# ��  &� ��  &�      B   , ��  &� ��  (# �3  (# �3  &� ��  &�      B   , �7  &� �7  (# ��  (# ��  &� �7  &�      B   , cx  $� cx  & d�  & d�  $� cx  $�      B   , e�  $� e�  & g  & g  $� e�  $�      B   , h  $� h  & i^  & i^  $� h  $�      B   , jb  $� jb  & k�  & k�  $� jb  $�      B   , l�  $� l�  & m�  & m�  $� l�  $�      B   , n�  $� n�  & pH  & pH  $� n�  $�      B   , qL  $� qL  & r�  & r�  $� qL  $�      B   , �  &� �  (# �  (# �  &� �  &�      B   , �  &� �  (# %  (# %  &� �  &�      B   , )  &� )  (# s  (# s  &� )  &�      B   , w  &� w  (# �  (# �  &� w  &�      B   ,  �  &�  �  (# "  (# "  &�  �  &�      B   , #  &� #  (# $]  (# $]  &� #  &�      B   , %a  &� %a  (# &�  (# &�  &� %a  &�      B   , '�  &� '�  (# (�  (# (�  &� '�  &�      B   , )�  &� )�  (# +G  (# +G  &� )�  &�      B   , ,K  &� ,K  (# -�  (# -�  &� ,K  &�      B   , G�  &� G�  '� I  '� I  &� G�  &�      B   , J  &� J  (# Kh  (# Kh  &� J  &�      B   , Ll  &� Ll  (# M�  (# M�  &� Ll  &�      B   , N�  &� N�  (# P  (# P  &� N�  &�      B   , Q  &� Q  (# RR  (# RR  &� Q  &�      B   , SV  &� SV  (# T�  (# T�  &� SV  &�      B   , U�  &� U�  (# V�  (# V�  &� U�  &�      B   , W�  &� W�  (# Y<  (# Y<  &� W�  &�      B   , Z@  &� Z@  (# [�  (# [�  &� Z@  &�      B   , \�  &� \�  (# ]�  (# ]�  &� \�  &�      B   , ^�  &� ^�  (# `&  (# `&  &� ^�  &�      B   , a*  &� a*  (# bt  (# bt  &� a*  &�      B   , cx  &� cx  (# d�  (# d�  &� cx  &�      B   , e�  &� e�  (# g  (# g  &� e�  &�      B   , h  &� h  (# i^  (# i^  &� h  &�      B   , jb  &� jb  (# k�  (# k�  &� jb  &�      B   , l�  &� l�  (# m�  (# m�  &� l�  &�      B   , n�  &� n�  (# pH  (# pH  &� n�  &�      B   , qL  &� qL  (# r�  (# r�  &� qL  &�      B   , �  $� �  & �  & �  $� �  $�      B   , �  $� �  & %  & %  $� �  $�      B   , )  $� )  & s  & s  $� )  $�      B   , w  $� w  & �  & �  $� w  $�      B   ,  �  $�  �  & "  & "  $�  �  $�      B   , #  $� #  & $]  & $]  $� #  $�      B   , %a  $� %a  & &�  & &�  $� %a  $�      B   , '�  $� '�  & (�  & (�  $� '�  $�      B   , )�  $� )�  & +G  & +G  $� )�  $�      B   , ,K  $� ,K  & -�  & -�  $� ,K  $�      B   , G�  $� G�  & I  & I  $� G�  $�      B   , J  $� J  & Kh  & Kh  $� J  $�      B   , Ll  $� Ll  & M�  & M�  $� Ll  $�      B   , N�  $� N�  & P  & P  $� N�  $�      B   , Q  $� Q  & RR  & RR  $� Q  $�      B   , SV  $� SV  & T�  & T�  $� SV  $�      B   , U�  $� U�  & V�  & V�  $� U�  $�      B   , W�  $� W�  & Y<  & Y<  $� W�  $�      B   , Z@  $� Z@  & [�  & [�  $� Z@  $�      B   , \�  $� \�  & ]�  & ]�  $� \�  $�      B   , ^�  $� ^�  & `&  & `&  $� ^�  $�      B   , a*  $� a*  & bt  & bt  $� a*  $�      B   ,  �E  &�  �E  (  ��  (  ��  &�  �E  &�      B   ,  �G  �  �G  #  ��  #  ��  �  �G  �      B   ,  ��  �  ��  #  ��  #  ��  �  ��  �      B   ,  ��  �  ��  #  �-  #  �-  �  ��  �      B   ,  �1  �  �1  #  �{  #  �{  �  �1  �      B   ,  �  �  �  #  ��  #  ��  �  �  �      B   ,  ��  �  ��  #  �  #  �  �  ��  �      B   ,  �  �  �  #  �e  #  �e  �  �  �      B   ,  �i  �  �i  #  γ  #  γ  �  �i  �      B   ,  Ϸ  �  Ϸ  #  �  #  �  �  Ϸ  �      B   ,  �  
�  �  �  �4  �  �4  
�  �  
�      B   ,  �V  
�  �V  �  ��  �  ��  
�  �V  
�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  ��  
�  ��  �  �  �  �  
�  ��  
�      B   ,  �@  
�  �@  �  �l  �  �l  
�  �@  
�      B   ,  Ǝ  
�  Ǝ  �  Ǻ  �  Ǻ  
�  Ǝ  
�      B   ,  ��  
�  ��  �  �  �  �  
�  ��  
�      B   ,  �*  
�  �*  �  �V  �  �V  
�  �*  
�      B   ,  �x  
�  �x  �  Τ  �  Τ  
�  �x  
�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  ��  �  ��  
�  �C  
�  �C  �  ��  �      B   ,  �G  �  �G  
�  ��  
�  ��  �  �G  �      B   ,  ��  �  ��  
�  ��  
�  ��  �  ��  �      B   ,  ��  �  ��  
�  �-  
�  �-  �  ��  �      B   ,  �1  �  �1  
�  �{  
�  �{  �  �1  �      B   ,  �  �  �  
�  ��  
�  ��  �  �  �      B   ,  ��  �  ��  
�  �  
�  �  �  ��  �      B   ,  �  �  �  
�  �e  
�  �e  �  �  �      B   ,  �i  �  �i  
�  γ  
�  γ  �  �i  �      B   ,  Ϸ  �  Ϸ  
�  �  
�  �  �  Ϸ  �      B   ,  �����  �  �  �4  �  �4����  �����      B   ,  �V����  �V  �  ��  �  ������  �V����      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  ������  ��  �  �  �  �����  ������      B   ,  �@����  �@  �  �l  �  �l����  �@����      B   ,  Ǝ����  Ǝ  �  Ǻ  �  Ǻ����  Ǝ����      B   ,  ������  ��  �  �  �  �����  ������      B   ,  �*����  �*  �  �V  �  �V����  �*����      B   ,  �x����  �x  �  Τ  �  Τ����  �x����      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  �����M  ������  �C����  �C���M  �����M      B   ,  �G���M  �G����  ������  �����M  �G���M      B   ,  �����M  ������  ������  �����M  �����M      B   ,  �����M  ������  �-����  �-���M  �����M      B   ,  �1���M  �1����  �{����  �{���M  �1���M      B   ,  ����M  �����  ������  �����M  ����M      B   ,  �����M  ������  �����  ����M  �����M      B   ,  ����M  �����  �e����  �e���M  ����M      B   ,  �i���M  �i����  γ����  γ���M  �i���M      B   ,  Ϸ���M  Ϸ����  �����  ����M  Ϸ���M      B   , 	�  &� 	�  (#   (#   &� 	�  &�      B   ,   &�   (# Q  (# Q  &�   &�      B   , U  &� U  (# �  (# �  &� U  &�      B   , �  &� �  (# �  (# �  &� �  &�      B   , �  &� �  (# ;  (# ;  &� �  &�      B   , ?  &� ?  (# �  (# �  &� ?  &�      B   ,  ��  �  ��  #  �C  #  �C  �  ��  �      B   ,  ��  &�  ��  (  ��  (  ��  &�  ��  &�      B   ,  ��  &�  ��  (  �+  (  �+  &�  ��  &�      B   ,  �/  &�  �/  (  �y  (  �y  &�  �/  &�      B   ,  �}  &�  �}  (  ��  (  ��  &�  �}  &�      B   ,  ��  &�  ��  (  �  (  �  &�  ��  &�      B   ,  �  &�  �  (  �c  (  �c  &�  �  &�      B   ,  �]  $�  �]  &  �  &  �  $�  �]  $�      B   ,  ��  $�  ��  &  ��  &  ��  $�  ��  $�      B   ,  ��  $�  ��  &  �/  &  �/  $�  ��  $�      B   ,  �3  $�  �3  &  �}  &  �}  $�  �3  $�      B   ,  �  $�  �  & �  & �  $�  �  $�      B   , �  $� �  &   &   $� �  $�      B   ,   $�   & g  & g  $�   $�      B   , k  $� k  & �  & �  $� k  $�      B   , 	�  $� 	�  &   &   $� 	�  $�      B   ,   $�   & Q  & Q  $�   $�      B   , U  $� U  & �  & �  $� U  $�      B   , �  $� �  & �  & �  $� �  $�      B   , �  $� �  & ;  & ;  $� �  $�      B   , ?  $� ?  & �  & �  $� ?  $�      B   ,  �]  &�  �]  '�  �  '�  �  &�  �]  &�      B   ,  ��  &�  ��  (#  ��  (#  ��  &�  ��  &�      B   ,  ��  &�  ��  (#  �/  (#  �/  &�  ��  &�      B   ,  �3  &�  �3  (#  �}  (#  �}  &�  �3  &�      B   ,  �  &�  �  (# �  (# �  &�  �  &�      B   , �  &� �  (#   (#   &� �  &�      B   ,   &�   (# g  (# g  &�   &�      B   , k  &� k  (# �  (# �  &� k  &�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  �  
�  �  �  �J  �  �J  
�  �  
�      B   ,  �l  
�  �l  �  ��  �  ��  
�  �l  
�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  ^�  
�  ^�  �  `  �  `  
�  ^�  
�      B   ,  a&  
�  a&  �  bR  �  bR  
�  a&  
�      B   ,  ct  
�  ct  �  d�  �  d�  
�  ct  
�      B   ,  e�  
�  e�  �  f�  �  f�  
�  e�  
�      B   ,  h  
�  h  �  i<  �  i<  
�  h  
�      B   ,  j^  
�  j^  �  k�  �  k�  
�  j^  
�      B   ,  l�  
�  l�  �  m�  �  m�  
�  l�  
�      B   ,  n�  
�  n�  �  p&  �  p&  
�  n�  
�      B   ,  qH  
�  qH  �  rt  �  rt  
�  qH  
�      B   ,  s�  
�  s�  �  t�  �  t�  
�  s�  
�      B   ,  u�  
�  u�  �  w  �  w  
�  u�  
�      B   ,  x2  
�  x2  �  y^  �  y^  
�  x2  
�      B   ,  z�  
�  z�  �  {�  �  {�  
�  z�  
�      B   ,  |�  
�  |�  �  }�  �  }�  
�  |�  
�      B   ,    
�    �  �H  �  �H  
�    
�      B   ,  �j  
�  �j  �  ��  �  ��  
�  �j  
�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  �  
�  �  �  �2  �  �2  
�  �  
�      B   ,  �T  
�  �T  �  ��  �  ��  
�  �T  
�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  ��  
�  ��  �  �  �  �  
�  ��  
�      B   ,  �>  
�  �>  �  �j  �  �j  
�  �>  
�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  ��  
�  ��  �  �  �  �  
�  ��  
�      B   ,  �(  
�  �(  �  �T  �  �T  
�  �(  
�      B   ,  �v  
�  �v  �  ��  �  ��  
�  �v  
�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  �  
�  �  �  �>  �  �>  
�  �  
�      B   ,  �`  
�  �`  �  ��  �  ��  
�  �`  
�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  ��  
�  ��  �  �(  �  �(  
�  ��  
�      B   ,  �J  
�  �J  �  �v  �  �v  
�  �J  
�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  ��  
�  ��  �  �  �  �  
�  ��  
�      B   ,  �4  
�  �4  �  �`  �  �`  
�  �4  
�      B   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      B   ,  �q  &�  �q  (  ��  (  ��  &�  �q  &�      B   ,  ��  &�  ��  (  �	  (  �	  &�  ��  &�      B   ,  �  &�  �  (  �W  (  �W  &�  �  &�      B   ,  �[  &�  �[  (  ��  (  ��  &�  �[  &�      B   ,  ��  &�  ��  (  ��  (  ��  &�  ��  &�      B   ,  ��  &�  ��  (  �A  (  �A  &�  ��  &�      B   ,  �  �  �  #  �M  #  �M  �  �  �      B   ,  �Q  �  �Q  #  ��  #  ��  �  �Q  �      B   ,  ��  �  ��  #  ��  #  ��  �  ��  �      B   ,  ��  �  ��  #  �7  #  �7  �  ��  �      B   ,  �;  �  �;  #  ��  #  ��  �  �;  �      B   ,  ��  �  ��  #  ��  #  ��  �  ��  �      B   ,  ��  �  ��  #  �!  #  �!  �  ��  �      B   ,  �%  �  �%  #  �o  #  �o  �  �%  �      B   ,  �s  �  �s  #  ��  #  ��  �  �s  �      B   ,  ��  �  ��  #  �  #  �  �  ��  �      B   ,  �  �  �  #  �Y  #  �Y  �  �  �      B   ,  �]  �  �]  #  ��  #  ��  �  �]  �      B   ,  ��  �  ��  #  ��  #  ��  �  ��  �      B   ,  ��  �  ��  #  �+  #  �+  �  ��  �      B   ,  �/  �  �/  #  �y  #  �y  �  �/  �      B   ,  �}  �  �}  #  ��  #  ��  �  �}  �      B   ,  ��  �  ��  #  �  #  �  �  ��  �      B   ,  �  �  �  #  �c  #  �c  �  �  �      B   ,  �g  �  �g  #  ��  #  ��  �  �g  �      B   ,  ��  �  ��  #  ��  #  ��  �  ��  �      B   ,  �?  &�  �?  (  ��  (  ��  &�  �?  &�      B   ,  ��  &�  ��  (  ��  (  ��  &�  ��  &�      B   ,  ��  &�  ��  (  �%  (  �%  &�  ��  &�      B   ,  �)  &�  �)  (  �s  (  �s  &�  �)  &�      B   ,  �w  &�  �w  (  ��  (  ��  &�  �w  &�      B   ,  ��  &�  ��  (  �  (  �  &�  ��  &�      B   ,  �  &�  �  (  �]  (  �]  &�  �  &�      B   ,  ��  &�  ��  (  �  (  �  &�  ��  &�      B   ,  �#  &�  �#  (  �m  (  �m  &�  �#  &�      B   ,  jO  �  jO  #  k�  #  k�  �  jO  �      B   ,  l�  �  l�  #  m�  #  m�  �  l�  �      B   ,  n�  �  n�  #  p5  #  p5  �  n�  �      B   ,  q9  �  q9  #  r�  #  r�  �  q9  �      B   ,  s�  �  s�  #  t�  #  t�  �  s�  �      B   ,  u�  �  u�  #  w  #  w  �  u�  �      B   ,  |�  �  |�  #  ~	  #  ~	  �  |�  �      B   ,    �    #  �W  #  �W  �    �      B   ,  �[  �  �[  #  ��  #  ��  �  �[  �      B   ,  ��  �  ��  #  ��  #  ��  �  ��  �      B   ,  ��  �  ��  #  �A  #  �A  �  ��  �      B   ,  �E  �  �E  #  ��  #  ��  �  �E  �      B   ,  ��  �  ��  #  ��  #  ��  �  ��  �      B   ,  x#  �  x#  #  ym  #  ym  �  x#  �      B   ,  zq  �  zq  #  {�  #  {�  �  zq  �      B   ,  a  �  a  #  ba  #  ba  �  a  �      B   ,  ce  �  ce  #  d�  #  d�  �  ce  �      B   ,  e�  �  e�  #  f�  #  f�  �  e�  �      B   ,  h  �  h  #  iK  #  iK  �  h  �      B   ,  ^�  �  ^�  #  `  #  `  �  ^�  �      B   ,  a  �  a  
�  ba  
�  ba  �  a  �      B   ,  ce  �  ce  
�  d�  
�  d�  �  ce  �      B   ,  e�  �  e�  
�  f�  
�  f�  �  e�  �      B   ,  h  �  h  
�  iK  
�  iK  �  h  �      B   ,  jO  �  jO  
�  k�  
�  k�  �  jO  �      B   ,  l�  �  l�  
�  m�  
�  m�  �  l�  �      B   ,  n�  �  n�  
�  p5  
�  p5  �  n�  �      B   ,  q9  �  q9  
�  r�  
�  r�  �  q9  �      B   ,  s�  �  s�  
�  t�  
�  t�  �  s�  �      B   ,  ^�����  ^�  �  `  �  `����  ^�����      B   ,  a&����  a&  �  bR  �  bR����  a&����      B   ,  ct����  ct  �  d�  �  d�����  ct����      B   ,  e�����  e�  �  f�  �  f�����  e�����      B   ,  h����  h  �  i<  �  i<����  h����      B   ,  j^����  j^  �  k�  �  k�����  j^����      B   ,  l�����  l�  �  m�  �  m�����  l�����      B   ,  n�����  n�  �  p&  �  p&����  n�����      B   ,  qH����  qH  �  rt  �  rt����  qH����      B   ,  s�����  s�  �  t�  �  t�����  s�����      B   ,  u�����  u�  �  w  �  w����  u�����      B   ,  x2����  x2  �  y^  �  y^����  x2����      B   ,  z�����  z�  �  {�  �  {�����  z�����      B   ,  |�����  |�  �  }�  �  }�����  |�����      B   ,  ����    �  �H  �  �H����  ����      B   ,  �j����  �j  �  ��  �  ������  �j����      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  �����  �  �  �2  �  �2����  �����      B   ,  �T����  �T  �  ��  �  ������  �T����      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  u�  �  u�  
�  w  
�  w  �  u�  �      B   ,  x#  �  x#  
�  ym  
�  ym  �  x#  �      B   ,  zq  �  zq  
�  {�  
�  {�  �  zq  �      B   ,  |�  �  |�  
�  ~	  
�  ~	  �  |�  �      B   ,    �    
�  �W  
�  �W  �    �      B   ,  �[  �  �[  
�  ��  
�  ��  �  �[  �      B   ,  ��  �  ��  
�  ��  
�  ��  �  ��  �      B   ,  ��  �  ��  
�  �A  
�  �A  �  ��  �      B   ,  �E  �  �E  
�  ��  
�  ��  �  �E  �      B   ,  ��  �  ��  
�  ��  
�  ��  �  ��  �      B   ,  ^����M  ^�����  `����  `���M  ^����M      B   ,  a���M  a����  ba����  ba���M  a���M      B   ,  ce���M  ce����  d�����  d����M  ce���M      B   ,  e����M  e�����  f�����  f����M  e����M      B   ,  h���M  h����  iK����  iK���M  h���M      B   ,  jO���M  jO����  k�����  k����M  jO���M      B   ,  l����M  l�����  m�����  m����M  l����M      B   ,  n����M  n�����  p5����  p5���M  n����M      B   ,  q9���M  q9����  r�����  r����M  q9���M      B   ,  s����M  s�����  t�����  t����M  s����M      B   ,  u����M  u�����  w����  w���M  u����M      B   ,  x#���M  x#����  ym����  ym���M  x#���M      B   ,  zq���M  zq����  {�����  {����M  zq���M      B   ,  |����M  |�����  ~	����  ~	���M  |����M      B   ,  ���M  ����  �W����  �W���M  ���M      B   ,  �[���M  �[����  ������  �����M  �[���M      B   ,  �����M  ������  ������  �����M  �����M      B   ,  �����M  ������  �A����  �A���M  �����M      B   ,  �E���M  �E����  ������  �����M  �E���M      B   ,  �����M  ������  ������  �����M  �����M      B   ,  ^�  �  ^�  
�  `  
�  `  �  ^�  �      B   ,  �J����  �J  �  �v  �  �v����  �J����      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  ������  ��  �  �  �  �����  ������      B   ,  �4����  �4  �  �`  �  �`����  �4����      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  �����  �  �  �J  �  �J����  �����      B   ,  �l����  �l  �  ��  �  ������  �l����      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  ��  �  ��  
�  �7  
�  �7  �  ��  �      B   ,  �;  �  �;  
�  ��  
�  ��  �  �;  �      B   ,  ��  �  ��  
�  ��  
�  ��  �  ��  �      B   ,  ��  �  ��  
�  �!  
�  �!  �  ��  �      B   ,  �%  �  �%  
�  �o  
�  �o  �  �%  �      B   ,  �s  �  �s  
�  ��  
�  ��  �  �s  �      B   ,  ��  �  ��  
�  �  
�  �  �  ��  �      B   ,  �  �  �  
�  �Y  
�  �Y  �  �  �      B   ,  �]  �  �]  
�  ��  
�  ��  �  �]  �      B   ,  ��  �  ��  
�  ��  
�  ��  �  ��  �      B   ,  ��  �  ��  
�  �+  
�  �+  �  ��  �      B   ,  �/  �  �/  
�  �y  
�  �y  �  �/  �      B   ,  �}  �  �}  
�  ��  
�  ��  �  �}  �      B   ,  ��  �  ��  
�  �  
�  �  �  ��  �      B   ,  �  �  �  
�  �c  
�  �c  �  �  �      B   ,  �g  �  �g  
�  ��  
�  ��  �  �g  �      B   ,  ��  �  ��  
�  ��  
�  ��  �  ��  �      B   ,  �  �  �  
�  �M  
�  �M  �  �  �      B   ,  �Q  �  �Q  
�  ��  
�  ��  �  �Q  �      B   ,  ��  �  ��  
�  ��  
�  ��  �  ��  �      B   ,  ������  ��  �  �  �  �����  ������      B   ,  �>����  �>  �  �j  �  �j����  �>����      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  ������  ��  �  �  �  �����  ������      B   ,  �(����  �(  �  �T  �  �T����  �(����      B   ,  �v����  �v  �  ��  �  ������  �v����      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  �����  �  �  �>  �  �>����  �����      B   ,  �`����  �`  �  ��  �  ������  �`����      B   ,  ������  ��  �  ��  �  ������  ������      B   ,  �����M  ������  �+����  �+���M  �����M      B   ,  �/���M  �/����  �y����  �y���M  �/���M      B   ,  �}���M  �}����  ������  �����M  �}���M      B   ,  �����M  ������  �����  ����M  �����M      B   ,  ����M  �����  �c����  �c���M  ����M      B   ,  �g���M  �g����  ������  �����M  �g���M      B   ,  �����M  ������  ������  �����M  �����M      B   ,  ����M  �����  �M����  �M���M  ����M      B   ,  �Q���M  �Q����  ������  �����M  �Q���M      B   ,  �����M  ������  ������  �����M  �����M      B   ,  �����M  ������  �7����  �7���M  �����M      B   ,  �;���M  �;����  ������  �����M  �;���M      B   ,  �����M  ������  ������  �����M  �����M      B   ,  �����M  ������  �!����  �!���M  �����M      B   ,  �%���M  �%����  �o����  �o���M  �%���M      B   ,  �s���M  �s����  ������  �����M  �s���M      B   ,  �����M  ������  �����  ����M  �����M      B   ,  ����M  �����  �Y����  �Y���M  ����M      B   ,  �]���M  �]����  ������  �����M  �]���M      B   ,  �����M  ������  ������  �����M  �����M      B   ,  ������  ��  �  �(  �  �(����  ������      B   ,  ^���ҍ  ^����{  `���{  `��ҍ  ^���ҍ      B   ,  a&��ҍ  a&���{  bR���{  bR��ҍ  a&��ҍ      B   ,  ct��ҍ  ct���{  d����{  d���ҍ  ct��ҍ      B   ,  e���ҍ  e����{  f����{  f���ҍ  e���ҍ      B   ,  h��ҍ  h���{  i<���{  i<��ҍ  h��ҍ      B   ,  j^��ҍ  j^���{  k����{  k���ҍ  j^��ҍ      B   ,  l���ҍ  l����{  m����{  m���ҍ  l���ҍ      B   ,  n���ҍ  n����{  p&���{  p&��ҍ  n���ҍ      B   ,  qH��ҍ  qH���{  rt���{  rt��ҍ  qH��ҍ      B   ,  s���ҍ  s����{  t����{  t���ҍ  s���ҍ      B   ,  u���ҍ  u����{  w���{  w��ҍ  u���ҍ      B   ,  x2��ҍ  x2���{  y^���{  y^��ҍ  x2��ҍ      B   ,  z���ҍ  z����{  {����{  {���ҍ  z���ҍ      B   ,  |���ҍ  |����{  }����{  }���ҍ  |���ҍ      B   ,  ��ҍ  ���{  �H���{  �H��ҍ  ��ҍ      B   ,  �j��ҍ  �j���{  �����{  ����ҍ  �j��ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ���ҍ  ����{  �2���{  �2��ҍ  ���ҍ      B   ,  �T��ҍ  �T���{  �����{  ����ҍ  �T��ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ����ҍ  �����{  ����{  ���ҍ  ����ҍ      B   ,  �>��ҍ  �>���{  �j���{  �j��ҍ  �>��ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ����ҍ  �����{  ����{  ���ҍ  ����ҍ      B   ,  �(��ҍ  �(���{  �T���{  �T��ҍ  �(��ҍ      B   ,  �v��ҍ  �v���{  �����{  ����ҍ  �v��ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ���ҍ  ����{  �>���{  �>��ҍ  ���ҍ      B   ,  �`��ҍ  �`���{  �����{  ����ҍ  �`��ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ����ҍ  �����{  �(���{  �(��ҍ  ����ҍ      B   ,  �J��ҍ  �J���{  �v���{  �v��ҍ  �J��ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ����ҍ  �����{  ����{  ���ҍ  ����ҍ      B   ,  �4��ҍ  �4���{  �`���{  �`��ҍ  �4��ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ���ҍ  ����{  �J���{  �J��ҍ  ���ҍ      B   ,  �l��ҍ  �l���{  �����{  ����ҍ  �l��ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ������  ������  �����  �����  ������      B   ,  �>����  �>����  �j����  �j����  �>����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  �����  �����  ������      B   ,  �(����  �(����  �T����  �T����  �(����      B   ,  �v����  �v����  ������  ������  �v����      B   ,  ������  ������  ������  ������  ������      B   ,  �����  �����  �>����  �>����  �����      B   ,  �`����  �`����  ������  ������  �`����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  �(����  �(����  ������      B   ,  �J����  �J����  �v����  �v����  �J����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  �����  �����  ������      B   ,  �4����  �4����  �`����  �`����  �4����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  ������  ������  ������      B   ,  �����  �����  �J����  �J����  �����      B   ,  �l����  �l����  ������  ������  �l����      B   ,  ������  ������  ������  ������  ������      B   ,  �����{  ������  �+����  �+���{  �����{      B   ,  �/���{  �/����  �y����  �y���{  �/���{      B   ,  �}���{  �}����  ������  �����{  �}���{      B   ,  �����{  ������  �����  ����{  �����{      B   ,  ����{  �����  �c����  �c���{  ����{      B   ,  �g���{  �g����  ������  �����{  �g���{      B   ,  �����{  ������  ������  �����{  �����{      B   ,  ����{  �����  �M����  �M���{  ����{      B   ,  �Q���{  �Q����  ������  �����{  �Q���{      B   ,  �����{  ������  ������  �����{  �����{      B   ,  �����{  ������  �7����  �7���{  �����{      B   ,  �;���{  �;����  ������  �����{  �;���{      B   ,  �����{  ������  ������  �����{  �����{      B   ,  �����{  ������  �!����  �!���{  �����{      B   ,  �%���{  �%����  �o����  �o���{  �%���{      B   ,  �s���{  �s����  ������  �����{  �s���{      B   ,  �����{  ������  �����  ����{  �����{      B   ,  ����{  �����  �Y����  �Y���{  ����{      B   ,  �]���{  �]����  ������  �����{  �]���{      B   ,  �����{  ������  ������  �����{  �����{      B   ,  ������  �����  �+���  �+����  ������      B   ,  �/����  �/���  �y���  �y����  �/����      B   ,  �}����  �}���  �����  ������  �}����      B   ,  ������  �����  ����  �����  ������      B   ,  �����  ����  �c���  �c����  �����      B   ,  �g����  �g���  �����  ������  �g����      B   ,  ������  �����  �����  ������  ������      B   ,  �����  ����  �M���  �M����  �����      B   ,  �Q����  �Q���  �����  ������  �Q����      B   ,  ������  �����  �����  ������  ������      B   ,  ������  �����  �7���  �7����  ������      B   ,  �;����  �;���  �����  ������  �;����      B   ,  ������  �����  �����  ������  ������      B   ,  ������  �����  �!���  �!����  ������      B   ,  �%����  �%���  �o���  �o����  �%����      B   ,  �s����  �s���  �����  ������  �s����      B   ,  ������  �����  ����  �����  ������      B   ,  �����  ����  �Y���  �Y����  �����      B   ,  �]����  �]���  �����  ������  �]����      B   ,  ������  �����  �����  ������  ������      B   ,  |����{  |�����  ~	����  ~	���{  |����{      B   ,  ���{  ����  �W����  �W���{  ���{      B   ,  �[���{  �[����  ������  �����{  �[���{      B   ,  �����{  ������  ������  �����{  �����{      B   ,  �����{  ������  �A����  �A���{  �����{      B   ,  �E���{  �E����  ������  �����{  �E���{      B   ,  �����{  ������  ������  �����{  �����{      B   ,  |�����  |�����  }�����  }�����  |�����      B   ,  ����  ����  �H����  �H����  ����      B   ,  ^�����  ^����  `���  `����  ^�����      B   ,  a����  a���  ba���  ba����  a����      B   ,  ce����  ce���  d����  d�����  ce����      B   ,  e�����  e����  f����  f�����  e�����      B   ,  h����  h���  iK���  iK����  h����      B   ,  jO����  jO���  k����  k�����  jO����      B   ,  l�����  l����  m����  m�����  l�����      B   ,  n�����  n����  p5���  p5����  n�����      B   ,  q9����  q9���  r����  r�����  q9����      B   ,  s�����  s����  t����  t�����  s�����      B   ,  u�����  u����  w���  w����  u�����      B   ,  x#����  x#���  ym���  ym����  x#����      B   ,  zq����  zq���  {����  {�����  zq����      B   ,  |�����  |����  ~	���  ~	����  |�����      B   ,  ����  ���  �W���  �W����  ����      B   ,  �[����  �[���  �����  ������  �[����      B   ,  ������  �����  �����  ������  ������      B   ,  ������  �����  �A���  �A����  ������      B   ,  �E����  �E���  �����  ������  �E����      B   ,  ������  �����  �����  ������  ������      B   ,  �j����  �j����  ������  ������  �j����      B   ,  ������  ������  ������  ������  ������      B   ,  �����  �����  �2����  �2����  �����      B   ,  �T����  �T����  ������  ������  �T����      B   ,  ������  ������  ������  ������  ������      B   ,  x2����  x2����  y^����  y^����  x2����      B   ,  z�����  z�����  {�����  {�����  z�����      B   ,  ^����{  ^�����  `����  `���{  ^����{      B   ,  a���{  a����  ba����  ba���{  a���{      B   ,  ce���{  ce����  d�����  d����{  ce���{      B   ,  e����{  e�����  f�����  f����{  e����{      B   ,  h���{  h����  iK����  iK���{  h���{      B   ,  jO���{  jO����  k�����  k����{  jO���{      B   ,  l����{  l�����  m�����  m����{  l����{      B   ,  n����{  n�����  p5����  p5���{  n����{      B   ,  q9���{  q9����  r�����  r����{  q9���{      B   ,  s����{  s�����  t�����  t����{  s����{      B   ,  u����{  u�����  w����  w���{  u����{      B   ,  x#���{  x#����  ym����  ym���{  x#���{      B   ,  zq���{  zq����  {�����  {����{  zq���{      B   ,  ^�����  ^�����  `����  `����  ^�����      B   ,  a&����  a&����  bR����  bR����  a&����      B   ,  ct����  ct����  d�����  d�����  ct����      B   ,  e�����  e�����  f�����  f�����  e�����      B   ,  h����  h����  i<����  i<����  h����      B   ,  j^����  j^����  k�����  k�����  j^����      B   ,  l�����  l�����  m�����  m�����  l�����      B   ,  n�����  n�����  p&����  p&����  n�����      B   ,  qH����  qH����  rt����  rt����  qH����      B   ,  s�����  s�����  t�����  t�����  s�����      B   ,  u�����  u�����  w����  w����  u�����      B   ,  x#���C  x#��ҍ  ym��ҍ  ym���C  x#���C      B   ,  zq���C  zq��ҍ  {���ҍ  {����C  zq���C      B   ,  |����C  |���ҍ  ~	��ҍ  ~	���C  |����C      B   ,  ���C  ��ҍ  �W��ҍ  �W���C  ���C      B   ,  �[���C  �[��ҍ  ����ҍ  �����C  �[���C      B   ,  �����C  ����ҍ  ����ҍ  �����C  �����C      B   ,  �����C  ����ҍ  �A��ҍ  �A���C  �����C      B   ,  �E���C  �E��ҍ  ����ҍ  �����C  �E���C      B   ,  �����C  ����ҍ  ����ҍ  �����C  �����C      B   ,  ^�����  ^����  `���  `����  ^�����      B   ,  a����  a���  ba���  ba����  a����      B   ,  ce����  ce���  d����  d�����  ce����      B   ,  e�����  e����  f����  f�����  e�����      B   ,  h����  h���  iK���  iK����  h����      B   ,  jO����  jO���  k����  k�����  jO����      B   ,  l�����  l����  m����  m�����  l�����      B   ,  n�����  n����  p5���  p5����  n�����      B   ,  q9����  q9���  r����  r�����  q9����      B   ,  s�����  s����  t����  t�����  s�����      B   ,  u�����  u����  w���  w����  u�����      B   ,  x#����  x#���  ym���  ym����  x#����      B   ,  zq����  zq���  {����  {�����  zq����      B   ,  |�����  |����  ~	���  ~	����  |�����      B   ,  ����  ���  �W���  �W����  ����      B   ,  �[����  �[���  �����  ������  �[����      B   ,  ������  �����  �����  ������  ������      B   ,  ������  �����  �A���  �A����  ������      B   ,  �E����  �E���  �����  ������  �E����      B   ,  ������  �����  �����  ������  ������      B   ,  ^����C  ^���ҍ  `��ҍ  `���C  ^����C      B   ,  a���C  a��ҍ  ba��ҍ  ba���C  a���C      B   ,  ce���C  ce��ҍ  d���ҍ  d����C  ce���C      B   ,  e����C  e���ҍ  f���ҍ  f����C  e����C      B   ,  h���C  h��ҍ  iK��ҍ  iK���C  h���C      B   ,  jO���C  jO��ҍ  k���ҍ  k����C  jO���C      B   ,  l����C  l���ҍ  m���ҍ  m����C  l����C      B   ,  n����C  n���ҍ  p5��ҍ  p5���C  n����C      B   ,  q9���C  q9��ҍ  r���ҍ  r����C  q9���C      B   ,  s����C  s���ҍ  t���ҍ  t����C  s����C      B   ,  u����C  u���ҍ  w��ҍ  w���C  u����C      B   ,  �;���C  �;��ҍ  ����ҍ  �����C  �;���C      B   ,  �����C  ����ҍ  ����ҍ  �����C  �����C      B   ,  �����C  ����ҍ  �!��ҍ  �!���C  �����C      B   ,  �%���C  �%��ҍ  �o��ҍ  �o���C  �%���C      B   ,  �s���C  �s��ҍ  ����ҍ  �����C  �s���C      B   ,  �����C  ����ҍ  ���ҍ  ����C  �����C      B   ,  ����C  ���ҍ  �Y��ҍ  �Y���C  ����C      B   ,  �]���C  �]��ҍ  ����ҍ  �����C  �]���C      B   ,  �����C  ����ҍ  ����ҍ  �����C  �����C      B   ,  ������  �����  �+���  �+����  ������      B   ,  �/����  �/���  �y���  �y����  �/����      B   ,  �}����  �}���  �����  ������  �}����      B   ,  ������  �����  ����  �����  ������      B   ,  �����  ����  �c���  �c����  �����      B   ,  �g����  �g���  �����  ������  �g����      B   ,  ������  �����  �����  ������  ������      B   ,  �����  ����  �M���  �M����  �����      B   ,  �Q����  �Q���  �����  ������  �Q����      B   ,  ������  �����  �����  ������  ������      B   ,  ������  �����  �7���  �7����  ������      B   ,  �;����  �;���  �����  ������  �;����      B   ,  ������  �����  �����  ������  ������      B   ,  ������  �����  �!���  �!����  ������      B   ,  �%����  �%���  �o���  �o����  �%����      B   ,  �s����  �s���  �����  ������  �s����      B   ,  ������  �����  ����  �����  ������      B   ,  �����  ����  �Y���  �Y����  �����      B   ,  �]����  �]���  �����  ������  �]����      B   ,  ������  �����  �����  ������  ������      B   ,  �����C  ����ҍ  �+��ҍ  �+���C  �����C      B   ,  �/���C  �/��ҍ  �y��ҍ  �y���C  �/���C      B   ,  �}���C  �}��ҍ  ����ҍ  �����C  �}���C      B   ,  �����C  ����ҍ  ���ҍ  ����C  �����C      B   ,  ����C  ���ҍ  �c��ҍ  �c���C  ����C      B   ,  �g���C  �g��ҍ  ����ҍ  �����C  �g���C      B   ,  �����C  ����ҍ  ����ҍ  �����C  �����C      B   ,  ����C  ���ҍ  �M��ҍ  �M���C  ����C      B   ,  �Q���C  �Q��ҍ  ����ҍ  �����C  �Q���C      B   ,  �����C  ����ҍ  ����ҍ  �����C  �����C      B   ,  �����C  ����ҍ  �7��ҍ  �7���C  �����C      B   ,  �G����  �G���  �����  ������  �G����      B   ,  ������  �����  �����  ������  ������      B   ,  ������  �����  �-���  �-����  ������      B   ,  �1����  �1���  �{���  �{����  �1����      B   ,  �����  ����  �����  ������  �����      B   ,  ������  �����  ����  �����  ������      B   ,  �����  ����  �e���  �e����  �����      B   ,  �i����  �i���  γ���  γ����  �i����      B   ,  Ϸ����  Ϸ���  ����  �����  Ϸ����      B   ,  �����C  ����ҍ  �C��ҍ  �C���C  �����C      B   ,  �G���C  �G��ҍ  ����ҍ  �����C  �G���C      B   ,  �����C  ����ҍ  ����ҍ  �����C  �����C      B   ,  �����C  ����ҍ  �-��ҍ  �-���C  �����C      B   ,  �1���C  �1��ҍ  �{��ҍ  �{���C  �1���C      B   ,  ����C  ���ҍ  ����ҍ  �����C  ����C      B   ,  �����C  ����ҍ  ���ҍ  ����C  �����C      B   ,  ����C  ���ҍ  �e��ҍ  �e���C  ����C      B   ,  �i���C  �i��ҍ  γ��ҍ  γ���C  �i���C      B   ,  Ϸ���C  Ϸ��ҍ  ���ҍ  ����C  Ϸ���C      B   ,  �����  �����  �4����  �4����  �����      B   ,  �V����  �V����  ������  ������  �V����      B   ,  ������  ������  ������  ������  ������      B   ,  ������  ������  �����  �����  ������      B   ,  �@����  �@����  �l����  �l����  �@����      B   ,  Ǝ����  Ǝ����  Ǻ����  Ǻ����  Ǝ����      B   ,  ������  ������  �����  �����  ������      B   ,  �*����  �*����  �V����  �V����  �*����      B   ,  �x����  �x����  Τ����  Τ����  �x����      B   ,  ������  ������  ������  ������  ������      B   ,  �����{  ������  �C����  �C���{  �����{      B   ,  �G���{  �G����  ������  �����{  �G���{      B   ,  �����{  ������  ������  �����{  �����{      B   ,  �����{  ������  �-����  �-���{  �����{      B   ,  �1���{  �1����  �{����  �{���{  �1���{      B   ,  ����{  �����  ������  �����{  ����{      B   ,  �����{  ������  �����  ����{  �����{      B   ,  ����{  �����  �e����  �e���{  ����{      B   ,  �i���{  �i����  γ����  γ���{  �i���{      B   ,  Ϸ���{  Ϸ����  �����  ����{  Ϸ���{      B   ,  ������  �����  �C���  �C����  ������      B   ,  �G����  �G���  �����  ������  �G����      B   ,  ������  �����  �����  ������  ������      B   ,  ������  �����  �-���  �-����  ������      B   ,  �1����  �1���  �{���  �{����  �1����      B   ,  �����  ����  �����  ������  �����      B   ,  ������  �����  ����  �����  ������      B   ,  �����  ����  �e���  �e����  �����      B   ,  �i����  �i���  γ���  γ����  �i����      B   ,  Ϸ����  Ϸ���  ����  �����  Ϸ����      B   ,  ���ҍ  ����{  �4���{  �4��ҍ  ���ҍ      B   ,  �V��ҍ  �V���{  �����{  ����ҍ  �V��ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ����ҍ  �����{  ����{  ���ҍ  ����ҍ      B   ,  �@��ҍ  �@���{  �l���{  �l��ҍ  �@��ҍ      B   ,  Ǝ��ҍ  Ǝ���{  Ǻ���{  Ǻ��ҍ  Ǝ��ҍ      B   ,  ����ҍ  �����{  ����{  ���ҍ  ����ҍ      B   ,  �*��ҍ  �*���{  �V���{  �V��ҍ  �*��ҍ      B   ,  �x��ҍ  �x���{  Τ���{  Τ��ҍ  �x��ҍ      B   ,  ����ҍ  �����{  �����{  ����ҍ  ����ҍ      B   ,  ������  �����  �C���  �C����  ������      B   ,  ^����g  ^�����  `����  `���g  ^����g      B   ,  a���g  a����  ba����  ba���g  a���g      B   ,  ce���g  ce����  d�����  d����g  ce���g      B   ,  e����g  e�����  f�����  f����g  e����g      B   ,  h���g  h����  iK����  iK���g  h���g      B   ,  jO���g  jO����  k�����  k����g  jO���g      B   ,  l����g  l�����  m�����  m����g  l����g      B   ,  n����g  n�����  p5����  p5���g  n����g      B   ,  q9���g  q9����  r�����  r����g  q9���g      B   ,  s����g  s�����  t�����  t����g  s����g      B   ,  u����g  u�����  w����  w���g  u����g      B   ,  x#���g  x#����  ym����  ym���g  x#���g      B   ,  zq���g  zq����  {�����  {����g  zq���g      B   ,  |����g  |�����  ~	����  ~	���g  |����g      B   ,  ���g  ����  �W����  �W���g  ���g      B   ,  �[���g  �[����  ������  �����g  �[���g      B   ,  �����g  ������  ������  �����g  �����g      B   ,  �����g  ������  �A����  �A���g  �����g      B   ,  �E���g  �E����  ������  �����g  �E���g      B   ,  �����g  ������  ������  �����g  �����g      B   ,  �����g  ������  �+����  �+���g  �����g      B   ,  �/���g  �/����  �y����  �y���g  �/���g      B   ,  �}���g  �}����  ������  �����g  �}���g      B   ,  �����g  ������  �����  ����g  �����g      B   ,  ����g  �����  �c����  �c���g  ����g      B   ,  �g���g  �g����  ������  �����g  �g���g      B   ,  �����g  ������  ������  �����g  �����g      B   ,  ����g  �����  �M����  �M���g  ����g      B   ,  �Q���g  �Q����  ������  �����g  �Q���g      B   ,  �����g  ������  ������  �����g  �����g      B   ,  �����g  ������  �7����  �7���g  �����g      B   ,  �;���g  �;����  ������  �����g  �;���g      B   ,  �����g  ������  ������  �����g  �����g      B   ,  �����g  ������  �!����  �!���g  �����g      B   ,  �%���g  �%����  �o����  �o���g  �%���g      B   ,  �s���g  �s����  ������  �����g  �s���g      B   ,  �����g  ������  �����  ����g  �����g      B   ,  ����g  �����  �Y����  �Y���g  ����g      B   ,  �]���g  �]����  ������  �����g  �]���g      B   ,  �����g  ������  ������  �����g  �����g      B   ,  �����g  ������  �C����  �C���g  �����g      B   ,  �G���g  �G����  ������  �����g  �G���g      B   ,  �����g  ������  ������  �����g  �����g      B   ,  �����g  ������  �-����  �-���g  �����g      B   ,  �1���g  �1����  �{����  �{���g  �1���g      B   ,  ����g  �����  ������  �����g  ����g      B   ,  �����g  ������  �����  ����g  �����g      B   ,  ����g  �����  �e����  �e���g  ����g      B   ,  �i���g  �i����  γ����  γ���g  �i���g      B   ,  Ϸ���g  Ϸ����  �����  ����g  Ϸ���g      B   ,  �����9  ������  �C����  �C���9  �����9      B   ,  �G���9  �G����  ������  �����9  �G���9      B   ,  �����9  ������  ������  �����9  �����9      B   ,  �����9  ������  �-����  �-���9  �����9      B   ,  �1���9  �1����  �{����  �{���9  �1���9      B   ,  ����9  �����  ������  �����9  ����9      B   ,  �����9  ������  �����  ����9  �����9      B   ,  ����9  �����  �e����  �e���9  ����9      B   ,  �i���9  �i����  γ����  γ���9  �i���9      B   ,  Ϸ���9  Ϸ����  �����  ����9  Ϸ���9      B   ,  �����q  ������  �C����  �C���q  �����q      B   ,  �G���q  �G����  ������  �����q  �G���q      B   ,  �����q  ������  ������  �����q  �����q      B   ,  �����q  ������  �-����  �-���q  �����q      B   ,  �1���q  �1����  �{����  �{���q  �1���q      B   ,  ����q  �����  ������  �����q  ����q      B   ,  �����q  ������  �����  ����q  �����q      B   ,  ����q  �����  �e����  �e���q  ����q      B   ,  �i���q  �i����  γ����  γ���q  �i���q      B   ,  Ϸ���q  Ϸ����  �����  ����q  Ϸ���q      B   ,  �����  ����q  �4���q  �4����  �����      B   ,  �V����  �V���q  �����q  ������  �V����      B   ,  ������  �����q  �����q  ������  ������      B   ,  ������  �����q  ����q  �����  ������      B   ,  �@����  �@���q  �l���q  �l����  �@����      B   ,  Ǝ����  Ǝ���q  Ǻ���q  Ǻ����  Ǝ����      B   ,  ������  �����q  ����q  �����  ������      B   ,  �*����  �*���q  �V���q  �V����  �*����      B   ,  �x����  �x���q  Τ���q  Τ����  �x����      B   ,  ������  �����q  �����q  ������  ������      B   ,  ^����9  ^�����  `����  `���9  ^����9      B   ,  a���9  a����  ba����  ba���9  a���9      B   ,  ce���9  ce����  d�����  d����9  ce���9      B   ,  e����9  e�����  f�����  f����9  e����9      B   ,  h���9  h����  iK����  iK���9  h���9      B   ,  jO���9  jO����  k�����  k����9  jO���9      B   ,  l����9  l�����  m�����  m����9  l����9      B   ,  n����9  n�����  p5����  p5���9  n����9      B   ,  q9���9  q9����  r�����  r����9  q9���9      B   ,  s����9  s�����  t�����  t����9  s����9      B   ,  u����9  u�����  w����  w���9  u����9      B   ,  x#���9  x#����  ym����  ym���9  x#���9      B   ,  zq���9  zq����  {�����  {����9  zq���9      B   ,  |����9  |�����  ~	����  ~	���9  |����9      B   ,  ���9  ����  �W����  �W���9  ���9      B   ,  �[���9  �[����  ������  �����9  �[���9      B   ,  �����9  ������  ������  �����9  �����9      B   ,  �����9  ������  �A����  �A���9  �����9      B   ,  �E���9  �E����  ������  �����9  �E���9      B   ,  �����9  ������  ������  �����9  �����9      B   ,  �����9  ������  �+����  �+���9  �����9      B   ,  �/���9  �/����  �y����  �y���9  �/���9      B   ,  �}���9  �}����  ������  �����9  �}���9      B   ,  �����9  ������  �����  ����9  �����9      B   ,  ����9  �����  �c����  �c���9  ����9      B   ,  �g���9  �g����  ������  �����9  �g���9      B   ,  �����9  ������  ������  �����9  �����9      B   ,  ����9  �����  �M����  �M���9  ����9      B   ,  �Q���9  �Q����  ������  �����9  �Q���9      B   ,  �����9  ������  ������  �����9  �����9      B   ,  �����9  ������  �7����  �7���9  �����9      B   ,  �;���9  �;����  ������  �����9  �;���9      B   ,  �����9  ������  ������  �����9  �����9      B   ,  �����9  ������  �!����  �!���9  �����9      B   ,  �%���9  �%����  �o����  �o���9  �%���9      B   ,  �s���9  �s����  ������  �����9  �s���9      B   ,  �����9  ������  �����  ����9  �����9      B   ,  ����9  �����  �Y����  �Y���9  ����9      B   ,  �]���9  �]����  ������  �����9  �]���9      B   ,  �����9  ������  ������  �����9  �����9      B   ,  �J����  �J���q  �v���q  �v����  �J����      B   ,  ������  �����q  �����q  ������  ������      B   ,  ������  �����q  ����q  �����  ������      B   ,  �4����  �4���q  �`���q  �`����  �4����      B   ,  ������  �����q  �����q  ������  ������      B   ,  ������  �����q  �����q  ������  ������      B   ,  �����  ����q  �J���q  �J����  �����      B   ,  �l����  �l���q  �����q  ������  �l����      B   ,  ������  �����q  �����q  ������  ������      B   ,  �����q  ������  �+����  �+���q  �����q      B   ,  �/���q  �/����  �y����  �y���q  �/���q      B   ,  �}���q  �}����  ������  �����q  �}���q      B   ,  �����q  ������  �����  ����q  �����q      B   ,  ����q  �����  �c����  �c���q  ����q      B   ,  �g���q  �g����  ������  �����q  �g���q      B   ,  �����q  ������  ������  �����q  �����q      B   ,  ����q  �����  �M����  �M���q  ����q      B   ,  �Q���q  �Q����  ������  �����q  �Q���q      B   ,  �����q  ������  ������  �����q  �����q      B   ,  �����q  ������  �7����  �7���q  �����q      B   ,  �;���q  �;����  ������  �����q  �;���q      B   ,  �����q  ������  ������  �����q  �����q      B   ,  �����q  ������  �!����  �!���q  �����q      B   ,  �%���q  �%����  �o����  �o���q  �%���q      B   ,  �s���q  �s����  ������  �����q  �s���q      B   ,  �����q  ������  �����  ����q  �����q      B   ,  ����q  �����  �Y����  �Y���q  ����q      B   ,  �]���q  �]����  ������  �����q  �]���q      B   ,  �����q  ������  ������  �����q  �����q      B   ,  ������  �����q  ����q  �����  ������      B   ,  �>����  �>���q  �j���q  �j����  �>����      B   ,  ������  �����q  �����q  ������  ������      B   ,  ������  �����q  ����q  �����  ������      B   ,  �(����  �(���q  �T���q  �T����  �(����      B   ,  �v����  �v���q  �����q  ������  �v����      B   ,  ������  �����q  �����q  ������  ������      B   ,  �����  ����q  �>���q  �>����  �����      B   ,  �`����  �`���q  �����q  ������  �`����      B   ,  ������  �����q  �����q  ������  ������      B   ,  ������  �����q  �(���q  �(����  ������      B   ,  e����q  e�����  f�����  f����q  e����q      B   ,  h���q  h����  iK����  iK���q  h���q      B   ,  jO���q  jO����  k�����  k����q  jO���q      B   ,  l����q  l�����  m�����  m����q  l����q      B   ,  n����q  n�����  p5����  p5���q  n����q      B   ,  q9���q  q9����  r�����  r����q  q9���q      B   ,  s����q  s�����  t�����  t����q  s����q      B   ,  u����q  u�����  w����  w���q  u����q      B   ,  ^�����  ^����q  `���q  `����  ^�����      B   ,  a&����  a&���q  bR���q  bR����  a&����      B   ,  ct����  ct���q  d����q  d�����  ct����      B   ,  e�����  e����q  f����q  f�����  e�����      B   ,  h����  h���q  i<���q  i<����  h����      B   ,  j^����  j^���q  k����q  k�����  j^����      B   ,  l�����  l����q  m����q  m�����  l�����      B   ,  n�����  n����q  p&���q  p&����  n�����      B   ,  qH����  qH���q  rt���q  rt����  qH����      B   ,  s�����  s����q  t����q  t�����  s�����      B   ,  u�����  u����q  w���q  w����  u�����      B   ,  x2����  x2���q  y^���q  y^����  x2����      B   ,  z�����  z����q  {����q  {�����  z�����      B   ,  |�����  |����q  }����q  }�����  |�����      B   ,  ����  ���q  �H���q  �H����  ����      B   ,  �j����  �j���q  �����q  ������  �j����      B   ,  ������  �����q  �����q  ������  ������      B   ,  �����  ����q  �2���q  �2����  �����      B   ,  �T����  �T���q  �����q  ������  �T����      B   ,  ������  �����q  �����q  ������  ������      B   ,  �����q  ������  �A����  �A���q  �����q      B   ,  �E���q  �E����  ������  �����q  �E���q      B   ,  �����q  ������  ������  �����q  �����q      B   ,  x#���q  x#����  ym����  ym���q  x#���q      B   ,  zq���q  zq����  {�����  {����q  zq���q      B   ,  |����q  |�����  ~	����  ~	���q  |����q      B   ,  ���q  ����  �W����  �W���q  ���q      B   ,  �[���q  �[����  ������  �����q  �[���q      B   ,  �����q  ������  ������  �����q  �����q      B   ,  a���q  a����  ba����  ba���q  a���q      B   ,  ce���q  ce����  d�����  d����q  ce���q      B   ,  ^����q  ^�����  `����  `���q  ^����q      B   ,  u���c�  u���g+  w3��g+  w3��c�  u���c�      B   ,  x7��c�  x7��g+  y���g+  y���c�  x7��c�      B   ,  z���c�  z���g+  {���g+  {���c�  z���c�      B   ,  |���c�  |���g+  ~��g+  ~��c�  |���c�      B   ,  !��c�  !��g+  �k��g+  �k��c�  !��c�      B   ,  �o��c�  �o��g+  ����g+  ����c�  �o��c�      B   ,  ����c�  ����g+  ���g+  ���c�  ����c�      B   ,  ���c�  ���g+  �U��g+  �U��c�  ���c�      B   ,  �Y��c�  �Y��g+  ����g+  ����c�  �Y��c�      B   ,  ����c�  ����g+  ����g+  ����c�  ����c�      B   ,  s���c�  s���g+  t���g+  t���c�  s���c�      B   ,  �C��c�  �C��g+  ����g+  ����c�  �C��c�      B   ,  ����c�  ����g+  ����g+  ����c�  ����c�      B   ,  ����c�  ����g+  �)��g+  �)��c�  ����c�      B   ,  ����f�  ����g+  ����g+  ����f�  ����f�      B   ,  ����f1  ����f�  ����f�  ����f1  ����f1      B   ,  ����f1  ����f�  ����f�  ����f1  ����f1      B   ,  ����d�  ����f1  ����f1  ����d�  ����d�      B   ,  ����d  ����d�  ����d�  ����d  ����d      B   ,  ����d  ����d�  ����d�  ����d  ����d      B   ,  ����c�  ����d  ����d  ����c�  ����c�      B   ,  ����f�  ����g+  �9��g+  �9��f�  ����f�      B   ,  ����f1  ����f�  �?��f�  �?��f1  ����f1      B   ,  ����f1  ����f�  �9��f�  �9��f1  ����f1      B   ,  ����d�  ����f1  �9��f1  �9��d�  ����d�      B   ,  ����d  ����d�  �?��d�  �?��d  ����d      B   ,  ����d  ����d�  �9��d�  �9��d  ����d      B   ,  ����c�  ����d  �9��d  �9��c�  ����c�      B   ,  �=��f�  �=��g+  ����g+  ����f�  �=��f�      B   ,  �=��f1  �=��f�  ����f�  ����f1  �=��f1      B   ,  �7��f1  �7��f�  ����f�  ����f1  �7��f1      B   ,  �=��d�  �=��f1  ����f1  ����d�  �=��d�      B   ,  �=��d  �=��d�  ����d�  ����d  �=��d      B   ,  �7��d  �7��d�  ����d�  ����d  �7��d      B   ,  �=��c�  �=��d  ����d  ����c�  �=��c�      B   ,  ����f�  ����g+  ����g+  ����f�  ����f�      B   ,  ����f1  ����f�  ����f�  ����f1  ����f1      B   ,  ����f1  ����f�  ����f�  ����f1  ����f1      B   ,  ����d�  ����f1  ����f1  ����d�  ����d�      B   ,  ����d  ����d�  ����d�  ����d  ����d      B   ,  ����d  ����d�  ����d�  ����d  ����d      B   ,  ����c�  ����d  ����d  ����c�  ����c�      B   ,  ����c�  ����g+  �?��g+  �?��c�  ����c�      B   ,  ����f1  ����f�  �)��f�  �)��f1  ����f1      B   ,  ����f1  ����f�  �#��f�  �#��f1  ����f1      B   ,  ����d�  ����f1  �#��f1  �#��d�  ����d�      B   ,  ����d  ����d�  �)��d�  �)��d  ����d      B   ,  ����d  ����d�  �#��d�  �#��d  ����d      B   ,  ����c�  ����d  �#��d  �#��c�  ����c�      B   ,  �'��f�  �'��g+  �q��g+  �q��f�  �'��f�      B   ,  �'��f1  �'��f�  �w��f�  �w��f1  �'��f1      B   ,  �!��f1  �!��f�  �q��f�  �q��f1  �!��f1      B   ,  �'��d�  �'��f1  �q��f1  �q��d�  �'��d�      B   ,  �'��d  �'��d�  �w��d�  �w��d  �'��d      B   ,  �!��d  �!��d�  �q��d�  �q��d  �!��d      B   ,  �'��c�  �'��d  �q��d  �q��c�  �'��c�      B   ,  �u��f�  �u��g+  ����g+  ����f�  �u��f�      B   ,  �u��f1  �u��f�  ����f�  ����f1  �u��f1      B   ,  �o��f1  �o��f�  ����f�  ����f1  �o��f1      B   ,  �u��d�  �u��f1  ����f1  ����d�  �u��d�      B   ,  �u��d  �u��d�  ����d�  ����d  �u��d      B   ,  �o��d  �o��d�  ����d�  ����d  �o��d      B   ,  �u��c�  �u��d  ����d  ����c�  �u��c�      B   ,  ����f�  ����g+  ���g+  ���f�  ����f�      B   ,  ����f1  ����f�  ���f�  ���f1  ����f1      B   ,  ����f1  ����f�  ���f�  ���f1  ����f1      B   ,  ����d�  ����f1  ���f1  ���d�  ����d�      B   ,  ����d  ����d�  ���d�  ���d  ����d      B   ,  ����d  ����d�  ���d�  ���d  ����d      B   ,  ����c�  ����d  ���d  ���c�  ����c�      B   ,  ���f�  ���g+  �[��g+  �[��f�  ���f�      B   ,  ���f1  ���f�  �a��f�  �a��f1  ���f1      B   ,  ���f1  ���f�  �[��f�  �[��f1  ���f1      B   ,  ���d�  ���f1  �[��f1  �[��d�  ���d�      B   ,  ���d  ���d�  �a��d�  �a��d  ���d      B   ,  ���d  ���d�  �[��d�  �[��d  ���d      B   ,  ���c�  ���d  �[��d  �[��c�  ���c�      B   ,  �_��f�  �_��g+  ����g+  ����f�  �_��f�      B   ,  �_��f1  �_��f�  ����f�  ����f1  �_��f1      B   ,  �Y��f1  �Y��f�  ����f�  ����f1  �Y��f1      B   ,  �_��d�  �_��f1  ����f1  ����d�  �_��d�      B   ,  �_��d  �_��d�  ����d�  ����d  �_��d      B   ,  �Y��d  �Y��d�  ����d�  ����d  �Y��d      B   ,  �_��c�  �_��d  ����d  ����c�  �_��c�      B   ,  ����f�  ����g+  ����g+  ����f�  ����f�      B   ,  ����f1  ����f�  ����f�  ����f1  ����f1      B   ,  ����f1  ����f�  ����f�  ����f1  ����f1      B   ,  ����d�  ����f1  ����f1  ����d�  ����d�      B   ,  ����d  ����d�  ����d�  ����d  ����d      B   ,  ����d  ����d�  ����d�  ����d  ����d      B   ,  ����c�  ����d  ����d  ����c�  ����c�      B   ,  ����f�  ����g+  �E��g+  �E��f�  ����f�      B   ,  ����f1  ����f�  �K��f�  �K��f1  ����f1      B   ,  ����f1  ����f�  �E��f�  �E��f1  ����f1      B   ,  ����d�  ����f1  �E��f1  �E��d�  ����d�      B   ,  ����d  ����d�  �K��d�  �K��d  ����d      B   ,  ����d  ����d�  �E��d�  �E��d  ����d      B   ,  ����c�  ����d  �E��d  �E��c�  ����c�      B   ,  �I��f�  �I��g+  ����g+  ����f�  �I��f�      B   ,  �I��f1  �I��f�  ����f�  ����f1  �I��f1      B   ,  �C��f1  �C��f�  ����f�  ����f1  �C��f1      B   ,  �I��d�  �I��f1  ����f1  ����d�  �I��d�      B   ,  �I��d  �I��d�  ����d�  ����d  �I��d      B   ,  �C��d  �C��d�  ����d�  ����d  �C��d      B   ,  �I��c�  �I��d  ����d  ����c�  �I��c�      B   ,  ����f�  ����g+  ����g+  ����f�  ����f�      B   ,  ����f1  ����f�  ����f�  ����f1  ����f1      B   ,  ����f1  ����f�  ����f�  ����f1  ����f1      B   ,  ����d�  ����f1  ����f1  ����d�  ����d�      B   ,  ����d  ����d�  ����d�  ����d  ����d      B   ,  ����d  ����d�  ����d�  ����d  ����d      B   ,  ����c�  ����d  ����d  ����c�  ����c�      B   ,  ����f�  ����g+  �#��g+  �#��f�  ����f�      B   ,  ����f1  ����f�  �5��f�  �5��f1  ����f1      B   ,  ����f1  ����f�  �/��f�  �/��f1  ����f1      B   ,  ����d�  ����f1  �/��f1  �/��d�  ����d�      B   ,  ����d  ����d�  �5��d�  �5��d  ����d      B   ,  ����d  ����d�  �/��d�  �/��d  ����d      B   ,  ����c�  ����d  �/��d  �/��c�  ����c�      B   ,  ����^  ����a  �v��a  �v��^  ����^      B   ,  ����]�  ����aO  �Z��aO  �Z��]�  ����]�      B   ,  �|��]�  �|��aO  �>��aO  �>��]�  �|��]�      B   ,  �`��]�  �`��aO  "��aO  "��]�  �`��]�      B   , D��]� D��aO ��aO ��]� D��]�      B   , (��]� (��aO ���aO ���]� (��]�      B   , ��]� ��aO ���aO ���]� ��]�      B   , 	���]� 	���aO ���aO ���]� 	���]�      B   , ���]� ���aO ���aO ���]� ���]�      B   , ���]� ���aO z��aO z��]� ���]�      B   , ���]� ���aO ^��aO ^��]� ���]�      B   ,  ����f�  ����g+  �/��g+  �/��f�  ����f�      B   , r ��`� r ��aO s���aO s���`� r ��`�      B   , r ��^� r ��`U s���`U s���^� r ��^�      B   , r ��]� r ��^9 s���^9 s���]� r ��]�      B   , ,��`U ,��`� |��`� |��`U ,��`U      B   , ���`U ���`� ���`� ���`U ���`U      B   , ,��^� ,��`U ���`U ���^� ,��^�      B   , ,��^9 ,��^� |��^� |��^9 ,��^9      B   , ���^9 ���^� ���^� ���^9 ���^9      B   , ,��]� ,��^9 ���^9 ���]� ,��]�      B   , !��`� !��aO "���aO "���`� !��`�      B   , !��`U !��`� !`��`� !`��`U !��`U      B   , "���`U "���`� "���`� "���`U "���`U      B   , !��^� !��`U "���`U "���^� !��^�      B   , !��^9 !��^� !`��^� !`��^9 !��^9      B   , "���^9 "���^� "���^� "���^9 "���^9      B   , !��]� !��^9 "���^9 "���]� !��]�      B   , #���`� #���aO %���aO %���`� #���`�      B   , #���`U #���`� $D��`� $D��`U #���`U      B   , %f��`U %f��`� %���`� %���`U %f��`U      B   , #���^� #���`U %���`U %���^� #���^�      B   , #���^9 #���^� $D��^� $D��^9 #���^9      B   , %f��^9 %f��^� %���^� %���^9 %f��^9      B   , #���]� #���^9 %���^9 %���]� #���]�      B   , &���`� &���aO (���aO (���`� &���`�      B   , &���`U &���`� '(��`� '(��`U &���`U      B   , (J��`U (J��`� (���`� (���`U (J��`U      B   , &���^� &���`U (���`U (���^� &���^�      B   , &���^9 &���^� '(��^� '(��^9 &���^9      B   , (J��^9 (J��^� (���^� (���^9 (J��^9      B   , &���]� &���^9 (���^9 (���]� &���]�      B   , )���`� )���aO +~��aO +~��`� )���`�      B   , )���`U )���`� *��`� *��`U )���`U      B   , +.��`U +.��`� +~��`� +~��`U +.��`U      B   , )���^� )���`U +~��`U +~��^� )���^�      B   , )���^9 )���^� *��^� *��^9 )���^9      B   , +.��^9 +.��^� +~��^� +~��^9 +.��^9      B   , )���]� )���^9 +~��^9 +~��]� )���]�      B   , ,���`� ,���aO .b��aO .b��`� ,���`�      B   , ,���`U ,���`� ,���`� ,���`U ,���`U      B   , .��`U .��`� .b��`� .b��`U .��`U      B   , ,���^� ,���`U .b��`U .b��^� ,���^�      B   , ,���^9 ,���^� ,���^� ,���^9 ,���^9      B   , .��^9 .��^� .b��^� .b��^9 .��^9      B   , ,���]� ,���^9 .b��^9 .b��]� ,���]�      B   , /���]� /���aO 1F��aO 1F��]� /���]�      B   , 2h��]� 2h��aO 4*��aO 4*��]� 2h��]�      B   , 5L��]� 5L��aO 7��aO 7��]� 5L��]�      B   , 80��]� 80��aO 9���aO 9���]� 80��]�      B   , ;��]� ;��aO <���aO <���]� ;��]�      B   , =���]� =���aO ?���aO ?���]� =���]�      B   , @���]� @���aO B���aO B���]� @���]�      B   , C���]� C���aO E���aO E���]� C���]�      B   , F���]� F���aO Hf��aO Hf��]� F���]�      B   , I���]� I���aO KJ��aO KJ��]� I���]�      B   , Ll��]� Ll��aO N.��aO N.��]� Ll��]�      B   , OP��]� OP��aO Q��aO Q��]� OP��]�      B   , R4��]� R4��aO S���aO S���]� R4��]�      B   , U��]� U��aO V���aO V���]� U��]�      B   , W���]� W���aO Y���aO Y���]� W���]�      B   , Z���]� Z���aO \���aO \���]� Z���]�      B   , ]���]� ]���aO _���aO _���]� ]���]�      B   , `���]� `���aO bj��aO bj��]� `���]�      B   , c���]� c���aO eN��aO eN��]� c���]�      B   , fp��]� fp��aO h2��aO h2��]� fp��]�      B   , iT��`� iT��aO k��aO k��`� iT��`�      B   , iT��`U iT��`� i���`� i���`U iT��`U      B   , j���`U j���`� k��`� k��`U j���`U      B   , iT��^� iT��`U k��`U k��^� iT��^�      B   , iT��^9 iT��^� i���^� i���^9 iT��^9      B   , j���^9 j���^� k��^� k��^9 j���^9      B   , iT��]� iT��^9 k��^9 k��]� iT��]�      B   , l8��`� l8��aO m���aO m���`� l8��`�      B   , l8��`U l8��`� l���`� l���`U l8��`U      B   , m���`U m���`� m���`� m���`U m���`U      B   , l8��^� l8��`U m���`U m���^� l8��^�      B   , l8��^9 l8��^� l���^� l���^9 l8��^9      B   , m���^9 m���^� m���^� m���^9 m���^9      B   , l8��]� l8��^9 m���^9 m���]� l8��]�      B   , o��`� o��aO p���aO p���`� o��`�      B   , o��`U o��`� ol��`� ol��`U o��`U      B   , p���`U p���`� p���`� p���`U p���`U      B   , o��^� o��`U p���`U p���^� o��^�      B   , o��^9 o��^� ol��^� ol��^9 o��^9      B   , p���^9 p���^� p���^� p���^9 p���^9      B   , o��]� o��^9 p���^9 p���]� o��]�      B   , d��]� d��aO &��aO &��]� d��]�      B   , r ��`U r ��`� rP��`� rP��`U r ��`U      B   , H��]� H��aO 
��aO 
��]� H��]�      B   , r ��^9 r ��^� rP��^� rP��^9 r ��^9      B   , ,��`� ,��aO ���aO ���`� ,��`�      B   , �@��`� �@��aO ���aO ���`� �@��`�      B   , �@��^� �@��`U ���`U ���^� �@��^�      B   , �@��]� �@��^9 ���^9 ���]� �@��]�      B   , t���`U t���`� u4��`� u4��`U t���`U      B   , vV��`U vV��`� v���`� v���`U vV��`U      B   , t���^� t���`U v���`U v���^� t���^�      B   , t���^9 t���^� u4��^� u4��^9 t���^9      B   , vV��^9 vV��^� v���^� v���^9 vV��^9      B   , t���]� t���^9 v���^9 v���]� t���]�      B   , w���]� w���aO y���aO y���]� w���]�      B   , z���]� z���aO |n��aO |n��]� z���]�      B   , }���]� }���aO R��aO R��]� }���]�      B   , �t��]� �t��aO �6��aO �6��]� �t��]�      B   , �X��`� �X��aO ���aO ���`� �X��`�      B   , �X��`U �X��`� ����`� ����`U �X��`U      B   , ����`U ����`� ���`� ���`U ����`U      B   , �X��^� �X��`U ���`U ���^� �X��^�      B   , �X��^9 �X��^� ����^� ����^9 �X��^9      B   , ����^9 ����^� ���^� ���^9 ����^9      B   , �X��]� �X��^9 ���^9 ���]� �X��]�      B   , �<��`� �<��aO ����aO ����`� �<��`�      B   , �<��`U �<��`� ����`� ����`U �<��`U      B   , ����`U ����`� ����`� ����`U ����`U      B   , �<��^� �<��`U ����`U ����^� �<��^�      B   , �<��^9 �<��^� ����^� ����^9 �<��^9      B   , ����^9 ����^� ����^� ����^9 ����^9      B   , �<��]� �<��^9 ����^9 ����]� �<��]�      B   , � ��`� � ��aO ����aO ����`� � ��`�      B   , � ��`U � ��`� �p��`� �p��`U � ��`U      B   , ����`U ����`� ����`� ����`U ����`U      B   , � ��^� � ��`U ����`U ����^� � ��^�      B   , � ��^9 � ��^� �p��^� �p��^9 � ��^9      B   , ����^9 ����^� ����^� ����^9 ����^9      B   , � ��]� � ��^9 ����^9 ����]� � ��]�      B   , ���`� ���aO ����aO ����`� ���`�      B   , ���`U ���`� �T��`� �T��`U ���`U      B   , �v��`U �v��`� ����`� ����`U �v��`U      B   , ���^� ���`U ����`U ����^� ���^�      B   , ���^9 ���^� �T��^� �T��^9 ���^9      B   , �v��^9 �v��^� ����^� ����^9 �v��^9      B   , ���]� ���^9 ����^9 ����]� ���]�      B   , ����`� ����aO ����aO ����`� ����`�      B   , ����`U ����`� �8��`� �8��`U ����`U      B   , �Z��`U �Z��`� ����`� ����`U �Z��`U      B   , ����^� ����`U ����`U ����^� ����^�      B   , ����^9 ����^� �8��^� �8��^9 ����^9      B   , �Z��^9 �Z��^� ����^� ����^9 �Z��^9      B   , ����]� ����^9 ����^9 ����]� ����]�      B   , ����`� ����aO ����aO ����`� ����`�      B   , ����`U ����`� ���`� ���`U ����`U      B   , �>��`U �>��`� ����`� ����`U �>��`U      B   , ����^� ����`U ����`U ����^� ����^�      B   , ����^9 ����^� ���^� ���^9 ����^9      B   , �>��^9 �>��^� ����^� ����^9 �>��^9      B   , ����]� ����^9 ����^9 ����]� ����]�      B   , ����`� ����aO �r��aO �r��`� ����`�      B   , ����`U ����`� � ��`� � ��`U ����`U      B   , �"��`U �"��`� �r��`� �r��`U �"��`U      B   , ����^� ����`U �r��`U �r��^� ����^�      B   , ����^9 ����^� � ��^� � ��^9 ����^9      B   , �"��^9 �"��^� �r��^� �r��^9 �"��^9      B   , ����]� ����^9 �r��^9 �r��]� ����]�      B   , ����`� ����aO �V��aO �V��`� ����`�      B   , ����`U ����`� ����`� ����`U ����`U      B   , ���`U ���`� �V��`� �V��`U ���`U      B   , ����^� ����`U �V��`U �V��^� ����^�      B   , ����^9 ����^� ����^� ����^9 ����^9      B   , ���^9 ���^� �V��^� �V��^9 ���^9      B   , ����]� ����^9 �V��^9 �V��]� ����]�      B   , �x��`� �x��aO �:��aO �:��`� �x��`�      B   , �x��`U �x��`� ����`� ����`U �x��`U      B   , ����`U ����`� �:��`� �:��`U ����`U      B   , �x��^� �x��`U �:��`U �:��^� �x��^�      B   , �x��^9 �x��^� ����^� ����^9 �x��^9      B   , ����^9 ����^� �:��^� �:��^9 ����^9      B   , �x��]� �x��^9 �:��^9 �:��]� �x��]�      B   , �\��`� �\��aO ���aO ���`� �\��`�      B   , �\��`U �\��`� ����`� ����`U �\��`U      B   , ����`U ����`� ���`� ���`U ����`U      B   , �\��^� �\��`U ���`U ���^� �\��^�      B   , �\��^9 �\��^� ����^� ����^9 �\��^9      B   , ����^9 ����^� ���^� ���^9 ����^9      B   , �\��]� �\��^9 ���^9 ���]� �\��]�      B   , sr��^9 sr��^� s���^� s���^9 sr��^9      B   , �@��`U �@��`� ����`� ����`U �@��`U      B   , sr��`U sr��`� s���`� s���`U sr��`U      B   , �@��^9 �@��^� ����^� ����^9 �@��^9      B   , t���`� t���aO v���aO v���`� t���`�      B   , �`��`� �`��aO �"��aO �"��`� �`��`�      B   , �`��`U �`��`� ����`� ����`U �`��`U      B   , �`��^� �`��`U �"��`U �"��^� �`��^�      B   , �`��^9 �`��^� ����^� ����^9 �`��^9      B   , �`��]� �`��^9 �"��^9 �"��]� �`��]�      B   , �$��^� �$��`U ����`U ����^� �$��^�      B   , �$��^9 �$��^� �t��^� �t��^9 �$��^9      B   , ����^9 ����^� ����^� ����^9 ����^9      B   , �$��]� �$��^9 ����^9 ����]� �$��]�      B   , ���`� ���aO ����aO ����`� ���`�      B   , ���`U ���`� �X��`� �X��`U ���`U      B   , �z��`U �z��`� ����`� ����`U �z��`U      B   , ���^� ���`U ����`U ����^� ���^�      B   , ���^9 ���^� �X��^� �X��^9 ���^9      B   , �z��^9 �z��^� ����^� ����^9 �z��^9      B   , ���]� ���^9 ����^9 ����]� ���]�      B   , ����`� ����aO ����aO ����`� ����`�      B   , ����`U ����`� �<��`� �<��`U ����`U      B   , �^��`U �^��`� ����`� ����`U �^��`U      B   , ����^� ����`U ����`U ����^� ����^�      B   , ����^9 ����^� �<��^� �<��^9 ����^9      B   , �^��^9 �^��^� ����^� ����^9 �^��^9      B   , ����]� ����^9 ����^9 ����]� ����]�      B   , ����`� ����aO ����aO ����`� ����`�      B   , ����`U ����`� � ��`� � ��`U ����`U      B   , �B��`U �B��`� ����`� ����`U �B��`U      B   , ����^� ����`U ����`U ����^� ����^�      B   , ����^9 ����^� � ��^� � ��^9 ����^9      B   , �B��^9 �B��^� ����^� ����^9 �B��^9      B   , ����]� ����^9 ����^9 ����]� ����]�      B   , ����`� ����aO �v��aO �v��`� ����`�      B   , ����`U ����`� ���`� ���`U ����`U      B   , �&��`U �&��`� �v��`� �v��`U �&��`U      B   , ����^� ����`U �v��`U �v��^� ����^�      B   , ����^9 ����^� ���^� ���^9 ����^9      B   , �&��^9 �&��^� �v��^� �v��^9 �&��^9      B   , ����]� ����^9 �v��^9 �v��]� ����]�      B   , ����`� ����aO �Z��aO �Z��`� ����`�      B   , ����`U ����`� ����`� ����`U ����`U      B   , �
��`U �
��`� �Z��`� �Z��`U �
��`U      B   , ����^� ����`U �Z��`U �Z��^� ����^�      B   , ����^9 ����^� ����^� ����^9 ����^9      B   , �
��^9 �
��^� �Z��^� �Z��^9 �
��^9      B   , ����]� ����^9 �Z��^9 �Z��]� ����]�      B   , �|��`� �|��aO �>��aO �>��`� �|��`�      B   , �|��`U �|��`� ����`� ����`U �|��`U      B   , ����`U ����`� �>��`� �>��`U ����`U      B   , �|��^� �|��`U �>��`U �>��^� �|��^�      B   , �|��^9 �|��^� ����^� ����^9 �|��^9      B   , ����^9 ����^� �>��^� �>��^9 ����^9      B   , �|��]� �|��^9 �>��^9 �>��]� �|��]�      B   , ����^9 ����^� ���^� ���^9 ����^9      B   , ����`U ����`� ���`� ���`U ����`U      B   , �$��`� �$��aO ����aO ����`� �$��`�      B   , �$��`U �$��`� �t��`� �t��`U �$��`U      B   , ����`U ����`� ����`� ����`U ����`U      B   , ����^9 ����^� �"��^� �"��^9 ����^9      B   , ����`U ����`� �"��`� �"��`U ����`U      B   , �D��`� �D��aO ���aO ���`� �D��`�      B   , �D��`U �D��`� ����`� ����`U �D��`U      B   , ����`U ����`� ���`� ���`U ����`U      B   , �D��^� �D��`U ���`U ���^� �D��^�      B   , �D��^9 �D��^� ����^� ����^9 �D��^9      B   , ����^9 ����^� ���^� ���^9 ����^9      B   , �D��]� �D��^9 ���^9 ���]� �D��]�      B   , �(��`� �(��aO ����aO ����`� �(��`�      B   , �(��`U �(��`� �x��`� �x��`U �(��`U      B   , ����`U ����`� ����`� ����`U ����`U      B   , �(��^� �(��`U ����`U ����^� �(��^�      B   , �(��^9 �(��^� �x��^� �x��^9 �(��^9      B   , ����^9 ����^� ����^� ����^9 ����^9      B   , �(��]� �(��^9 ����^9 ����]� �(��]�      B   , ���`� ���aO ����aO ����`� ���`�      B   , ���`U ���`� �\��`� �\��`U ���`U      B   , �~��`U �~��`� ����`� ����`U �~��`U      B   , ���^� ���`U ����`U ����^� ���^�      B   , ���^9 ���^� �\��^� �\��^9 ���^9      B   , �~��^9 �~��^� ����^� ����^9 �~��^9      B   , ���]� ���^9 ����^9 ����]� ���]�      B   , ����`� ����aO Ĳ��aO Ĳ��`� ����`�      B   , ����`U ����`� �@��`� �@��`U ����`U      B   , �b��`U �b��`� Ĳ��`� Ĳ��`U �b��`U      B   , ����^� ����`U Ĳ��`U Ĳ��^� ����^�      B   , ����^9 ����^� �@��^� �@��^9 ����^9      B   , �b��^9 �b��^� Ĳ��^� Ĳ��^9 �b��^9      B   , ����]� ����^9 Ĳ��^9 Ĳ��]� ����]�      B   , ����`� ����aO ǖ��aO ǖ��`� ����`�      B   , ����`U ����`� �$��`� �$��`U ����`U      B   , �F��`U �F��`� ǖ��`� ǖ��`U �F��`U      B   , ����^� ����`U ǖ��`U ǖ��^� ����^�      B   , ����^9 ����^� �$��^� �$��^9 ����^9      B   , �F��^9 �F��^� ǖ��^� ǖ��^9 �F��^9      B   , ����]� ����^9 ǖ��^9 ǖ��]� ����]�      B   , ȸ��`� ȸ��aO �z��aO �z��`� ȸ��`�      B   , ȸ��`U ȸ��`� ���`� ���`U ȸ��`U      B   , �*��`U �*��`� �z��`� �z��`U �*��`U      B   , ȸ��^� ȸ��`U �z��`U �z��^� ȸ��^�      B   , ȸ��^9 ȸ��^� ���^� ���^9 ȸ��^9      B   , �*��^9 �*��^� �z��^� �z��^9 �*��^9      B   , ȸ��]� ȸ��^9 �z��^9 �z��]� ȸ��]�      B   , ˜��`� ˜��aO �^��aO �^��`� ˜��`�      B   , ˜��`U ˜��`� ����`� ����`U ˜��`U      B   , ���`U ���`� �^��`� �^��`U ���`U      B   , ˜��^� ˜��`U �^��`U �^��^� ˜��^�      B   , ˜��^9 ˜��^� ����^� ����^9 ˜��^9      B   , ���^9 ���^� �^��^� �^��^9 ���^9      B   , ˜��]� ˜��^9 �^��^9 �^��]� ˜��]�      B  , , �  ') �  '� 9  '� 9  ') �  ')      B  , , �  % �  %� 9  %� 9  % �  %      B  , , ��  2� ��  3� �b  3� �b  2� ��  2�      B  , , ��  1� ��  2A �b  2A �b  1� ��  1�      B  , , ��  0C ��  0� �b  0� �b  0C ��  0C      B  , , ��  .� ��  /� �b  /� �b  .� ��  .�      B  , , ��  -� ��  .E �b  .E �b  -� ��  -�      B  , , ��  ,G ��  ,� �b  ,� �b  ,G ��  ,G      B  , , ��  *� ��  +� �b  +� �b  *� ��  *�      B  , , ��  )� ��  *I �b  *I �b  )� ��  )�      B  , , ��  "� ��  #A �b  #A �b  "� ��  "�      B  , , ��  !C ��  !� �b  !� �b  !C ��  !C      B  , , ��  � ��   � �b   � �b  � ��  �      B  , , ��  � ��  E �b  E �b  � ��  �      B  , , ��  G ��  � �b  � �b  G ��  G      B  , , ��  � ��  � �b  � �b  � ��  �      B  , , ��  � ��  I �b  I �b  � ��  �      B  , , ��  K ��  � �b  � �b  K ��  K      B  , , ��  1� ��  2A �n  2A �n  1� ��  1�      B  , , ��  0C ��  0� �n  0� �n  0C ��  0C      B  , , ��  .� ��  /� �n  /� �n  .� ��  .�      B  , , ��  -� ��  .E �n  .E �n  -� ��  -�      B  , , ��  ,G ��  ,� �n  ,� �n  ,G ��  ,G      B  , , ��  *� ��  +� �n  +� �n  *� ��  *�      B  , , ��  )� ��  *I �n  *I �n  )� ��  )�      B  , , ��  % ��  %� ��  %� ��  % ��  %      B  , , �-  % �-  %� ��  %� ��  % �-  %      B  , , �{  % �{  %� �%  %� �%  % �{  %      B  , , ��  % ��  %� �s  %� �s  % ��  %      B  , , �  % �  %� ��  %� ��  % �  %      B  , , �e  % �e  %� �  %� �  % �e  %      B  , , ��  % ��  %� �]  %� �]  % ��  %      B  , , �  % �  %� ��  %� ��  % �  %      B  , , �O  % �O  %� ��  %� ��  % �O  %      B  , , ��  % ��  %� �G  %� �G  % ��  %      B  , , ��  % ��  %� ��  %� ��  % ��  %      B  , , �9  % �9  %� ��  %� ��  % �9  %      B  , , ��  % ��  %� �1  %� �1  % ��  %      B  , , ��  % ��  %� �  %� �  % ��  %      B  , , �#  % �#  %� ��  %� ��  % �#  %      B  , , �q  % �q  %� �  %� �  % �q  %      B  , , ƿ  % ƿ  %� �i  %� �i  % ƿ  %      B  , , �  % �  %� ɷ  %� ɷ  % �  %      B  , , �[  % �[  %� �  %� �  % �[  %      B  , , ͩ  % ͩ  %� �S  %� �S  % ͩ  %      B  , , ��  "� ��  #A �n  #A �n  "� ��  "�      B  , , ��  !C ��  !� �n  !� �n  !C ��  !C      B  , , ��  2� ��  3� �n  3� �n  2� ��  2�      B  , , ��  � ��   � �n   � �n  � ��  �      B  , , ��  � ��  E �n  E �n  � ��  �      B  , , ��  G ��  � �n  � �n  G ��  G      B  , , ��  � ��  � �n  � �n  � ��  �      B  , , ��  � ��  I �n  I �n  � ��  �      B  , , ��  K ��  � �n  � �n  K ��  K      B  , , ̂  .� ̂  /� �,  /� �,  .� ̂  .�      B  , , ��  .� ��  /� �z  /� �z  .� ��  .�      B  , , ̂  2� ̂  3� �,  3� �,  2� ̂  2�      B  , , �  -� �  .E ��  .E ��  -� �  -�      B  , , �`  -� �`  .E �
  .E �
  -� �`  -�      B  , , ��  -� ��  .E �X  .E �X  -� ��  -�      B  , , ��  -� ��  .E ��  .E ��  -� ��  -�      B  , , �J  -� �J  .E ��  .E ��  -� �J  -�      B  , , Ř  -� Ř  .E �B  .E �B  -� Ř  -�      B  , , ��  -� ��  .E Ȑ  .E Ȑ  -� ��  -�      B  , , �4  -� �4  .E ��  .E ��  -� �4  -�      B  , , ̂  -� ̂  .E �,  .E �,  -� ̂  -�      B  , , ��  -� ��  .E �z  .E �z  -� ��  -�      B  , , ��  2� ��  3� �z  3� �z  2� ��  2�      B  , , �  ,G �  ,� ��  ,� ��  ,G �  ,G      B  , , �`  ,G �`  ,� �
  ,� �
  ,G �`  ,G      B  , , ��  ,G ��  ,� �X  ,� �X  ,G ��  ,G      B  , , ��  ,G ��  ,� ��  ,� ��  ,G ��  ,G      B  , , �J  ,G �J  ,� ��  ,� ��  ,G �J  ,G      B  , , Ř  ,G Ř  ,� �B  ,� �B  ,G Ř  ,G      B  , , ��  ,G ��  ,� Ȑ  ,� Ȑ  ,G ��  ,G      B  , , �4  ,G �4  ,� ��  ,� ��  ,G �4  ,G      B  , , ̂  ,G ̂  ,� �,  ,� �,  ,G ̂  ,G      B  , , ��  ,G ��  ,� �z  ,� �z  ,G ��  ,G      B  , , Ř  2� Ř  3� �B  3� �B  2� Ř  2�      B  , , �  *� �  +� ��  +� ��  *� �  *�      B  , , �`  *� �`  +� �
  +� �
  *� �`  *�      B  , , ��  *� ��  +� �X  +� �X  *� ��  *�      B  , , ��  *� ��  +� ��  +� ��  *� ��  *�      B  , , �J  *� �J  +� ��  +� ��  *� �J  *�      B  , , Ř  *� Ř  +� �B  +� �B  *� Ř  *�      B  , , ��  *� ��  +� Ȑ  +� Ȑ  *� ��  *�      B  , , �4  *� �4  +� ��  +� ��  *� �4  *�      B  , , ̂  *� ̂  +� �,  +� �,  *� ̂  *�      B  , , ��  *� ��  +� �z  +� �z  *� ��  *�      B  , , �  1� �  2A ��  2A ��  1� �  1�      B  , , �  )� �  *I ��  *I ��  )� �  )�      B  , , �`  )� �`  *I �
  *I �
  )� �`  )�      B  , , ��  )� ��  *I �X  *I �X  )� ��  )�      B  , , ��  )� ��  *I ��  *I ��  )� ��  )�      B  , , �J  )� �J  *I ��  *I ��  )� �J  )�      B  , , Ř  )� Ř  *I �B  *I �B  )� Ř  )�      B  , , ��  )� ��  *I Ȑ  *I Ȑ  )� ��  )�      B  , , �4  )� �4  *I ��  *I ��  )� �4  )�      B  , , ̂  )� ̂  *I �,  *I �,  )� ̂  )�      B  , , ��  )� ��  *I �z  *I �z  )� ��  )�      B  , , ��  ') ��  '� ��  '� ��  ') ��  ')      B  , , �9  ') �9  '� ��  '� ��  ') �9  ')      B  , , ��  ') ��  '� �1  '� �1  ') ��  ')      B  , , ��  ') ��  '� �  '� �  ') ��  ')      B  , , �#  ') �#  '� ��  '� ��  ') �#  ')      B  , , �q  ') �q  '� �  '� �  ') �q  ')      B  , , ƿ  ') ƿ  '� �i  '� �i  ') ƿ  ')      B  , , �  ') �  '� ɷ  '� ɷ  ') �  ')      B  , , �[  ') �[  '� �  '� �  ') �[  ')      B  , , ͩ  ') ͩ  '� �S  '� �S  ') ͩ  ')      B  , , �`  1� �`  2A �
  2A �
  1� �`  1�      B  , , ��  1� ��  2A �X  2A �X  1� ��  1�      B  , , ��  1� ��  2A ��  2A ��  1� ��  1�      B  , , �J  1� �J  2A ��  2A ��  1� �J  1�      B  , , Ř  1� Ř  2A �B  2A �B  1� Ř  1�      B  , , ��  1� ��  2A Ȑ  2A Ȑ  1� ��  1�      B  , , �4  1� �4  2A ��  2A ��  1� �4  1�      B  , , ̂  1� ̂  2A �,  2A �,  1� ̂  1�      B  , , ��  1� ��  2A �z  2A �z  1� ��  1�      B  , , ��  2� ��  3� Ȑ  3� Ȑ  2� ��  2�      B  , , �  0C �  0� ��  0� ��  0C �  0C      B  , , �`  0C �`  0� �
  0� �
  0C �`  0C      B  , , ��  0C ��  0� �X  0� �X  0C ��  0C      B  , , ��  0C ��  0� ��  0� ��  0C ��  0C      B  , , �J  0C �J  0� ��  0� ��  0C �J  0C      B  , , Ř  0C Ř  0� �B  0� �B  0C Ř  0C      B  , , ��  0C ��  0� Ȑ  0� Ȑ  0C ��  0C      B  , , �4  0C �4  0� ��  0� ��  0C �4  0C      B  , , ̂  0C ̂  0� �,  0� �,  0C ̂  0C      B  , , ��  0C ��  0� �z  0� �z  0C ��  0C      B  , , �4  2� �4  3� ��  3� ��  2� �4  2�      B  , , �  .� �  /� ��  /� ��  .� �  .�      B  , , �`  .� �`  /� �
  /� �
  .� �`  .�      B  , , ��  .� ��  /� �X  /� �X  .� ��  .�      B  , , �  2� �  3� ��  3� ��  2� �  2�      B  , , ��  .� ��  /� ��  /� ��  .� ��  .�      B  , , �`  2� �`  3� �
  3� �
  2� �`  2�      B  , , �J  .� �J  /� ��  /� ��  .� �J  .�      B  , , ��  2� ��  3� �X  3� �X  2� ��  2�      B  , , Ř  .� Ř  /� �B  /� �B  .� Ř  .�      B  , , ��  2� ��  3� ��  3� ��  2� ��  2�      B  , , ��  .� ��  /� Ȑ  /� Ȑ  .� ��  .�      B  , , �J  2� �J  3� ��  3� ��  2� �J  2�      B  , , �4  .� �4  /� ��  /� ��  .� �4  .�      B  , , �  1� �  2A ��  2A ��  1� �  1�      B  , , �T  1� �T  2A ��  2A ��  1� �T  1�      B  , , ��  2� ��  3� ��  3� ��  2� ��  2�      B  , , �  -� �  .E ��  .E ��  -� �  -�      B  , , �T  -� �T  .E ��  .E ��  -� �T  -�      B  , , ��  2� ��  3� ��  3� ��  2� ��  2�      B  , , �  )� �  *I ��  *I ��  )� �  )�      B  , , �T  )� �T  *I ��  *I ��  )� �T  )�      B  , , ��  )� ��  *I �L  *I �L  )� ��  )�      B  , , ��  )� ��  *I ��  *I ��  )� ��  )�      B  , , �>  )� �>  *I ��  *I ��  )� �>  )�      B  , , ��  )� ��  *I �6  *I �6  )� ��  )�      B  , , ��  )� ��  *I ��  *I ��  )� ��  )�      B  , , �(  )� �(  *I ��  *I ��  )� �(  )�      B  , , �v  )� �v  *I �   *I �   )� �v  )�      B  , , ��  -� ��  .E �L  .E �L  -� ��  -�      B  , , ��  -� ��  .E ��  .E ��  -� ��  -�      B  , , �>  -� �>  .E ��  .E ��  -� �>  -�      B  , , ��  -� ��  .E �6  .E �6  -� ��  -�      B  , , ��  -� ��  .E ��  .E ��  -� ��  -�      B  , , �(  -� �(  .E ��  .E ��  -� �(  -�      B  , , �v  -� �v  .E �   .E �   -� �v  -�      B  , , ��  1� ��  2A �L  2A �L  1� ��  1�      B  , , ��  1� ��  2A ��  2A ��  1� ��  1�      B  , , �>  1� �>  2A ��  2A ��  1� �>  1�      B  , , ��  1� ��  2A �6  2A �6  1� ��  1�      B  , , ��  ') ��  '� ��  '� ��  ') ��  ')      B  , , �-  ') �-  '� ��  '� ��  ') �-  ')      B  , , �{  ') �{  '� �%  '� �%  ') �{  ')      B  , , ��  ') ��  '� �s  '� �s  ') ��  ')      B  , , �  ') �  '� ��  '� ��  ') �  ')      B  , , �e  ') �e  '� �  '� �  ') �e  ')      B  , , ��  ') ��  '� �]  '� �]  ') ��  ')      B  , , �  ') �  '� ��  '� ��  ') �  ')      B  , , �O  ') �O  '� ��  '� ��  ') �O  ')      B  , , ��  ') ��  '� �G  '� �G  ') ��  ')      B  , , ��  1� ��  2A ��  2A ��  1� ��  1�      B  , , �(  1� �(  2A ��  2A ��  1� �(  1�      B  , , �v  1� �v  2A �   2A �   1� �v  1�      B  , , �  2� �  3� ��  3� ��  2� �  2�      B  , , �T  2� �T  3� ��  3� ��  2� �T  2�      B  , , ��  2� ��  3� �L  3� �L  2� ��  2�      B  , , �  .� �  /� ��  /� ��  .� �  .�      B  , , �>  2� �>  3� ��  3� ��  2� �>  2�      B  , , �  ,G �  ,� ��  ,� ��  ,G �  ,G      B  , , �T  ,G �T  ,� ��  ,� ��  ,G �T  ,G      B  , , ��  ,G ��  ,� �L  ,� �L  ,G ��  ,G      B  , , ��  ,G ��  ,� ��  ,� ��  ,G ��  ,G      B  , , �>  ,G �>  ,� ��  ,� ��  ,G �>  ,G      B  , , ��  ,G ��  ,� �6  ,� �6  ,G ��  ,G      B  , , ��  ,G ��  ,� ��  ,� ��  ,G ��  ,G      B  , , �(  ,G �(  ,� ��  ,� ��  ,G �(  ,G      B  , , �v  ,G �v  ,� �   ,� �   ,G �v  ,G      B  , , �T  .� �T  /� ��  /� ��  .� �T  .�      B  , , ��  .� ��  /� �L  /� �L  .� ��  .�      B  , , ��  .� ��  /� ��  /� ��  .� ��  .�      B  , , �>  .� �>  /� ��  /� ��  .� �>  .�      B  , , ��  .� ��  /� �6  /� �6  .� ��  .�      B  , , ��  .� ��  /� ��  /� ��  .� ��  .�      B  , , �(  .� �(  /� ��  /� ��  .� �(  .�      B  , , �v  .� �v  /� �   /� �   .� �v  .�      B  , , �  0C �  0� ��  0� ��  0C �  0C      B  , , �T  0C �T  0� ��  0� ��  0C �T  0C      B  , , ��  0C ��  0� �L  0� �L  0C ��  0C      B  , , ��  2� ��  3� �6  3� �6  2� ��  2�      B  , , �  *� �  +� ��  +� ��  *� �  *�      B  , , �(  2� �(  3� ��  3� ��  2� �(  2�      B  , , �T  *� �T  +� ��  +� ��  *� �T  *�      B  , , �v  2� �v  3� �   3� �   2� �v  2�      B  , , ��  *� ��  +� �L  +� �L  *� ��  *�      B  , , ��  *� ��  +� ��  +� ��  *� ��  *�      B  , , �>  *� �>  +� ��  +� ��  *� �>  *�      B  , , ��  *� ��  +� �6  +� �6  *� ��  *�      B  , , ��  *� ��  +� ��  +� ��  *� ��  *�      B  , , �(  *� �(  +� ��  +� ��  *� �(  *�      B  , , �v  *� �v  +� �   +� �   *� �v  *�      B  , , ��  0C ��  0� ��  0� ��  0C ��  0C      B  , , �>  0C �>  0� ��  0� ��  0C �>  0C      B  , , ��  0C ��  0� �6  0� �6  0C ��  0C      B  , , ��  0C ��  0� ��  0� ��  0C ��  0C      B  , , �(  0C �(  0� ��  0� ��  0C �(  0C      B  , , �v  0C �v  0� �   0� �   0C �v  0C      B  , , �>  !C �>  !� ��  !� ��  !C �>  !C      B  , , ��  !C ��  !� �6  !� �6  !C ��  !C      B  , , ��  !C ��  !� ��  !� ��  !C ��  !C      B  , , �(  !C �(  !� ��  !� ��  !C �(  !C      B  , , �v  !C �v  !� �   !� �   !C �v  !C      B  , , ��  "� ��  #A �L  #A �L  "� ��  "�      B  , , ��  "� ��  #A ��  #A ��  "� ��  "�      B  , , �  � �   � ��   � ��  � �  �      B  , , �T  � �T   � ��   � ��  � �T  �      B  , , ��  � ��   � �L   � �L  � ��  �      B  , , ��  � ��   � ��   � ��  � ��  �      B  , , �>  � �>   � ��   � ��  � �>  �      B  , , ��  � ��   � �6   � �6  � ��  �      B  , , ��  � ��   � ��   � ��  � ��  �      B  , , �(  � �(   � ��   � ��  � �(  �      B  , , �v  � �v   � �    � �   � �v  �      B  , , �>  "� �>  #A ��  #A ��  "� �>  "�      B  , , ��  "� ��  #A �6  #A �6  "� ��  "�      B  , , �  � �  E ��  E ��  � �  �      B  , , �T  � �T  E ��  E ��  � �T  �      B  , , ��  � ��  E �L  E �L  � ��  �      B  , , ��  � ��  E ��  E ��  � ��  �      B  , , �>  � �>  E ��  E ��  � �>  �      B  , , ��  � ��  E �6  E �6  � ��  �      B  , , ��  � ��  E ��  E ��  � ��  �      B  , , �(  � �(  E ��  E ��  � �(  �      B  , , �v  � �v  E �   E �   � �v  �      B  , , ��  "� ��  #A ��  #A ��  "� ��  "�      B  , , �(  "� �(  #A ��  #A ��  "� �(  "�      B  , , �  G �  � ��  � ��  G �  G      B  , , �T  G �T  � ��  � ��  G �T  G      B  , , ��  G ��  � �L  � �L  G ��  G      B  , , ��  G ��  � ��  � ��  G ��  G      B  , , �>  G �>  � ��  � ��  G �>  G      B  , , ��  G ��  � �6  � �6  G ��  G      B  , , ��  G ��  � ��  � ��  G ��  G      B  , , �(  G �(  � ��  � ��  G �(  G      B  , , �v  G �v  � �   � �   G �v  G      B  , , �v  "� �v  #A �   #A �   "� �v  "�      B  , , �  "� �  #A ��  #A ��  "� �  "�      B  , , �  � �  � ��  � ��  � �  �      B  , , �T  � �T  � ��  � ��  � �T  �      B  , , ��  � ��  � �L  � �L  � ��  �      B  , , ��  � ��  � ��  � ��  � ��  �      B  , , �>  � �>  � ��  � ��  � �>  �      B  , , ��  � ��  � �6  � �6  � ��  �      B  , , ��  � ��  � ��  � ��  � ��  �      B  , , �(  � �(  � ��  � ��  � �(  �      B  , , �v  � �v  � �   � �   � �v  �      B  , , �T  "� �T  #A ��  #A ��  "� �T  "�      B  , , �  !C �  !� ��  !� ��  !C �  !C      B  , , �  � �  I ��  I ��  � �  �      B  , , �T  � �T  I ��  I ��  � �T  �      B  , , ��  � ��  I �L  I �L  � ��  �      B  , , ��  � ��  I ��  I ��  � ��  �      B  , , �>  � �>  I ��  I ��  � �>  �      B  , , ��  � ��  I �6  I �6  � ��  �      B  , , ��  � ��  I ��  I ��  � ��  �      B  , , �(  � �(  I ��  I ��  � �(  �      B  , , �v  � �v  I �   I �   � �v  �      B  , , �T  !C �T  !� ��  !� ��  !C �T  !C      B  , , ��  !C ��  !� �L  !� �L  !C ��  !C      B  , , �  K �  � ��  � ��  K �  K      B  , , �T  K �T  � ��  � ��  K �T  K      B  , , ��  K ��  � �L  � �L  K ��  K      B  , , ��  K ��  � ��  � ��  K ��  K      B  , , �>  K �>  � ��  � ��  K �>  K      B  , , ��  K ��  � �6  � �6  K ��  K      B  , , ��  K ��  � ��  � ��  K ��  K      B  , , �(  K �(  � ��  � ��  K �(  K      B  , , �v  K �v  � �   � �   K �v  K      B  , , ��  !C ��  !� ��  !� ��  !C ��  !C      B  , , �4  "� �4  #A ��  #A ��  "� �4  "�      B  , , ̂  "� ̂  #A �,  #A �,  "� ̂  "�      B  , , ��  "� ��  #A �z  #A �z  "� ��  "�      B  , , �  "� �  #A ��  #A ��  "� �  "�      B  , , �  !C �  !� ��  !� ��  !C �  !C      B  , , �  � �   � ��   � ��  � �  �      B  , , �`  � �`   � �
   � �
  � �`  �      B  , , �  G �  � ��  � ��  G �  G      B  , , �`  G �`  � �
  � �
  G �`  G      B  , , ��  G ��  � �X  � �X  G ��  G      B  , , ��  G ��  � ��  � ��  G ��  G      B  , , �J  G �J  � ��  � ��  G �J  G      B  , , Ř  G Ř  � �B  � �B  G Ř  G      B  , , ��  G ��  � Ȑ  � Ȑ  G ��  G      B  , , �4  G �4  � ��  � ��  G �4  G      B  , , ̂  G ̂  � �,  � �,  G ̂  G      B  , , ��  G ��  � �z  � �z  G ��  G      B  , , ��  � ��   � �X   � �X  � ��  �      B  , , ��  � ��   � ��   � ��  � ��  �      B  , , �J  � �J   � ��   � ��  � �J  �      B  , , Ř  � Ř   � �B   � �B  � Ř  �      B  , , ��  � ��   � Ȑ   � Ȑ  � ��  �      B  , , �4  � �4   � ��   � ��  � �4  �      B  , , ̂  � ̂   � �,   � �,  � ̂  �      B  , , ��  � ��   � �z   � �z  � ��  �      B  , , �`  !C �`  !� �
  !� �
  !C �`  !C      B  , , ��  !C ��  !� �X  !� �X  !C ��  !C      B  , , ��  !C ��  !� ��  !� ��  !C ��  !C      B  , , �  � �  � ��  � ��  � �  �      B  , , �`  � �`  � �
  � �
  � �`  �      B  , , ��  � ��  � �X  � �X  � ��  �      B  , , ��  � ��  � ��  � ��  � ��  �      B  , , �J  � �J  � ��  � ��  � �J  �      B  , , Ř  � Ř  � �B  � �B  � Ř  �      B  , , ��  � ��  � Ȑ  � Ȑ  � ��  �      B  , , �4  � �4  � ��  � ��  � �4  �      B  , , ̂  � ̂  � �,  � �,  � ̂  �      B  , , ��  � ��  � �z  � �z  � ��  �      B  , , �J  !C �J  !� ��  !� ��  !C �J  !C      B  , , Ř  !C Ř  !� �B  !� �B  !C Ř  !C      B  , , ��  !C ��  !� Ȑ  !� Ȑ  !C ��  !C      B  , , �4  !C �4  !� ��  !� ��  !C �4  !C      B  , , ̂  !C ̂  !� �,  !� �,  !C ̂  !C      B  , , ��  !C ��  !� �z  !� �z  !C ��  !C      B  , , �`  "� �`  #A �
  #A �
  "� �`  "�      B  , , ��  "� ��  #A �X  #A �X  "� ��  "�      B  , , �  � �  E ��  E ��  � �  �      B  , , �`  � �`  E �
  E �
  � �`  �      B  , , ��  � ��  E �X  E �X  � ��  �      B  , , �  � �  I ��  I ��  � �  �      B  , , �`  � �`  I �
  I �
  � �`  �      B  , , ��  � ��  I �X  I �X  � ��  �      B  , , ��  � ��  I ��  I ��  � ��  �      B  , , �J  � �J  I ��  I ��  � �J  �      B  , , Ř  � Ř  I �B  I �B  � Ř  �      B  , , ��  � ��  I Ȑ  I Ȑ  � ��  �      B  , , �4  � �4  I ��  I ��  � �4  �      B  , , ̂  � ̂  I �,  I �,  � ̂  �      B  , , ��  � ��  I �z  I �z  � ��  �      B  , , ��  � ��  E ��  E ��  � ��  �      B  , , �J  � �J  E ��  E ��  � �J  �      B  , , Ř  � Ř  E �B  E �B  � Ř  �      B  , , ��  � ��  E Ȑ  E Ȑ  � ��  �      B  , , �4  � �4  E ��  E ��  � �4  �      B  , , ̂  � ̂  E �,  E �,  � ̂  �      B  , , ��  � ��  E �z  E �z  � ��  �      B  , , ��  "� ��  #A ��  #A ��  "� ��  "�      B  , , �J  "� �J  #A ��  #A ��  "� �J  "�      B  , , Ř  "� Ř  #A �B  #A �B  "� Ř  "�      B  , , ��  "� ��  #A Ȑ  #A Ȑ  "� ��  "�      B  , , �  K �  � ��  � ��  K �  K      B  , , �`  K �`  � �
  � �
  K �`  K      B  , , ��  K ��  � �X  � �X  K ��  K      B  , , ��  K ��  � ��  � ��  K ��  K      B  , , �J  K �J  � ��  � ��  K �J  K      B  , , Ř  K Ř  � �B  � �B  K Ř  K      B  , , ��  K ��  � Ȑ  � Ȑ  K ��  K      B  , , �4  K �4  � ��  � ��  K �4  K      B  , , ̂  K ̂  � �,  � �,  K ̂  K      B  , , ��  K ��  � �z  � �z  K ��  K      B  , , s�  % s�  %� t�  %� t�  % s�  %      B  , , v8  % v8  %� v�  %� v�  % v8  %      B  , , x�  % x�  %� y0  %� y0  % x�  %      B  , , z�  % z�  %� {~  %� {~  % z�  %      B  , , }"  % }"  %� }�  %� }�  % }"  %      B  , , ��  % ��  %� �Q  %� �Q  % ��  %      B  , , ��  % ��  %� ��  %� ��  % ��  %      B  , , �C  % �C  %� ��  %� ��  % �C  %      B  , , ��  % ��  %� �;  %� �;  % ��  %      B  , , �j  1� �j  2A �  2A �  1� �j  1�      B  , , �j  )� �j  *I �  *I �  )� �j  )�      B  , , �j  0C �j  0� �  0� �  0C �j  0C      B  , , �j  -� �j  .E �  .E �  -� �j  -�      B  , , �j  .� �j  /� �  /� �  .� �j  .�      B  , , ��  ') ��  '� �Q  '� �Q  ') ��  ')      B  , , ��  ') ��  '� ��  '� ��  ') ��  ')      B  , , �C  ') �C  '� ��  '� ��  ') �C  ')      B  , , ��  ') ��  '� �;  '� �;  ') ��  ')      B  , , �j  *� �j  +� �  +� �  *� �j  *�      B  , , �j  2� �j  3� �  3� �  2� �j  2�      B  , , �j  ,G �j  ,� �  ,� �  ,G �j  ,G      B  , , {�  .� {�  /� |�  /� |�  .� {�  .�      B  , , ~I  .� ~I  /� ~�  /� ~�  .� ~I  .�      B  , , r�  0C r�  0� sm  0� sm  0C r�  0C      B  , , s�  ') s�  '� t�  '� t�  ') s�  ')      B  , , v8  ') v8  '� v�  '� v�  ') v8  ')      B  , , x�  ') x�  '� y0  '� y0  ') x�  ')      B  , , z�  ') z�  '� {~  '� {~  ') z�  ')      B  , , }"  ') }"  '� }�  '� }�  ') }"  ')      B  , , u  0C u  0� u�  0� u�  0C u  0C      B  , , w_  0C w_  0� x	  0� x	  0C w_  0C      B  , , y�  0C y�  0� zW  0� zW  0C y�  0C      B  , , {�  0C {�  0� |�  0� |�  0C {�  0C      B  , , r�  *� r�  +� sm  +� sm  *� r�  *�      B  , , u  *� u  +� u�  +� u�  *� u  *�      B  , , w_  *� w_  +� x	  +� x	  *� w_  *�      B  , , y�  *� y�  +� zW  +� zW  *� y�  *�      B  , , {�  *� {�  +� |�  +� |�  *� {�  *�      B  , , ~I  *� ~I  +� ~�  +� ~�  *� ~I  *�      B  , , ~I  0C ~I  0� ~�  0� ~�  0C ~I  0C      B  , , r�  1� r�  2A sm  2A sm  1� r�  1�      B  , , u  1� u  2A u�  2A u�  1� u  1�      B  , , w_  1� w_  2A x	  2A x	  1� w_  1�      B  , , y�  1� y�  2A zW  2A zW  1� y�  1�      B  , , {�  1� {�  2A |�  2A |�  1� {�  1�      B  , , ~I  1� ~I  2A ~�  2A ~�  1� ~I  1�      B  , , ~I  )� ~I  *I ~�  *I ~�  )� ~I  )�      B  , , r�  2� r�  3� sm  3� sm  2� r�  2�      B  , , u  2� u  3� u�  3� u�  2� u  2�      B  , , w_  2� w_  3� x	  3� x	  2� w_  2�      B  , , y�  2� y�  3� zW  3� zW  2� y�  2�      B  , , {�  2� {�  3� |�  3� |�  2� {�  2�      B  , , ~I  2� ~I  3� ~�  3� ~�  2� ~I  2�      B  , , r�  -� r�  .E sm  .E sm  -� r�  -�      B  , , u  -� u  .E u�  .E u�  -� u  -�      B  , , w_  -� w_  .E x	  .E x	  -� w_  -�      B  , , y�  -� y�  .E zW  .E zW  -� y�  -�      B  , , {�  -� {�  .E |�  .E |�  -� {�  -�      B  , , ~I  -� ~I  .E ~�  .E ~�  -� ~I  -�      B  , , {�  )� {�  *I |�  *I |�  )� {�  )�      B  , , r�  .� r�  /� sm  /� sm  .� r�  .�      B  , , u  .� u  /� u�  /� u�  .� u  .�      B  , , w_  .� w_  /� x	  /� x	  .� w_  .�      B  , , r�  ,G r�  ,� sm  ,� sm  ,G r�  ,G      B  , , u  ,G u  ,� u�  ,� u�  ,G u  ,G      B  , , w_  ,G w_  ,� x	  ,� x	  ,G w_  ,G      B  , , y�  ,G y�  ,� zW  ,� zW  ,G y�  ,G      B  , , {�  ,G {�  ,� |�  ,� |�  ,G {�  ,G      B  , , ~I  ,G ~I  ,� ~�  ,� ~�  ,G ~I  ,G      B  , , y�  .� y�  /� zW  /� zW  .� y�  .�      B  , , r�  )� r�  *I sm  *I sm  )� r�  )�      B  , , u  )� u  *I u�  *I u�  )� u  )�      B  , , w_  )� w_  *I x	  *I x	  )� w_  )�      B  , , y�  )� y�  *I zW  *I zW  )� y�  )�      B  , , {�  � {�  I |�  I |�  � {�  �      B  , , ~I  � ~I  I ~�  I ~�  � ~I  �      B  , , w_  � w_  � x	  � x	  � w_  �      B  , , y�  � y�  � zW  � zW  � y�  �      B  , , {�  � {�  � |�  � |�  � {�  �      B  , , ~I  � ~I  � ~�  � ~�  � ~I  �      B  , , r�  � r�   � sm   � sm  � r�  �      B  , , u  � u   � u�   � u�  � u  �      B  , , w_  � w_   � x	   � x	  � w_  �      B  , , y�  � y�   � zW   � zW  � y�  �      B  , , {�  � {�   � |�   � |�  � {�  �      B  , , ~I  � ~I   � ~�   � ~�  � ~I  �      B  , , y�  !C y�  !� zW  !� zW  !C y�  !C      B  , , {�  !C {�  !� |�  !� |�  !C {�  !C      B  , , ~I  !C ~I  !� ~�  !� ~�  !C ~I  !C      B  , , r�  G r�  � sm  � sm  G r�  G      B  , , u  G u  � u�  � u�  G u  G      B  , , w_  G w_  � x	  � x	  G w_  G      B  , , y�  G y�  � zW  � zW  G y�  G      B  , , {�  G {�  � |�  � |�  G {�  G      B  , , ~I  G ~I  � ~�  � ~�  G ~I  G      B  , , y�  "� y�  #A zW  #A zW  "� y�  "�      B  , , r�  K r�  � sm  � sm  K r�  K      B  , , u  K u  � u�  � u�  K u  K      B  , , w_  K w_  � x	  � x	  K w_  K      B  , , y�  K y�  � zW  � zW  K y�  K      B  , , {�  K {�  � |�  � |�  K {�  K      B  , , ~I  K ~I  � ~�  � ~�  K ~I  K      B  , , {�  "� {�  #A |�  #A |�  "� {�  "�      B  , , ~I  "� ~I  #A ~�  #A ~�  "� ~I  "�      B  , , r�  "� r�  #A sm  #A sm  "� r�  "�      B  , , u  "� u  #A u�  #A u�  "� u  "�      B  , , w_  "� w_  #A x	  #A x	  "� w_  "�      B  , , r�  !C r�  !� sm  !� sm  !C r�  !C      B  , , u  !C u  !� u�  !� u�  !C u  !C      B  , , w_  !C w_  !� x	  !� x	  !C w_  !C      B  , , r�  � r�  � sm  � sm  � r�  �      B  , , u  � u  � u�  � u�  � u  �      B  , , r�  � r�  I sm  I sm  � r�  �      B  , , r�  � r�  E sm  E sm  � r�  �      B  , , u  � u  E u�  E u�  � u  �      B  , , w_  � w_  E x	  E x	  � w_  �      B  , , y�  � y�  E zW  E zW  � y�  �      B  , , {�  � {�  E |�  E |�  � {�  �      B  , , ~I  � ~I  E ~�  E ~�  � ~I  �      B  , , u  � u  I u�  I u�  � u  �      B  , , w_  � w_  I x	  I x	  � w_  �      B  , , y�  � y�  I zW  I zW  � y�  �      B  , , �j  K �j  � �  � �  K �j  K      B  , , �j  � �j  I �  I �  � �j  �      B  , , �j  � �j   � �   � �  � �j  �      B  , , �j  !C �j  !� �  !� �  !C �j  !C      B  , , �j  � �j  E �  E �  � �j  �      B  , , �j  G �j  � �  � �  G �j  G      B  , , �j  "� �j  #A �  #A �  "� �j  "�      B  , , �j  � �j  � �  � �  � �j  �      B  , , H   % H   %� H�  %� H�  % H   %      B  , , Jn  % Jn  %� K  %� K  % Jn  %      B  , , L�  % L�  %� Mf  %� Mf  % L�  %      B  , , O
  % O
  %� O�  %� O�  % O
  %      B  , , QX  % QX  %� R  %� R  % QX  %      B  , , S�  % S�  %� TP  %� TP  % S�  %      B  , , U�  % U�  %� V�  %� V�  % U�  %      B  , , XB  % XB  %� X�  %� X�  % XB  %      B  , , Z�  % Z�  %� [:  %� [:  % Z�  %      B  , , \�  % \�  %� ]�  %� ]�  % \�  %      B  , , _,  % _,  %� _�  %� _�  % _,  %      B  , , az  % az  %� b$  %� b$  % az  %      B  , , c�  % c�  %� dr  %� dr  % c�  %      B  , , f  % f  %� f�  %� f�  % f  %      B  , , hd  % hd  %� i  %� i  % hd  %      B  , , j�  % j�  %� k\  %� k\  % j�  %      B  , , m   % m   %� m�  %� m�  % m   %      B  , , oN  % oN  %� o�  %� o�  % oN  %      B  , , q�  % q�  %� rF  %� rF  % q�  %      B  , , [�  0C [�  0� \a  0� \a  0C [�  0C      B  , , ^  0C ^  0� ^�  0� ^�  0C ^  0C      B  , , `S  0C `S  0� `�  0� `�  0C `S  0C      B  , , b�  0C b�  0� cK  0� cK  0C b�  0C      B  , , d�  0C d�  0� e�  0� e�  0C d�  0C      B  , , g=  0C g=  0� g�  0� g�  0C g=  0C      B  , , i�  0C i�  0� j5  0� j5  0C i�  0C      B  , , k�  0C k�  0� l�  0� l�  0C k�  0C      B  , , n'  0C n'  0� n�  0� n�  0C n'  0C      B  , , pu  0C pu  0� q  0� q  0C pu  0C      B  , , [�  ,G [�  ,� \a  ,� \a  ,G [�  ,G      B  , , ^  ,G ^  ,� ^�  ,� ^�  ,G ^  ,G      B  , , `S  ,G `S  ,� `�  ,� `�  ,G `S  ,G      B  , , b�  ,G b�  ,� cK  ,� cK  ,G b�  ,G      B  , , d�  ,G d�  ,� e�  ,� e�  ,G d�  ,G      B  , , g=  ,G g=  ,� g�  ,� g�  ,G g=  ,G      B  , , i�  ,G i�  ,� j5  ,� j5  ,G i�  ,G      B  , , k�  ,G k�  ,� l�  ,� l�  ,G k�  ,G      B  , , n'  ,G n'  ,� n�  ,� n�  ,G n'  ,G      B  , , pu  ,G pu  ,� q  ,� q  ,G pu  ,G      B  , , [�  1� [�  2A \a  2A \a  1� [�  1�      B  , , ^  1� ^  2A ^�  2A ^�  1� ^  1�      B  , , `S  1� `S  2A `�  2A `�  1� `S  1�      B  , , b�  1� b�  2A cK  2A cK  1� b�  1�      B  , , d�  1� d�  2A e�  2A e�  1� d�  1�      B  , , g=  1� g=  2A g�  2A g�  1� g=  1�      B  , , i�  1� i�  2A j5  2A j5  1� i�  1�      B  , , k�  1� k�  2A l�  2A l�  1� k�  1�      B  , , n'  1� n'  2A n�  2A n�  1� n'  1�      B  , , pu  1� pu  2A q  2A q  1� pu  1�      B  , , [�  *� [�  +� \a  +� \a  *� [�  *�      B  , , ^  *� ^  +� ^�  +� ^�  *� ^  *�      B  , , `S  *� `S  +� `�  +� `�  *� `S  *�      B  , , b�  *� b�  +� cK  +� cK  *� b�  *�      B  , , d�  *� d�  +� e�  +� e�  *� d�  *�      B  , , g=  *� g=  +� g�  +� g�  *� g=  *�      B  , , i�  *� i�  +� j5  +� j5  *� i�  *�      B  , , k�  *� k�  +� l�  +� l�  *� k�  *�      B  , , n'  *� n'  +� n�  +� n�  *� n'  *�      B  , , pu  *� pu  +� q  +� q  *� pu  *�      B  , , [�  .� [�  /� \a  /� \a  .� [�  .�      B  , , ^  .� ^  /� ^�  /� ^�  .� ^  .�      B  , , `S  .� `S  /� `�  /� `�  .� `S  .�      B  , , b�  .� b�  /� cK  /� cK  .� b�  .�      B  , , d�  .� d�  /� e�  /� e�  .� d�  .�      B  , , g=  .� g=  /� g�  /� g�  .� g=  .�      B  , , i�  .� i�  /� j5  /� j5  .� i�  .�      B  , , k�  .� k�  /� l�  /� l�  .� k�  .�      B  , , n'  .� n'  /� n�  /� n�  .� n'  .�      B  , , pu  .� pu  /� q  /� q  .� pu  .�      B  , , [�  )� [�  *I \a  *I \a  )� [�  )�      B  , , ^  )� ^  *I ^�  *I ^�  )� ^  )�      B  , , `S  )� `S  *I `�  *I `�  )� `S  )�      B  , , b�  )� b�  *I cK  *I cK  )� b�  )�      B  , , d�  )� d�  *I e�  *I e�  )� d�  )�      B  , , g=  )� g=  *I g�  *I g�  )� g=  )�      B  , , i�  )� i�  *I j5  *I j5  )� i�  )�      B  , , k�  )� k�  *I l�  *I l�  )� k�  )�      B  , , n'  )� n'  *I n�  *I n�  )� n'  )�      B  , , pu  )� pu  *I q  *I q  )� pu  )�      B  , , [�  2� [�  3� \a  3� \a  2� [�  2�      B  , , ^  2� ^  3� ^�  3� ^�  2� ^  2�      B  , , `S  2� `S  3� `�  3� `�  2� `S  2�      B  , , b�  2� b�  3� cK  3� cK  2� b�  2�      B  , , d�  2� d�  3� e�  3� e�  2� d�  2�      B  , , g=  2� g=  3� g�  3� g�  2� g=  2�      B  , , i�  2� i�  3� j5  3� j5  2� i�  2�      B  , , k�  2� k�  3� l�  3� l�  2� k�  2�      B  , , n'  2� n'  3� n�  3� n�  2� n'  2�      B  , , pu  2� pu  3� q  3� q  2� pu  2�      B  , , \�  ') \�  '� ]�  '� ]�  ') \�  ')      B  , , _,  ') _,  '� _�  '� _�  ') _,  ')      B  , , az  ') az  '� b$  '� b$  ') az  ')      B  , , c�  ') c�  '� dr  '� dr  ') c�  ')      B  , , f  ') f  '� f�  '� f�  ') f  ')      B  , , hd  ') hd  '� i  '� i  ') hd  ')      B  , , j�  ') j�  '� k\  '� k\  ') j�  ')      B  , , m   ') m   '� m�  '� m�  ') m   ')      B  , , oN  ') oN  '� o�  '� o�  ') oN  ')      B  , , q�  ') q�  '� rF  '� rF  ') q�  ')      B  , , [�  -� [�  .E \a  .E \a  -� [�  -�      B  , , ^  -� ^  .E ^�  .E ^�  -� ^  -�      B  , , `S  -� `S  .E `�  .E `�  -� `S  -�      B  , , b�  -� b�  .E cK  .E cK  -� b�  -�      B  , , d�  -� d�  .E e�  .E e�  -� d�  -�      B  , , g=  -� g=  .E g�  .E g�  -� g=  -�      B  , , i�  -� i�  .E j5  .E j5  -� i�  -�      B  , , k�  -� k�  .E l�  .E l�  -� k�  -�      B  , , n'  -� n'  .E n�  .E n�  -� n'  -�      B  , , pu  -� pu  .E q  .E q  -� pu  -�      B  , , W  *� W  +� W�  +� W�  *� W  *�      B  , , Yi  *� Yi  +� Z  +� Z  *� Yi  *�      B  , , W  ,G W  ,� W�  ,� W�  ,G W  ,G      B  , , M�  1� M�  2A N�  2A N�  1� M�  1�      B  , , P1  1� P1  2A P�  2A P�  1� P1  1�      B  , , R  1� R  2A S)  2A S)  1� R  1�      B  , , T�  1� T�  2A Uw  2A Uw  1� T�  1�      B  , , W  1� W  2A W�  2A W�  1� W  1�      B  , , Yi  1� Yi  2A Z  2A Z  1� Yi  1�      B  , , W  2� W  3� W�  3� W�  2� W  2�      B  , , Yi  2� Yi  3� Z  3� Z  2� Yi  2�      B  , , Yi  ,G Yi  ,� Z  ,� Z  ,G Yi  ,G      B  , , P1  0C P1  0� P�  0� P�  0C P1  0C      B  , , R  0C R  0� S)  0� S)  0C R  0C      B  , , M�  .� M�  /� N�  /� N�  .� M�  .�      B  , , P1  .� P1  /� P�  /� P�  .� P1  .�      B  , , R  .� R  /� S)  /� S)  .� R  .�      B  , , T�  .� T�  /� Uw  /� Uw  .� T�  .�      B  , , W  .� W  /� W�  /� W�  .� W  .�      B  , , Yi  .� Yi  /� Z  /� Z  .� Yi  .�      B  , , T�  0C T�  0� Uw  0� Uw  0C T�  0C      B  , , H   ') H   '� H�  '� H�  ') H   ')      B  , , Jn  ') Jn  '� K  '� K  ') Jn  ')      B  , , L�  ') L�  '� Mf  '� Mf  ') L�  ')      B  , , O
  ') O
  '� O�  '� O�  ') O
  ')      B  , , QX  ') QX  '� R  '� R  ') QX  ')      B  , , S�  ') S�  '� TP  '� TP  ') S�  ')      B  , , U�  ') U�  '� V�  '� V�  ') U�  ')      B  , , XB  ') XB  '� X�  '� X�  ') XB  ')      B  , , Z�  ') Z�  '� [:  '� [:  ') Z�  ')      B  , , W  0C W  0� W�  0� W�  0C W  0C      B  , , Yi  0C Yi  0� Z  0� Z  0C Yi  0C      B  , , M�  ,G M�  ,� N�  ,� N�  ,G M�  ,G      B  , , P1  ,G P1  ,� P�  ,� P�  ,G P1  ,G      B  , , R  ,G R  ,� S)  ,� S)  ,G R  ,G      B  , , T�  ,G T�  ,� Uw  ,� Uw  ,G T�  ,G      B  , , M�  *� M�  +� N�  +� N�  *� M�  *�      B  , , P1  *� P1  +� P�  +� P�  *� P1  *�      B  , , R  *� R  +� S)  +� S)  *� R  *�      B  , , M�  2� M�  3� N�  3� N�  2� M�  2�      B  , , M�  -� M�  .E N�  .E N�  -� M�  -�      B  , , P1  -� P1  .E P�  .E P�  -� P1  -�      B  , , R  -� R  .E S)  .E S)  -� R  -�      B  , , T�  -� T�  .E Uw  .E Uw  -� T�  -�      B  , , W  -� W  .E W�  .E W�  -� W  -�      B  , , Yi  -� Yi  .E Z  .E Z  -� Yi  -�      B  , , P1  2� P1  3� P�  3� P�  2� P1  2�      B  , , R  2� R  3� S)  3� S)  2� R  2�      B  , , T�  2� T�  3� Uw  3� Uw  2� T�  2�      B  , , M�  )� M�  *I N�  *I N�  )� M�  )�      B  , , P1  )� P1  *I P�  *I P�  )� P1  )�      B  , , R  )� R  *I S)  *I S)  )� R  )�      B  , , T�  )� T�  *I Uw  *I Uw  )� T�  )�      B  , , W  )� W  *I W�  *I W�  )� W  )�      B  , , Yi  )� Yi  *I Z  *I Z  )� Yi  )�      B  , , T�  *� T�  +� Uw  +� Uw  *� T�  *�      B  , , M�  0C M�  0� N�  0� N�  0C M�  0C      B  , , W  G W  � W�  � W�  G W  G      B  , , M�  � M�  I N�  I N�  � M�  �      B  , , P1  � P1  I P�  I P�  � P1  �      B  , , R  � R  I S)  I S)  � R  �      B  , , T�  � T�  I Uw  I Uw  � T�  �      B  , , W  � W  I W�  I W�  � W  �      B  , , Yi  � Yi  I Z  I Z  � Yi  �      B  , , Yi  G Yi  � Z  � Z  G Yi  G      B  , , T�  !C T�  !� Uw  !� Uw  !C T�  !C      B  , , W  !C W  !� W�  !� W�  !C W  !C      B  , , Yi  !C Yi  !� Z  !� Z  !C Yi  !C      B  , , M�  � M�  E N�  E N�  � M�  �      B  , , P1  � P1  E P�  E P�  � P1  �      B  , , R  � R  E S)  E S)  � R  �      B  , , T�  � T�  E Uw  E Uw  � T�  �      B  , , W  � W  E W�  E W�  � W  �      B  , , Yi  � Yi  E Z  E Z  � Yi  �      B  , , Yi  "� Yi  #A Z  #A Z  "� Yi  "�      B  , , M�  "� M�  #A N�  #A N�  "� M�  "�      B  , , P1  "� P1  #A P�  #A P�  "� P1  "�      B  , , R  "� R  #A S)  #A S)  "� R  "�      B  , , T�  "� T�  #A Uw  #A Uw  "� T�  "�      B  , , W  "� W  #A W�  #A W�  "� W  "�      B  , , M�  !C M�  !� N�  !� N�  !C M�  !C      B  , , P1  !C P1  !� P�  !� P�  !C P1  !C      B  , , R  !C R  !� S)  !� S)  !C R  !C      B  , , M�  � M�   � N�   � N�  � M�  �      B  , , P1  � P1   � P�   � P�  � P1  �      B  , , R  � R   � S)   � S)  � R  �      B  , , T�  � T�   � Uw   � Uw  � T�  �      B  , , M�  K M�  � N�  � N�  K M�  K      B  , , P1  K P1  � P�  � P�  K P1  K      B  , , R  K R  � S)  � S)  K R  K      B  , , T�  K T�  � Uw  � Uw  K T�  K      B  , , W  K W  � W�  � W�  K W  K      B  , , Yi  K Yi  � Z  � Z  K Yi  K      B  , , W  � W   � W�   � W�  � W  �      B  , , Yi  � Yi   � Z   � Z  � Yi  �      B  , , M�  G M�  � N�  � N�  G M�  G      B  , , P1  G P1  � P�  � P�  G P1  G      B  , , R  G R  � S)  � S)  G R  G      B  , , T�  G T�  � Uw  � Uw  G T�  G      B  , , M�  � M�  � N�  � N�  � M�  �      B  , , P1  � P1  � P�  � P�  � P1  �      B  , , R  � R  � S)  � S)  � R  �      B  , , T�  � T�  � Uw  � Uw  � T�  �      B  , , W  � W  � W�  � W�  � W  �      B  , , Yi  � Yi  � Z  � Z  � Yi  �      B  , , d�  "� d�  #A e�  #A e�  "� d�  "�      B  , , g=  "� g=  #A g�  #A g�  "� g=  "�      B  , , [�  � [�  � \a  � \a  � [�  �      B  , , ^  � ^  � ^�  � ^�  � ^  �      B  , , `S  � `S  � `�  � `�  � `S  �      B  , , b�  � b�  � cK  � cK  � b�  �      B  , , d�  � d�  � e�  � e�  � d�  �      B  , , g=  � g=  � g�  � g�  � g=  �      B  , , i�  � i�  � j5  � j5  � i�  �      B  , , k�  � k�  � l�  � l�  � k�  �      B  , , n'  � n'  � n�  � n�  � n'  �      B  , , pu  � pu  � q  � q  � pu  �      B  , , i�  "� i�  #A j5  #A j5  "� i�  "�      B  , , k�  "� k�  #A l�  #A l�  "� k�  "�      B  , , n'  "� n'  #A n�  #A n�  "� n'  "�      B  , , [�  !C [�  !� \a  !� \a  !C [�  !C      B  , , ^  !C ^  !� ^�  !� ^�  !C ^  !C      B  , , `S  !C `S  !� `�  !� `�  !C `S  !C      B  , , [�  G [�  � \a  � \a  G [�  G      B  , , [�  � [�  I \a  I \a  � [�  �      B  , , ^  � ^  I ^�  I ^�  � ^  �      B  , , `S  � `S  I `�  I `�  � `S  �      B  , , b�  � b�  I cK  I cK  � b�  �      B  , , d�  � d�  I e�  I e�  � d�  �      B  , , g=  � g=  I g�  I g�  � g=  �      B  , , i�  � i�  I j5  I j5  � i�  �      B  , , k�  � k�  I l�  I l�  � k�  �      B  , , n'  � n'  I n�  I n�  � n'  �      B  , , pu  � pu  I q  I q  � pu  �      B  , , ^  G ^  � ^�  � ^�  G ^  G      B  , , `S  G `S  � `�  � `�  G `S  G      B  , , b�  G b�  � cK  � cK  G b�  G      B  , , d�  G d�  � e�  � e�  G d�  G      B  , , g=  G g=  � g�  � g�  G g=  G      B  , , i�  G i�  � j5  � j5  G i�  G      B  , , k�  G k�  � l�  � l�  G k�  G      B  , , n'  G n'  � n�  � n�  G n'  G      B  , , pu  G pu  � q  � q  G pu  G      B  , , b�  !C b�  !� cK  !� cK  !C b�  !C      B  , , d�  !C d�  !� e�  !� e�  !C d�  !C      B  , , [�  � [�   � \a   � \a  � [�  �      B  , , ^  � ^   � ^�   � ^�  � ^  �      B  , , `S  � `S   � `�   � `�  � `S  �      B  , , b�  � b�   � cK   � cK  � b�  �      B  , , d�  � d�   � e�   � e�  � d�  �      B  , , g=  � g=   � g�   � g�  � g=  �      B  , , i�  � i�   � j5   � j5  � i�  �      B  , , [�  � [�  E \a  E \a  � [�  �      B  , , ^  � ^  E ^�  E ^�  � ^  �      B  , , `S  � `S  E `�  E `�  � `S  �      B  , , b�  � b�  E cK  E cK  � b�  �      B  , , d�  � d�  E e�  E e�  � d�  �      B  , , g=  � g=  E g�  E g�  � g=  �      B  , , i�  � i�  E j5  E j5  � i�  �      B  , , k�  � k�  E l�  E l�  � k�  �      B  , , n'  � n'  E n�  E n�  � n'  �      B  , , pu  � pu  E q  E q  � pu  �      B  , , k�  � k�   � l�   � l�  � k�  �      B  , , [�  K [�  � \a  � \a  K [�  K      B  , , ^  K ^  � ^�  � ^�  K ^  K      B  , , `S  K `S  � `�  � `�  K `S  K      B  , , b�  K b�  � cK  � cK  K b�  K      B  , , d�  K d�  � e�  � e�  K d�  K      B  , , g=  K g=  � g�  � g�  K g=  K      B  , , i�  K i�  � j5  � j5  K i�  K      B  , , k�  K k�  � l�  � l�  K k�  K      B  , , n'  K n'  � n�  � n�  K n'  K      B  , , pu  K pu  � q  � q  K pu  K      B  , , n'  � n'   � n�   � n�  � n'  �      B  , , pu  � pu   � q   � q  � pu  �      B  , , g=  !C g=  !� g�  !� g�  !C g=  !C      B  , , i�  !C i�  !� j5  !� j5  !C i�  !C      B  , , k�  !C k�  !� l�  !� l�  !C k�  !C      B  , , n'  !C n'  !� n�  !� n�  !C n'  !C      B  , , pu  !C pu  !� q  !� q  !C pu  !C      B  , , pu  "� pu  #A q  #A q  "� pu  "�      B  , , [�  "� [�  #A \a  #A \a  "� [�  "�      B  , , ^  "� ^  #A ^�  #A ^�  "� ^  "�      B  , , `S  "� `S  #A `�  #A `�  "� `S  "�      B  , , b�  "� b�  #A cK  #A cK  "� b�  "�      B  , , *M  % *M  %� *�  %� *�  % *M  %      B  , , ,�  % ,�  %� -E  %� -E  % ,�  %      B  , , ,�  ') ,�  '� -E  '� -E  ') ,�  ')      B  , , �  % �  %� �  %� �  % �  %      B  , , +  % +  %� �  %� �  % +  %      B  , , y  % y  %� #  %� #  % y  %      B  , , �  % �  %� q  %� q  % �  %      B  , , !  % !  %� !�  %� !�  % !  %      B  , , #c  % #c  %� $  %� $  % #c  %      B  , , %�  % %�  %� &[  %� &[  % %�  %      B  , , '�  % '�  %� (�  %� (�  % '�  %      B  , , -�  *� -�  +� .l  +� .l  *� -�  *�      B  , , -�  ,G -�  ,� .l  ,� .l  ,G -�  ,G      B  , , -�  .� -�  /� .l  /� .l  .� -�  .�      B  , , -�  1� -�  2A .l  2A .l  1� -�  1�      B  , , -�  2� -�  3� .l  3� .l  2� -�  2�      B  , , -�  -� -�  .E .l  .E .l  -� -�  -�      B  , , -�  )� -�  *I .l  *I .l  )� -�  )�      B  , , -�  0C -�  0� .l  0� .l  0C -�  0C      B  , ,   1�   2A �  2A �  1�   1�      B  , , R  1� R  2A �  2A �  1� R  1�      B  , , �  0C �  0� `  0� `  0C �  0C      B  , ,   0C   0� �  0� �  0C   0C      B  , , R  0C R  0� �  0� �  0C R  0C      B  , , �  0C �  0� J  0� J  0C �  0C      B  , , �  -� �  .E `  .E `  -� �  -�      B  , ,   -�   .E �  .E �  -�   -�      B  , , R  -� R  .E �  .E �  -� R  -�      B  , , �  -� �  .E J  .E J  -� �  -�      B  , , �  -� �  .E  �  .E  �  -� �  -�      B  , , "<  -� "<  .E "�  .E "�  -� "<  -�      B  , , �  2� �  3� `  3� `  2� �  2�      B  , , �  ') �  '� �  '� �  ') �  ')      B  , , +  ') +  '� �  '� �  ') +  ')      B  , , y  ') y  '� #  '� #  ') y  ')      B  , , �  ') �  '� q  '� q  ') �  ')      B  , , !  ') !  '� !�  '� !�  ') !  ')      B  , , #c  ') #c  '� $  '� $  ') #c  ')      B  , , %�  ') %�  '� &[  '� &[  ') %�  ')      B  , , '�  ') '�  '� (�  '� (�  ') '�  ')      B  , , *M  ') *M  '� *�  '� *�  ') *M  ')      B  , , +t  ,G +t  ,� ,  ,� ,  ,G +t  ,G      B  , , �  1� �  2A J  2A J  1� �  1�      B  , , �  1� �  2A  �  2A  �  1� �  1�      B  , , "<  1� "<  2A "�  2A "�  1� "<  1�      B  , , )&  1� )&  2A )�  2A )�  1� )&  1�      B  , , +t  1� +t  2A ,  2A ,  1� +t  1�      B  , , "<  ,G "<  ,� "�  ,� "�  ,G "<  ,G      B  , , "<  2� "<  3� "�  3� "�  2� "<  2�      B  , , $�  2� $�  3� %4  3� %4  2� $�  2�      B  , , &�  2� &�  3� '�  3� '�  2� &�  2�      B  , , )&  2� )&  3� )�  3� )�  2� )&  2�      B  , , �  .� �  /� `  /� `  .� �  .�      B  , ,   .�   /� �  /� �  .�   .�      B  , , R  .� R  /� �  /� �  .� R  .�      B  , , �  .� �  /� J  /� J  .� �  .�      B  , , �  .� �  /�  �  /�  �  .� �  .�      B  , , �  *� �  +� `  +� `  *� �  *�      B  , ,   *�   +� �  +� �  *�   *�      B  , , R  *� R  +� �  +� �  *� R  *�      B  , , �  *� �  +� J  +� J  *� �  *�      B  , , �  *� �  +�  �  +�  �  *� �  *�      B  , , "<  *� "<  +� "�  +� "�  *� "<  *�      B  , , $�  *� $�  +� %4  +� %4  *� $�  *�      B  , , &�  *� &�  +� '�  +� '�  *� &�  *�      B  , , )&  *� )&  +� )�  +� )�  *� )&  *�      B  , , +t  *� +t  +� ,  +� ,  *� +t  *�      B  , , +t  2� +t  3� ,  3� ,  2� +t  2�      B  , , "<  .� "<  /� "�  /� "�  .� "<  .�      B  , , �  )� �  *I `  *I `  )� �  )�      B  , ,   )�   *I �  *I �  )�   )�      B  , , $�  -� $�  .E %4  .E %4  -� $�  -�      B  , , &�  -� &�  .E '�  .E '�  -� &�  -�      B  , , )&  -� )&  .E )�  .E )�  -� )&  -�      B  , , +t  -� +t  .E ,  .E ,  -� +t  -�      B  , , $�  .� $�  /� %4  /� %4  .� $�  .�      B  , , R  )� R  *I �  *I �  )� R  )�      B  , , �  )� �  *I J  *I J  )� �  )�      B  , , �  )� �  *I  �  *I  �  )� �  )�      B  , , "<  )� "<  *I "�  *I "�  )� "<  )�      B  , , $�  )� $�  *I %4  *I %4  )� $�  )�      B  , , &�  )� &�  *I '�  *I '�  )� &�  )�      B  , , )&  )� )&  *I )�  *I )�  )� )&  )�      B  , , +t  )� +t  *I ,  *I ,  )� +t  )�      B  , , &�  .� &�  /� '�  /� '�  .� &�  .�      B  , , $�  1� $�  2A %4  2A %4  1� $�  1�      B  , , &�  1� &�  2A '�  2A '�  1� &�  1�      B  , , �  ,G �  ,� `  ,� `  ,G �  ,G      B  , ,   ,G   ,� �  ,� �  ,G   ,G      B  , , R  ,G R  ,� �  ,� �  ,G R  ,G      B  , , �  ,G �  ,� J  ,� J  ,G �  ,G      B  , , �  ,G �  ,�  �  ,�  �  ,G �  ,G      B  , , �  0C �  0�  �  0�  �  0C �  0C      B  , , "<  0C "<  0� "�  0� "�  0C "<  0C      B  , , $�  0C $�  0� %4  0� %4  0C $�  0C      B  , , &�  0C &�  0� '�  0� '�  0C &�  0C      B  , , )&  0C )&  0� )�  0� )�  0C )&  0C      B  , , +t  0C +t  0� ,  0� ,  0C +t  0C      B  , , )&  .� )&  /� )�  /� )�  .� )&  .�      B  , ,   2�   3� �  3� �  2�   2�      B  , , +t  .� +t  /� ,  /� ,  .� +t  .�      B  , , $�  ,G $�  ,� %4  ,� %4  ,G $�  ,G      B  , , &�  ,G &�  ,� '�  ,� '�  ,G &�  ,G      B  , , )&  ,G )&  ,� )�  ,� )�  ,G )&  ,G      B  , , R  2� R  3� �  3� �  2� R  2�      B  , , �  2� �  3� J  3� J  2� �  2�      B  , , �  2� �  3�  �  3�  �  2� �  2�      B  , , �  1� �  2A `  2A `  1� �  1�      B  , , �  "� �  #A  �  #A  �  "� �  "�      B  , , "<  "� "<  #A "�  #A "�  "� "<  "�      B  , , $�  "� $�  #A %4  #A %4  "� $�  "�      B  , , &�  "� &�  #A '�  #A '�  "� &�  "�      B  , , )&  !C )&  !� )�  !� )�  !C )&  !C      B  , ,   !C   !� �  !� �  !C   !C      B  , , +t  !C +t  !� ,  !� ,  !C +t  !C      B  , , R  !C R  !� �  !� �  !C R  !C      B  , , �  � �   � `   � `  � �  �      B  , ,   �    � �   � �  �   �      B  , , �  !C �  !� J  !� J  !C �  !C      B  , , �  !C �  !�  �  !�  �  !C �  !C      B  , , R  � R   � �   � �  � R  �      B  , , �  � �   � J   � J  � �  �      B  , , �  � �   �  �   �  �  � �  �      B  , , "<  � "<   � "�   � "�  � "<  �      B  , , �  � �  � `  � `  � �  �      B  , ,   �   � �  � �  �   �      B  , , R  � R  � �  � �  � R  �      B  , , �  � �  � J  � J  � �  �      B  , , �  � �  �  �  �  �  � �  �      B  , , "<  � "<  � "�  � "�  � "<  �      B  , , $�  � $�  � %4  � %4  � $�  �      B  , , &�  � &�  � '�  � '�  � &�  �      B  , , )&  � )&  � )�  � )�  � )&  �      B  , , +t  � +t  � ,  � ,  � +t  �      B  , , )&  "� )&  #A )�  #A )�  "� )&  "�      B  , , +t  "� +t  #A ,  #A ,  "� +t  "�      B  , , �  K �  � `  � `  K �  K      B  , ,   K   � �  � �  K   K      B  , , R  K R  � �  � �  K R  K      B  , , �  K �  � J  � J  K �  K      B  , , �  K �  �  �  �  �  K �  K      B  , , "<  K "<  � "�  � "�  K "<  K      B  , , $�  K $�  � %4  � %4  K $�  K      B  , , &�  K &�  � '�  � '�  K &�  K      B  , , )&  K )&  � )�  � )�  K )&  K      B  , , +t  K +t  � ,  � ,  K +t  K      B  , , "<  !C "<  !� "�  !� "�  !C "<  !C      B  , , �  � �  I `  I `  � �  �      B  , ,   �   I �  I �  �   �      B  , , R  � R  I �  I �  � R  �      B  , , �  G �  � `  � `  G �  G      B  , ,   G   � �  � �  G   G      B  , , R  G R  � �  � �  G R  G      B  , , �  G �  � J  � J  G �  G      B  , , �  G �  �  �  �  �  G �  G      B  , , "<  G "<  � "�  � "�  G "<  G      B  , , $�  G $�  � %4  � %4  G $�  G      B  , , &�  G &�  � '�  � '�  G &�  G      B  , , )&  G )&  � )�  � )�  G )&  G      B  , , +t  G +t  � ,  � ,  G +t  G      B  , , $�  � $�   � %4   � %4  � $�  �      B  , , &�  � &�   � '�   � '�  � &�  �      B  , , )&  � )&   � )�   � )�  � )&  �      B  , , +t  � +t   � ,   � ,  � +t  �      B  , , �  � �  I J  I J  � �  �      B  , , �  � �  I  �  I  �  � �  �      B  , , "<  � "<  I "�  I "�  � "<  �      B  , , $�  � $�  I %4  I %4  � $�  �      B  , , &�  � &�  I '�  I '�  � &�  �      B  , , )&  � )&  I )�  I )�  � )&  �      B  , , +t  � +t  I ,  I ,  � +t  �      B  , , $�  !C $�  !� %4  !� %4  !C $�  !C      B  , , �  � �  E `  E `  � �  �      B  , ,   �   E �  E �  �   �      B  , , R  � R  E �  E �  � R  �      B  , , �  � �  E J  E J  � �  �      B  , , �  � �  E  �  E  �  � �  �      B  , , "<  � "<  E "�  E "�  � "<  �      B  , , �  !C �  !� `  !� `  !C �  !C      B  , , $�  � $�  E %4  E %4  � $�  �      B  , , &�  � &�  E '�  E '�  � &�  �      B  , , )&  � )&  E )�  E )�  � )&  �      B  , , +t  � +t  E ,  E ,  � +t  �      B  , , &�  !C &�  !� '�  !� '�  !C &�  !C      B  , , �  "� �  #A `  #A `  "� �  "�      B  , ,   "�   #A �  #A �  "�   "�      B  , , R  "� R  #A �  #A �  "� R  "�      B  , , �  "� �  #A J  #A J  "� �  "�      B  , , -�  � -�  I .l  I .l  � -�  �      B  , , -�  "� -�  #A .l  #A .l  "� -�  "�      B  , , -�  G -�  � .l  � .l  G -�  G      B  , , -�  � -�  E .l  E .l  � -�  �      B  , , -�  !C -�  !� .l  !� .l  !C -�  !C      B  , , -�  � -�  � .l  � .l  � -�  �      B  , , -�  K -�  � .l  � .l  K -�  K      B  , , -�  � -�   � .l   � .l  � -�  �      B  , ,  �  �  �  �  ��  �  ��  �  �  �      B  , ,  �G  '.  �G  '�  ��  '�  ��  '.  �G  '.      B  , ,  �  '  �  �  ��  �  ��  '  �  '      B  , ,  [�����  [����G  \b���G  \b����  [�����      B  , ,  �h����  �h���G  ����G  �����  �h����      B  , ,  �����  ����I  �����I  ������  �����      B  , ,  �����  �����  ������  ������  �����      B  , ,  ����/  �����  ������  �����/  ����/      B  , ,  ����  �����  ������  �����  ����      B  , ,  ���ϕ  ����?  �����?  ����ϕ  ���ϕ      B  , ,  �����  ���·  ����·  ������  �����      B  , ,  ����%  �����  ������  �����%  ����%      B  , ,  ����  ���ʽ  ����ʽ  �����  ����      B  , ,  ��  %  ��  %�  �C  %�  �C  %  ��  %      B  , ,  ��  %  ��  %�  ��  %�  ��  %  ��  %      B  , ,  �5  %  �5  %�  ��  %�  ��  %  �5  %      B  , ,  ��  %  ��  %�  �-  %�  �-  %  ��  %      B  , ,  �  %  �  %� {  %� {  %  �  %      B  , ,   %   %� �  %� �  %   %      B  , , m  % m  %�   %�   % m  %      B  , , �  % �  %� e  %� e  % �  %      B  , , 
	  % 
	  %� 
�  %� 
�  % 
	  %      B  , , W  % W  %�   %�   % W  %      B  , , �  % �  %� O  %� O  % �  %      B  , , �  % �  %� �  %� �  % �  %      B  , , A  % A  %� �  %� �  % A  %      B  , , A  ') A  '� �  '� �  ') A  ')      B  , ,  ��  .�  ��  /�  T  /�  T  .�  ��  .�      B  , , �  .� �  /� �  /� �  .� �  .�      B  , , F  .� F  /� �  /� �  .� F  .�      B  , , �  .� �  /� >  /� >  .� �  .�      B  , , �  .� �  /� 	�  /� 	�  .� �  .�      B  , , 0  .� 0  /� �  /� �  .� 0  .�      B  , , ~  .� ~  /� (  /� (  .� ~  .�      B  , , �  .� �  /� v  /� v  .� �  .�      B  , ,   1�   2A �  2A �  1�   1�      B  , ,   .�   /� �  /� �  .�   .�      B  , , h  .� h  /�   /�   .� h  .�      B  , ,  ��  0C  ��  0�  T  0�  T  0C  ��  0C      B  , , �  0C �  0� �  0� �  0C �  0C      B  , , F  0C F  0� �  0� �  0C F  0C      B  , , �  0C �  0� >  0� >  0C �  0C      B  , , �  0C �  0� 	�  0� 	�  0C �  0C      B  , , 0  0C 0  0� �  0� �  0C 0  0C      B  , , ~  0C ~  0� (  0� (  0C ~  0C      B  , , �  0C �  0� v  0� v  0C �  0C      B  , ,   0C   0� �  0� �  0C   0C      B  , , h  0C h  0�   0�   0C h  0C      B  , ,  ��  )�  ��  *I  T  *I  T  )�  ��  )�      B  , , �  )� �  *I �  *I �  )� �  )�      B  , , F  )� F  *I �  *I �  )� F  )�      B  , , �  )� �  *I >  *I >  )� �  )�      B  , , �  )� �  *I 	�  *I 	�  )� �  )�      B  , , 0  )� 0  *I �  *I �  )� 0  )�      B  , , ~  )� ~  *I (  *I (  )� ~  )�      B  , , �  )� �  *I v  *I v  )� �  )�      B  , ,   )�   *I �  *I �  )�   )�      B  , , h  )� h  *I   *I   )� h  )�      B  , ,  ��  -�  ��  .E  T  .E  T  -�  ��  -�      B  , , �  -� �  .E �  .E �  -� �  -�      B  , , F  -� F  .E �  .E �  -� F  -�      B  , , �  -� �  .E >  .E >  -� �  -�      B  , , �  -� �  .E 	�  .E 	�  -� �  -�      B  , , 0  -� 0  .E �  .E �  -� 0  -�      B  , , ~  -� ~  .E (  .E (  -� ~  -�      B  , , �  -� �  .E v  .E v  -� �  -�      B  , ,   -�   .E �  .E �  -�   -�      B  , , h  -� h  .E   .E   -� h  -�      B  , ,  ��  *�  ��  +�  T  +�  T  *�  ��  *�      B  , , �  *� �  +� �  +� �  *� �  *�      B  , , F  *� F  +� �  +� �  *� F  *�      B  , , �  *� �  +� >  +� >  *� �  *�      B  , , �  *� �  +� 	�  +� 	�  *� �  *�      B  , , 0  *� 0  +� �  +� �  *� 0  *�      B  , , ~  *� ~  +� (  +� (  *� ~  *�      B  , , �  *� �  +� v  +� v  *� �  *�      B  , ,   *�   +� �  +� �  *�   *�      B  , , h  *� h  +�   +�   *� h  *�      B  , ,  ��  ,G  ��  ,�  T  ,�  T  ,G  ��  ,G      B  , , �  ,G �  ,� �  ,� �  ,G �  ,G      B  , , F  ,G F  ,� �  ,� �  ,G F  ,G      B  , ,   2�   3� �  3� �  2�   2�      B  , , h  2� h  3�   3�   2� h  2�      B  , , ~  1� ~  2A (  2A (  1� ~  1�      B  , , �  1� �  2A v  2A v  1� �  1�      B  , ,  ��  ')  ��  '�  �-  '�  �-  ')  ��  ')      B  , ,  �  ')  �  '� {  '� {  ')  �  ')      B  , ,   ')   '� �  '� �  ')   ')      B  , , m  ') m  '�   '�   ') m  ')      B  , , �  ') �  '� e  '� e  ') �  ')      B  , , 
	  ') 
	  '� 
�  '� 
�  ') 
	  ')      B  , , W  ') W  '�   '�   ') W  ')      B  , , �  ') �  '� O  '� O  ') �  ')      B  , , �  ') �  '� �  '� �  ') �  ')      B  , , �  ,G �  ,� >  ,� >  ,G �  ,G      B  , , �  ,G �  ,� 	�  ,� 	�  ,G �  ,G      B  , , 0  ,G 0  ,� �  ,� �  ,G 0  ,G      B  , , ~  ,G ~  ,� (  ,� (  ,G ~  ,G      B  , , �  ,G �  ,� v  ,� v  ,G �  ,G      B  , ,   ,G   ,� �  ,� �  ,G   ,G      B  , , h  ,G h  ,�   ,�   ,G h  ,G      B  , ,  ��  1�  ��  2A  T  2A  T  1�  ��  1�      B  , , �  1� �  2A �  2A �  1� �  1�      B  , , F  1� F  2A �  2A �  1� F  1�      B  , , �  1� �  2A >  2A >  1� �  1�      B  , , �  1� �  2A 	�  2A 	�  1� �  1�      B  , , 0  1� 0  2A �  2A �  1� 0  1�      B  , , h  1� h  2A   2A   1� h  1�      B  , ,  ��  2�  ��  3�  T  3�  T  2�  ��  2�      B  , , �  2� �  3� �  3� �  2� �  2�      B  , , F  2� F  3� �  3� �  2� F  2�      B  , , �  2� �  3� >  3� >  2� �  2�      B  , , �  2� �  3� 	�  3� 	�  2� �  2�      B  , , 0  2� 0  3� �  3� �  2� 0  2�      B  , , ~  2� ~  3� (  3� (  2� ~  2�      B  , , �  2� �  3� v  3� v  2� �  2�      B  , ,  �\  -�  �\  .E  �  .E  �  -�  �\  -�      B  , ,  �\  0C  �\  0�  �  0�  �  0C  �\  0C      B  , ,  �\  2�  �\  3�  �  3�  �  2�  �\  2�      B  , ,  �\  )�  �\  *I  �  *I  �  )�  �\  )�      B  , ,  �\  .�  �\  /�  �  /�  �  .�  �\  .�      B  , ,  �\  1�  �\  2A  �  2A  �  1�  �\  1�      B  , ,  �\  *�  �\  +�  �  +�  �  *�  �\  *�      B  , ,  ��  ')  ��  '�  ��  '�  ��  ')  ��  ')      B  , ,  �5  ')  �5  '�  ��  '�  ��  ')  �5  ')      B  , ,  �\  ,G  �\  ,�  �  ,�  �  ,G  �\  ,G      B  , ,  ��  ')  ��  '�  �C  '�  �C  ')  ��  ')      B  , ,  �\  G  �\  �  �  �  �  G  �\  G      B  , ,  �\  "�  �\  #A  �  #A  �  "�  �\  "�      B  , ,  �\  �  �\  I  �  I  �  �  �\  �      B  , ,  �\  �  �\  E  �  E  �  �  �\  �      B  , ,  �\  �  �\  �  �  �  �  �  �\  �      B  , ,  �\  �  �\   �  �   �  �  �  �\  �      B  , ,  �\  !C  �\  !�  �  !�  �  !C  �\  !C      B  , ,  �\  K  �\  �  �  �  �  K  �\  K      B  , , �  � �  � �  � �  � �  �      B  , , F  � F  � �  � �  � F  �      B  , ,  ��  !C  ��  !�  T  !�  T  !C  ��  !C      B  , , �  !C �  !� �  !� �  !C �  !C      B  , , �  � �  � >  � >  � �  �      B  , ,  ��  K  ��  �  T  �  T  K  ��  K      B  , , �  K �  � �  � �  K �  K      B  , , F  K F  � �  � �  K F  K      B  , , �  K �  � >  � >  K �  K      B  , , �  K �  � 	�  � 	�  K �  K      B  , , 0  K 0  � �  � �  K 0  K      B  , , ~  K ~  � (  � (  K ~  K      B  , , �  K �  � v  � v  K �  K      B  , ,   K   � �  � �  K   K      B  , , h  K h  �   �   K h  K      B  , , F  !C F  !� �  !� �  !C F  !C      B  , , �  !C �  !� >  !� >  !C �  !C      B  , , �  !C �  !� 	�  !� 	�  !C �  !C      B  , , 0  !C 0  !� �  !� �  !C 0  !C      B  , , ~  !C ~  !� (  !� (  !C ~  !C      B  , , �  !C �  !� v  !� v  !C �  !C      B  , ,   !C   !� �  !� �  !C   !C      B  , , h  !C h  !�   !�   !C h  !C      B  , ,  ��  "�  ��  #A  T  #A  T  "�  ��  "�      B  , ,  ��  �  ��  E  T  E  T  �  ��  �      B  , , �  � �  E �  E �  � �  �      B  , , F  � F  E �  E �  � F  �      B  , , �  � �  E >  E >  � �  �      B  , , �  � �  E 	�  E 	�  � �  �      B  , , 0  � 0  E �  E �  � 0  �      B  , , ~  � ~  E (  E (  � ~  �      B  , ,  ��  G  ��  �  T  �  T  G  ��  G      B  , , �  G �  � �  � �  G �  G      B  , , F  G F  � �  � �  G F  G      B  , , �  G �  � >  � >  G �  G      B  , , �  G �  � 	�  � 	�  G �  G      B  , , 0  G 0  � �  � �  G 0  G      B  , , ~  G ~  � (  � (  G ~  G      B  , , �  G �  � v  � v  G �  G      B  , ,   G   � �  � �  G   G      B  , , h  G h  �   �   G h  G      B  , , �  � �  E v  E v  � �  �      B  , ,   �   E �  E �  �   �      B  , , h  � h  E   E   � h  �      B  , , �  "� �  #A �  #A �  "� �  "�      B  , , F  "� F  #A �  #A �  "� F  "�      B  , , �  "� �  #A >  #A >  "� �  "�      B  , , �  "� �  #A 	�  #A 	�  "� �  "�      B  , , 0  "� 0  #A �  #A �  "� 0  "�      B  , , ~  "� ~  #A (  #A (  "� ~  "�      B  , , �  "� �  #A v  #A v  "� �  "�      B  , ,   "�   #A �  #A �  "�   "�      B  , , h  "� h  #A   #A   "� h  "�      B  , , �  � �  � 	�  � 	�  � �  �      B  , , 0  � 0  � �  � �  � 0  �      B  , , ~  � ~  � (  � (  � ~  �      B  , , �  � �  � v  � v  � �  �      B  , ,   �   � �  � �  �   �      B  , , h  � h  �   �   � h  �      B  , , ~  � ~   � (   � (  � ~  �      B  , , �  � �   � v   � v  � �  �      B  , ,   �    � �   � �  �   �      B  , , h  � h   �    �   � h  �      B  , , F  � F   � �   � �  � F  �      B  , , �  � �   � >   � >  � �  �      B  , , �  � �   � 	�   � 	�  � �  �      B  , , 0  � 0   � �   � �  � 0  �      B  , ,  ��  �  ��   �  T   �  T  �  ��  �      B  , , �  � �   � �   � �  � �  �      B  , ,  ��  �  ��  I  T  I  T  �  ��  �      B  , , �  � �  I �  I �  � �  �      B  , , F  � F  I �  I �  � F  �      B  , , �  � �  I >  I >  � �  �      B  , , �  � �  I 	�  I 	�  � �  �      B  , , 0  � 0  I �  I �  � 0  �      B  , , ~  � ~  I (  I (  � ~  �      B  , , �  � �  I v  I v  � �  �      B  , ,   �   I �  I �  �   �      B  , , h  � h  I   I   � h  �      B  , ,  ��  �  ��  �  T  �  T  �  ��  �      B  , ,  �^  �  �^  �  �  �  �  �  �^  �      B  , ,  ʲ  �  ʲ  �  �\  �  �\  �  ʲ  �      B  , ,  �  �  �  �  ̰  �  ̰  �  �  �      B  , ,  �Z  �  �Z  �  �  �  �  �  �Z  �      B  , ,  ��  '.  ��  '�  �?  '�  �?  '.  ��  '.      B  , ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      B  , ,  �1  '.  �1  '�  ��  '�  ��  '.  �1  '.      B  , ,  �  '.  �  '�  �)  '�  �)  '.  �  '.      B  , ,  ��  '.  ��  '�  �w  '�  �w  '.  ��  '.      B  , ,  �  '.  �  '�  ��  '�  ��  '.  �  '.      B  , ,  �i  '.  �i  '�  �  '�  �  '.  �i  '.      B  , ,  ή  �  ή  �  �X  �  �X  �  ή  �      B  , ,  �  �  �  �  Ь  �  Ь  �  �  �      B  , ,  �V  �  �V  �  �   �  �   �  �V  �      B  , ,  �n  �  �n  �  �  �  �  �  �n  �      B  , ,  ��  �  ��  �  �l  �  �l  �  ��  �      B  , ,  �  �  �  �  ��  �  ��  �  �  �      B  , ,  �j  �  �j  �  �  �  �  �  �j  �      B  , ,  ��  �  ��  �  �h  �  �h  �  ��  �      B  , ,  �n  '  �n  �  �  �  �  '  �n  '      B  , ,  ��  '  ��  �  �l  �  �l  '  ��  '      B  , ,  �  '  �  �  ��  �  ��  '  �  '      B  , ,  �j  '  �j  �  �  �  �  '  �j  '      B  , ,  ��  '  ��  �  �h  �  �h  '  ��  '      B  , ,  �  '  �  �  ��  �  ��  '  �  '      B  , ,  �f  '  �f  �  �  �  �  '  �f  '      B  , ,  º  '  º  �  �d  �  �d  '  º  '      B  , ,  �  '  �  �  ĸ  �  ĸ  '  �  '      B  , ,  �b  '  �b  �  �  �  �  '  �b  '      B  , ,  ƶ  '  ƶ  �  �`  �  �`  '  ƶ  '      B  , ,  �
  '  �
  �  ȴ  �  ȴ  '  �
  '      B  , ,  �^  '  �^  �  �  �  �  '  �^  '      B  , ,  ʲ  '  ʲ  �  �\  �  �\  '  ʲ  '      B  , ,  �  '  �  �  ̰  �  ̰  '  �  '      B  , ,  �Z  '  �Z  �  �  �  �  '  �Z  '      B  , ,  �h  )  �h  �  �  �  �  )  �h  )      B  , ,  �h  �  �h    �    �  �  �h  �      B  , ,  ή  '  ή  �  �X  �  �X  '  ή  '      B  , ,  �  '  �  �  Ь  �  Ь  '  �  '      B  , ,  �V  '  �V  �  �   �  �   '  �V  '      B  , ,  �  �  �  �  ��  �  ��  �  �  �      B  , ,  �f  �  �f  �  �  �  �  �  �f  �      B  , ,  º  �  º  �  �d  �  �d  �  º  �      B  , ,  �  �  �  �  ĸ  �  ĸ  �  �  �      B  , ,  �b  �  �b  �  �  �  �  �  �b  �      B  , ,  ƶ  �  ƶ  �  �`  �  �`  �  ƶ  �      B  , ,  �
  �  �
  �  ȴ  �  ȴ  �  �
  �      B  , ,  ��  �  ��    ��    ��  �  ��  �      B  , ,  �I  �  �I    ��    ��  �  �I  �      B  , ,  ��  �  ��    �A    �A  �  ��  �      B  , ,  ��  �  ��    ��    ��  �  ��  �      B  , ,  �3  �  �3    ��    ��  �  �3  �      B  , ,  ā  �  ā    �+    �+  �  ā  �      B  , ,  ��  �  ��    �y    �y  �  ��  �      B  , ,  �  �  �    ��    ��  �  �  �      B  , ,  �k  �  �k    �    �  �  �k  �      B  , ,  ͹  �  ͹    �c    �c  �  ͹  �      B  , ,  �  �  �    б    б  �  �  �      B  , ,  �h  9  �h  �  �  �  �  9  �h  9      B  , ,  �.  �  �.  e  ��  e  ��  �  �.  �      B  , ,  �h  �  �h  3  �  3  �  �  �h  �      B  , ,  �.  g  �.    ��    ��  g  �.  g      B  , ,  �h  5  �h  �  �  �  �  5  �h  5      B  , ,  �h  
�  �h  �  �  �  �  
�  �h  
�      B  , ,  �  	�  �  
�  б  
�  б  	�  �  	�      B  , ,  �h  	�  �h  
7  �  
7  �  	�  �h  	�      B  , ,  �.  �  �.  ]  ��  ]  ��  �  �.  �      B  , ,  �h  �  �h  +  �  +  �  �  �h  �      B  , ,  �.  _  �.  	  ��  	  ��  _  �.  _      B  , ,  �h  -  �h  �  �  �  �  -  �h  -      B  , ,  �.    �.  �  ��  �  ��    �.        B  , ,  �h  �  �h  �  �  �  �  �  �h  �      B  , ,  �.  �  �.  a  ��  a  ��  �  �.  �      B  , ,  �h  �  �h  /  �  /  �  �  �h  �      B  , ,  �.  c  �.    ��    ��  c  �.  c      B  , ,  �h  1  �h  �  �  �  �  1  �h  1      B  , ,  �.    �.  �  ��  �  ��    �.        B  , ,  �h  �  �h  �  �  �  �  �  �h  �      B  , ,  Ũ  �  Ũ  a  �R  a  �R  �  Ũ  �      B  , ,  ��  �  ��  a  Ƞ  a  Ƞ  �  ��  �      B  , ,  �D  �  �D  a  ��  a  ��  �  �D  �      B  , ,  ̒  �  ̒  a  �<  a  �<  �  ̒  �      B  , ,  ��  �  ��  a  ϊ  a  ϊ  �  ��  �      B  , ,  �Z  _  �Z  	  �  	  �  _  �Z  _      B  , ,  Ũ  _  Ũ  	  �R  	  �R  _  Ũ  _      B  , ,  �"  c  �"    ��    ��  c  �"  c      B  , ,  �p  c  �p    �    �  c  �p  c      B  , ,  ��  c  ��    �h    �h  c  ��  c      B  , ,  �  c  �    ��    ��  c  �  c      B  , ,  �Z  c  �Z    �    �  c  �Z  c      B  , ,  Ũ  c  Ũ    �R    �R  c  Ũ  c      B  , ,  ��  c  ��    Ƞ    Ƞ  c  ��  c      B  , ,  �D  c  �D    ��    ��  c  �D  c      B  , ,  ̒  c  ̒    �<    �<  c  ̒  c      B  , ,  ��  c  ��    ϊ    ϊ  c  ��  c      B  , ,  ��  _  ��  	  Ƞ  	  Ƞ  _  ��  _      B  , ,  �D  _  �D  	  ��  	  ��  _  �D  _      B  , ,  �"    �"  �  ��  �  ��    �"        B  , ,  �p    �p  �  �  �  �    �p        B  , ,  ��    ��  �  �h  �  �h    ��        B  , ,  �    �  �  ��  �  ��    �        B  , ,  �Z    �Z  �  �  �  �    �Z        B  , ,  Ũ    Ũ  �  �R  �  �R    Ũ        B  , ,  ��    ��  �  Ƞ  �  Ƞ    ��        B  , ,  �D    �D  �  ��  �  ��    �D        B  , ,  ̒    ̒  �  �<  �  �<    ̒        B  , ,  ��    ��  �  ϊ  �  ϊ    ��        B  , ,  ̒  _  ̒  	  �<  	  �<  _  ̒  _      B  , ,  ��  _  ��  	  ϊ  	  ϊ  _  ��  _      B  , ,  �"  �  �"  e  ��  e  ��  �  �"  �      B  , ,  �p  �  �p  e  �  e  �  �  �p  �      B  , ,  ��  �  ��  e  �h  e  �h  �  ��  �      B  , ,  �  �  �  e  ��  e  ��  �  �  �      B  , ,  �Z  �  �Z  e  �  e  �  �  �Z  �      B  , ,  Ũ  �  Ũ  e  �R  e  �R  �  Ũ  �      B  , ,  ��  �  ��  e  Ƞ  e  Ƞ  �  ��  �      B  , ,  �D  �  �D  e  ��  e  ��  �  �D  �      B  , ,  ̒  �  ̒  e  �<  e  �<  �  ̒  �      B  , ,  ��  �  ��  e  ϊ  e  ϊ  �  ��  �      B  , ,  �"  _  �"  	  ��  	  ��  _  �"  _      B  , ,  �p  _  �p  	  �  	  �  _  �p  _      B  , ,  �"  g  �"    ��    ��  g  �"  g      B  , ,  �p  g  �p    �    �  g  �p  g      B  , ,  ��  g  ��    �h    �h  g  ��  g      B  , ,  �  g  �    ��    ��  g  �  g      B  , ,  �Z  g  �Z    �    �  g  �Z  g      B  , ,  Ũ  g  Ũ    �R    �R  g  Ũ  g      B  , ,  ��  g  ��    Ƞ    Ƞ  g  ��  g      B  , ,  �D  g  �D    ��    ��  g  �D  g      B  , ,  ̒  g  ̒    �<    �<  g  ̒  g      B  , ,  ��  g  ��    ϊ    ϊ  g  ��  g      B  , ,  �"    �"  �  ��  �  ��    �"        B  , ,  �p    �p  �  �  �  �    �p        B  , ,  ��    ��  �  �h  �  �h    ��        B  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      B  , ,  �I  	�  �I  
�  ��  
�  ��  	�  �I  	�      B  , ,  ��  	�  ��  
�  �A  
�  �A  	�  ��  	�      B  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      B  , ,  �3  	�  �3  
�  ��  
�  ��  	�  �3  	�      B  , ,  ā  	�  ā  
�  �+  
�  �+  	�  ā  	�      B  , ,  ��  	�  ��  
�  �y  
�  �y  	�  ��  	�      B  , ,  �  	�  �  
�  ��  
�  ��  	�  �  	�      B  , ,  �k  	�  �k  
�  �  
�  �  	�  �k  	�      B  , ,  ͹  	�  ͹  
�  �c  
�  �c  	�  ͹  	�      B  , ,  �    �  �  ��  �  ��    �        B  , ,  �Z    �Z  �  �  �  �    �Z        B  , ,  Ũ    Ũ  �  �R  �  �R    Ũ        B  , ,  ��    ��  �  Ƞ  �  Ƞ    ��        B  , ,  �D    �D  �  ��  �  ��    �D        B  , ,  ̒    ̒  �  �<  �  �<    ̒        B  , ,  ��    ��  �  ϊ  �  ϊ    ��        B  , ,  ��  _  ��  	  �h  	  �h  _  ��  _      B  , ,  �  _  �  	  ��  	  ��  _  �  _      B  , ,  �"  �  �"  a  ��  a  ��  �  �"  �      B  , ,  �p  �  �p  a  �  a  �  �  �p  �      B  , ,  ��  �  ��  a  �h  a  �h  �  ��  �      B  , ,  �  �  �  a  ��  a  ��  �  �  �      B  , ,  �Z  �  �Z  a  �  a  �  �  �Z  �      B  , ,  �"  �  �"  ]  ��  ]  ��  �  �"  �      B  , ,  �p  �  �p  ]  �  ]  �  �  �p  �      B  , ,  ��  �  ��  ]  �h  ]  �h  �  ��  �      B  , ,  �  �  �  ]  ��  ]  ��  �  �  �      B  , ,  �Z  �  �Z  ]  �  ]  �  �  �Z  �      B  , ,  Ũ  �  Ũ  ]  �R  ]  �R  �  Ũ  �      B  , ,  ��  �  ��  ]  Ƞ  ]  Ƞ  �  ��  �      B  , ,  �D  �  �D  ]  ��  ]  ��  �  �D  �      B  , ,  ̒  �  ̒  ]  �<  ]  �<  �  ̒  �      B  , ,  ��  �  ��  ]  ϊ  ]  ϊ  �  ��  �      B  , ,  �"    �"  �  ��  �  ��    �"        B  , ,  �p    �p  �  �  �  �    �p        B  , ,  ��    ��  �  �h  �  �h    ��        B  , ,  �    �  �  ��  �  ��    �        B  , ,  �Z    �Z  �  �  �  �    �Z        B  , ,  Ũ    Ũ  �  �R  �  �R    Ũ        B  , ,  ��    ��  �  Ƞ  �  Ƞ    ��        B  , ,  �D    �D  �  ��  �  ��    �D        B  , ,  ̒    ̒  �  �<  �  �<    ̒        B  , ,  ��    ��  �  ϊ  �  ϊ    ��        B  , ,  �"  �  �"  a  ��  a  ��  �  �"  �      B  , ,  �p  �  �p  a  �  a  �  �  �p  �      B  , ,  ��  �  ��  a  �h  a  �h  �  ��  �      B  , ,  �  �  �  a  ��  a  ��  �  �  �      B  , ,  �Z  �  �Z  a  �  a  �  �  �Z  �      B  , ,  Ũ  �  Ũ  a  �R  a  �R  �  Ũ  �      B  , ,  ��  �  ��  a  Ƞ  a  Ƞ  �  ��  �      B  , ,  �D  �  �D  a  ��  a  ��  �  �D  �      B  , ,  ̒  �  ̒  a  �<  a  �<  �  ̒  �      B  , ,  ��  �  ��  a  ϊ  a  ϊ  �  ��  �      B  , ,  �"  c  �"    ��    ��  c  �"  c      B  , ,  �p  c  �p    �    �  c  �p  c      B  , ,  ��  c  ��    �h    �h  c  ��  c      B  , ,  �  c  �    ��    ��  c  �  c      B  , ,  �Z  c  �Z    �    �  c  �Z  c      B  , ,  Ũ  c  Ũ    �R    �R  c  Ũ  c      B  , ,  ��  c  ��    Ƞ    Ƞ  c  ��  c      B  , ,  �D  c  �D    ��    ��  c  �D  c      B  , ,  ̒  c  ̒    �<    �<  c  ̒  c      B  , ,  ��  c  ��    ϊ    ϊ  c  ��  c      B  , ,  �"     �"   �  ��   �  ��     �"         B  , ,  �p     �p   �  �   �  �     �p         B  , ,  ��     ��   �  �h   �  �h     ��         B  , ,  �     �   �  ��   �  ��     �         B  , ,  �Z     �Z   �  �   �  �     �Z         B  , ,  Ũ     Ũ   �  �R   �  �R     Ũ         B  , ,  ��     ��   �  Ƞ   �  Ƞ     ��         B  , ,  �D     �D   �  ��   �  ��     �D         B  , ,  ̒     ̒   �  �<   �  �<     ̒         B  , ,  ��     ��   �  ϊ   �  ϊ     ��         B  , ,  �"����  �"���e  �����e  ������  �"����      B  , ,  �p����  �p���e  ����e  �����  �p����      B  , ,  ������  �����e  �h���e  �h����  ������      B  , ,  �����  ����e  �����e  ������  �����      B  , ,  �Z����  �Z���e  ����e  �����  �Z����      B  , ,  Ũ����  Ũ���e  �R���e  �R����  Ũ����      B  , ,  ������  �����e  Ƞ���e  Ƞ����  ������      B  , ,  �D����  �D���e  �����e  ������  �D����      B  , ,  ̒����  ̒���e  �<���e  �<����  ̒����      B  , ,  ������  �����e  ϊ���e  ϊ����  ������      B  , ,  �"���g  �"���  �����  �����g  �"���g      B  , ,  �p���g  �p���  ����  ����g  �p���g      B  , ,  �����g  �����  �h���  �h���g  �����g      B  , ,  ����g  ����  �����  �����g  ����g      B  , ,  �Z���g  �Z���  ����  ����g  �Z���g      B  , ,  Ũ���g  Ũ���  �R���  �R���g  Ũ���g      B  , ,  �����g  �����  Ƞ���  Ƞ���g  �����g      B  , ,  �D���g  �D���  �����  �����g  �D���g      B  , ,  ̒���g  ̒���  �<���  �<���g  ̒���g      B  , ,  �����g  �����  ϊ���  ϊ���g  �����g      B  , ,  �"���  �"����  ������  �����  �"���      B  , ,  �p���  �p����  �����  ����  �p���      B  , ,  �����  ������  �h����  �h���  �����      B  , ,  ����  �����  ������  �����  ����      B  , ,  �Z���  �Z����  �����  ����  �Z���      B  , ,  Ũ���  Ũ����  �R����  �R���  Ũ���      B  , ,  �����  ������  Ƞ����  Ƞ���  �����      B  , ,  �D���  �D����  ������  �����  �D���      B  , ,  ̒���  ̒����  �<����  �<���  ̒���      B  , ,  �����  ������  ϊ����  ϊ���  �����      B  , ,  �"  _  �"  	  ��  	  ��  _  �"  _      B  , ,  �p  _  �p  	  �  	  �  _  �p  _      B  , ,  ��  _  ��  	  �h  	  �h  _  ��  _      B  , ,  �  _  �  	  ��  	  ��  _  �  _      B  , ,  �Z  _  �Z  	  �  	  �  _  �Z  _      B  , ,  Ũ  _  Ũ  	  �R  	  �R  _  Ũ  _      B  , ,  ��  _  ��  	  Ƞ  	  Ƞ  _  ��  _      B  , ,  �D  _  �D  	  ��  	  ��  _  �D  _      B  , ,  ̒  _  ̒  	  �<  	  �<  _  ̒  _      B  , ,  ��  _  ��  	  ϊ  	  ϊ  _  ��  _      B  , ,  �.  �  �.  a  ��  a  ��  �  �.  �      B  , ,  �h  �  �h  �  �  �  �  �  �h  �      B  , ,  �.  _  �.  	  ��  	  ��  _  �.  _      B  , ,  �h  �  �h  ;  �  ;  �  �  �h  �      B  , ,  �h  �  �h  �  �  �  �  �  �h  �      B  , ,  �.���  �.����  ������  �����  �.���      B  , ,  �h���E  �h����  �����  ����E  �h���E      B  , ,  �h����  �h����  �����  �����  �h����      B  , ,  �.  c  �.    ��    ��  c  �.  c      B  , ,  �h  �  �h  ?  �  ?  �  �  �h  �      B  , ,  �.    �.  �  ��  �  ��    �.        B  , ,  �.���g  �.���  �����  �����g  �.���g      B  , ,  �h����  �h���C  ����C  �����  �h����      B  , ,  �.     �.   �  ��   �  ��     �.         B  , ,  �.����  �.���e  �����e  ������  �.����      B  , ,  �h����  �h����  �����  �����  �h����      B  , ,  �h   A  �h   �  �   �  �   A  �h   A      B  , ,  �h  =  �h  �  �  �  �  =  �h  =      B  , ,  ��    ��  �  �f  �  �f    ��        B  , ,  ��  �  ��  a  �f  a  �f  �  ��  �      B  , ,  ��  �  ��  �  �H  �  �H  �  ��  �      B  , ,  ��  c  ��    �f    �f  c  ��  c      B  , ,  ��    ��  �  �f  �  �f    ��        B  , ,  ��  �  ��  e  �f  e  �f  �  ��  �      B  , ,  ��  g  ��    �f    �f  g  ��  g      B  , ,  ��  '  ��  �  �H  �  �H  '  ��  '      B  , ,  ��  _  ��  	  �f  	  �f  _  ��  _      B  , ,  ��    ��  �  �f  �  �f    ��        B  , ,  ��  �  ��  a  �f  a  �f  �  ��  �      B  , ,  ��  c  ��    �f    �f  c  ��  c      B  , ,  ��     ��   �  �f   �  �f     ��         B  , ,  ��  �  ��  ]  �f  ]  �f  �  ��  �      B  , ,  ������  �����e  �f���e  �f����  ������      B  , ,  �����g  �����  �f���  �f���g  �����g      B  , ,  �����  ������  �f����  �f���  �����      B  , ,  ��  _  ��  	  �f  	  �f  _  ��  _      B  , ,  ��  �  ��  �  �@  �  �@  �  ��  �      B  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      B  , ,  �>  �  �>  �  ��  �  ��  �  �>  �      B  , ,  �c  '.  �c  '�  �  '�  �  '.  �c  '.      B  , ,  ��  �  ��  �  �<  �  �<  �  ��  �      B  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      B  , ,  �:  �  �:  �  ��  �  ��  �  �:  �      B  , ,  ��  �  ��  �  �8  �  �8  �  ��  �      B  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      B  , ,  �6  �  �6  �  ��  �  ��  �  �6  �      B  , ,  ��  �  ��  �  �4  �  �4  �  ��  �      B  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      B  , ,  �2  �  �2  �  ��  �  ��  �  �2  �      B  , ,  ��  �  ��  �  �0  �  �0  �  ��  �      B  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      B  , ,  �.  �  �.  �  ��  �  ��  �  �.  �      B  , ,  �%  '.  �%  '�  ��  '�  ��  '.  �%  '.      B  , ,  ��  �  ��  �  �,  �  �,  �  ��  �      B  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      B  , ,  �*  �  �*  �  ��  �  ��  �  �*  �      B  , ,  �~  �  �~  �  �(  �  �(  �  �~  �      B  , ,  ��  �  ��  �  �|  �  �|  �  ��  �      B  , ,  �&  �  �&  �  ��  �  ��  �  �&  �      B  , ,  �z  �  �z  �  �$  �  �$  �  �z  �      B  , ,  ��  �  ��  �  �x  �  �x  �  ��  �      B  , ,  �"  �  �"  �  ��  �  ��  �  �"  �      B  , ,  �v  �  �v  �  �   �  �   �  �v  �      B  , ,  ��  �  ��  �  �t  �  �t  �  ��  �      B  , ,  �  �  �  �  ��  �  ��  �  �  �      B  , ,  �s  '.  �s  '�  �  '�  �  '.  �s  '.      B  , ,  �r  �  �r  �  �  �  �  �  �r  �      B  , ,  ��  �  ��  �  �p  �  �p  �  ��  �      B  , ,  �y  '.  �y  '�  �#  '�  �#  '.  �y  '.      B  , ,  ��  '.  ��  '�  �9  '�  �9  '.  ��  '.      B  , ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      B  , ,  �+  '.  �+  '�  ��  '�  ��  '.  �+  '.      B  , ,  ��  '.  ��  '�  �k  '�  �k  '.  ��  '.      B  , ,  �  '.  �  '�  ��  '�  ��  '.  �  '.      B  , ,  ��  '  ��  �  ��  �  ��  '  ��  '      B  , ,  �F  '  �F  �  ��  �  ��  '  �F  '      B  , ,  ��  '  ��  �  �D  �  �D  '  ��  '      B  , ,  ��  '  ��  �  ��  �  ��  '  ��  '      B  , ,  �B  '  �B  �  ��  �  ��  '  �B  '      B  , ,  ��  '  ��  �  �@  �  �@  '  ��  '      B  , ,  ��  '  ��  �  ��  �  ��  '  ��  '      B  , ,  �>  '  �>  �  ��  �  ��  '  �>  '      B  , ,  ��  '  ��  �  �<  �  �<  '  ��  '      B  , ,  ��  '  ��  �  ��  �  ��  '  ��  '      B  , ,  �]  '.  �]  '�  �  '�  �  '.  �]  '.      B  , ,  �:  '  �:  �  ��  �  ��  '  �:  '      B  , ,  ��  '  ��  �  �8  �  �8  '  ��  '      B  , ,  ��  '  ��  �  ��  �  ��  '  ��  '      B  , ,  �6  '  �6  �  ��  �  ��  '  �6  '      B  , ,  ��  '  ��  �  �4  �  �4  '  ��  '      B  , ,  ��  '  ��  �  ��  �  ��  '  ��  '      B  , ,  �2  '  �2  �  ��  �  ��  '  �2  '      B  , ,  ��  '  ��  �  �0  �  �0  '  ��  '      B  , ,  ��  '  ��  �  ��  �  ��  '  ��  '      B  , ,  �.  '  �.  �  ��  �  ��  '  �.  '      B  , ,  ��  '  ��  �  �,  �  �,  '  ��  '      B  , ,  ��  '  ��  �  ��  �  ��  '  ��  '      B  , ,  ��  '.  ��  '�  �U  '�  �U  '.  ��  '.      B  , ,  �*  '  �*  �  ��  �  ��  '  �*  '      B  , ,  �~  '  �~  �  �(  �  �(  '  �~  '      B  , ,  ��  '  ��  �  �|  �  �|  '  ��  '      B  , ,  �&  '  �&  �  ��  �  ��  '  �&  '      B  , ,  �z  '  �z  �  �$  �  �$  '  �z  '      B  , ,  ��  '  ��  �  �x  �  �x  '  ��  '      B  , ,  �"  '  �"  �  ��  �  ��  '  �"  '      B  , ,  �v  '  �v  �  �   �  �   '  �v  '      B  , ,  ��  '  ��  �  �t  �  �t  '  ��  '      B  , ,  �  '  �  �  ��  �  ��  '  �  '      B  , ,  �r  '  �r  �  �  �  �  '  �r  '      B  , ,  ��  '  ��  �  �p  �  �p  '  ��  '      B  , ,  ��  '.  ��  '�  �q  '�  �q  '.  ��  '.      B  , ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      B  , ,  �  '.  �  '�  ��  '�  ��  '.  �  '.      B  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      B  , ,  �F  �  �F  �  ��  �  ��  �  �F  �      B  , ,  ��  �  ��  �  �D  �  �D  �  ��  �      B  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      B  , ,  �B  �  �B  �  ��  �  ��  �  �B  �      B  , ,  ��  '  ��  �  ��  �  ��  '  ��  '      B  , ,  �N  '  �N  �  ��  �  ��  '  �N  '      B  , ,  ��  '  ��  �  �L  �  �L  '  ��  '      B  , ,  ��  '  ��  �  ��  �  ��  '  ��  '      B  , ,  �J  '  �J  �  ��  �  ��  '  �J  '      B  , ,  {  �  {  �  {�  �  {�  �  {  �      B  , ,  |V  �  |V  �  }   �  }   �  |V  �      B  , ,  }�  �  }�  �  ~T  �  ~T  �  }�  �      B  , ,  ~�  �  ~�  �  �  �  �  �  ~�  �      B  , ,  �R  �  �R  �  ��  �  ��  �  �R  �      B  , ,  ��  �  ��  �  �P  �  �P  �  ��  �      B  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      B  , ,  �J  �  �J  �  ��  �  ��  �  �J  �      B  , ,  s
  �  s
  �  s�  �  s�  �  s
  �      B  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      B  , ,  �N  �  �N  �  ��  �  ��  �  �N  �      B  , ,  ��  �  ��  �  �L  �  �L  �  ��  �      B  , ,  t^  �  t^  �  u  �  u  �  t^  �      B  , ,  u�  �  u�  �  v\  �  v\  �  u�  �      B  , ,  w  �  w  �  w�  �  w�  �  w  �      B  , ,  xZ  �  xZ  �  y  �  y  �  xZ  �      B  , ,  ]�  '  ]�  �  ^t  �  ^t  '  ]�  '      B  , ,  _  '  _  �  _�  �  _�  '  _  '      B  , ,  `r  '  `r  �  a  �  a  '  `r  '      B  , ,  a�  '  a�  �  bp  �  bp  '  a�  '      B  , ,  c  '  c  �  c�  �  c�  '  c  '      B  , ,  dn  '  dn  �  e  �  e  '  dn  '      B  , ,  y�  �  y�  �  zX  �  zX  �  y�  �      B  , ,  e�  '  e�  �  fl  �  fl  '  e�  '      B  , ,  g  '  g  �  g�  �  g�  '  g  '      B  , ,  hj  '  hj  �  i  �  i  '  hj  '      B  , ,  i�  '  i�  �  jh  �  jh  '  i�  '      B  , ,  k  '  k  �  k�  �  k�  '  k  '      B  , ,  lf  '  lf  �  m  �  m  '  lf  '      B  , ,  m�  '  m�  �  nd  �  nd  '  m�  '      B  , ,  o  '  o  �  o�  �  o�  '  o  '      B  , ,  pb  '  pb  �  q  �  q  '  pb  '      B  , ,  q�  '  q�  �  r`  �  r`  '  q�  '      B  , ,  s
  '  s
  �  s�  �  s�  '  s
  '      B  , ,  t^  '  t^  �  u  �  u  '  t^  '      B  , ,  u�  '  u�  �  v\  �  v\  '  u�  '      B  , ,  w  '  w  �  w�  �  w�  '  w  '      B  , ,  xZ  '  xZ  �  y  �  y  '  xZ  '      B  , ,  ]�  �  ]�  �  ^t  �  ^t  �  ]�  �      B  , ,  _  �  _  �  _�  �  _�  �  _  �      B  , ,  [�  )  [�  �  \b  �  \b  )  [�  )      B  , ,  `r  �  `r  �  a  �  a  �  `r  �      B  , ,  [�  �  [�    \b    \b  �  [�  �      B  , ,  a�  �  a�  �  bp  �  bp  �  a�  �      B  , ,  y�  '  y�  �  zX  �  zX  '  y�  '      B  , ,  {  '  {  �  {�  �  {�  '  {  '      B  , ,  |V  '  |V  �  }   �  }   '  |V  '      B  , ,  }�  '  }�  �  ~T  �  ~T  '  }�  '      B  , ,  c  �  c  �  c�  �  c�  �  c  �      B  , ,  ~�  '  ~�  �  �  �  �  '  ~�  '      B  , ,  dn  �  dn  �  e  �  e  �  dn  �      B  , ,  e�  �  e�  �  fl  �  fl  �  e�  �      B  , ,  g  �  g  �  g�  �  g�  �  g  �      B  , ,  hj  �  hj  �  i  �  i  �  hj  �      B  , ,  i�  �  i�  �  jh  �  jh  �  i�  �      B  , ,  k  �  k  �  k�  �  k�  �  k  �      B  , ,  lf  �  lf  �  m  �  m  �  lf  �      B  , ,  m�  �  m�  �  nd  �  nd  �  m�  �      B  , ,  o  �  o  �  o�  �  o�  �  o  �      B  , ,  pb  �  pb  �  q  �  q  �  pb  �      B  , ,  q�  �  q�  �  r`  �  r`  �  q�  �      B  , ,  �R  '  �R  �  ��  �  ��  '  �R  '      B  , ,  ��  '  ��  �  �P  �  �P  '  ��  '      B  , ,  r�  g  r�    sZ    sZ  g  r�  g      B  , ,  r�  c  r�    sZ    sZ  c  r�  c      B  , ,  r�    r�  �  sZ  �  sZ    r�        B  , ,  [�  9  [�  �  \b  �  \b  9  [�  9      B  , ,  _  �  _    _�    _�  �  _  �      B  , ,  ag  �  ag    b    b  �  ag  �      B  , ,  c�  �  c�    d_    d_  �  c�  �      B  , ,  f  �  f    f�    f�  �  f  �      B  , ,  hQ  �  hQ    h�    h�  �  hQ  �      B  , ,  j�  �  j�    kI    kI  �  j�  �      B  , ,  l�  �  l�    m�    m�  �  l�  �      B  , ,  o;  �  o;    o�    o�  �  o;  �      B  , ,  q�  �  q�    r3    r3  �  q�  �      B  , ,  s�  �  s�    t�    t�  �  s�  �      B  , ,  v%  �  v%    v�    v�  �  v%  �      B  , ,  xs  �  xs    y    y  �  xs  �      B  , ,  z�  �  z�    {k    {k  �  z�  �      B  , ,  }  �  }    }�    }�  �  }  �      B  , ,  ]  �  ]    �    �  �  ]  �      B  , ,  ��  �  ��    �U    �U  �  ��  �      B  , ,  ��  �  ��    ��    ��  �  ��  �      B  , ,  �G  �  �G    ��    ��  �  �G  �      B  , ,  ��  �  ��    �?    �?  �  ��  �      B  , ,  r�  _  r�  	  sZ  	  sZ  _  r�  _      B  , ,  r�    r�  �  sZ  �  sZ    r�        B  , ,  r�    r�  �  sZ  �  sZ    r�        B  , ,  r�  �  r�  a  sZ  a  sZ  �  r�  �      B  , ,  r�  �  r�  a  sZ  a  sZ  �  r�  �      B  , ,  r�  c  r�    sZ    sZ  c  r�  c      B  , ,  r�  �  r�  ]  sZ  ]  sZ  �  r�  �      B  , ,  r�     r�   �  sZ   �  sZ     r�         B  , ,  r�����  r����e  sZ���e  sZ����  r�����      B  , ,  r����g  r����  sZ���  sZ���g  r����g      B  , ,  r�  �  r�  e  sZ  e  sZ  �  r�  �      B  , ,  r����  r�����  sZ����  sZ���  r����      B  , ,  r�  _  r�  	  sZ  	  sZ  _  r�  _      B  , ,  ��    ��  �  �.  �  �.    ��        B  , ,  t�  g  t�    u�    u�  g  t�  g      B  , ,  wL  g  wL    w�    w�  g  wL  g      B  , ,  y�  g  y�    zD    zD  g  y�  g      B  , ,  {�  g  {�    |�    |�  g  {�  g      B  , ,  ~6  g  ~6    ~�    ~�  g  ~6  g      B  , ,  ��  g  ��    �.    �.  g  ��  g      B  , ,  ��  g  ��    �|    �|  g  ��  g      B  , ,  �   g  �     ��    ��  g  �   g      B  , ,  �n  g  �n    �    �  g  �n  g      B  , ,  ��    ��  �  �|  �  �|    ��        B  , ,  t�  c  t�    u�    u�  c  t�  c      B  , ,  wL  c  wL    w�    w�  c  wL  c      B  , ,  s�  	�  s�  
�  t�  
�  t�  	�  s�  	�      B  , ,  v%  	�  v%  
�  v�  
�  v�  	�  v%  	�      B  , ,  xs  	�  xs  
�  y  
�  y  	�  xs  	�      B  , ,  z�  	�  z�  
�  {k  
�  {k  	�  z�  	�      B  , ,  }  	�  }  
�  }�  
�  }�  	�  }  	�      B  , ,  ]  	�  ]  
�  �  
�  �  	�  ]  	�      B  , ,  t�    t�  �  u�  �  u�    t�        B  , ,  wL    wL  �  w�  �  w�    wL        B  , ,  ��  	�  ��  
�  �U  
�  �U  	�  ��  	�      B  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      B  , ,  t�    t�  �  u�  �  u�    t�        B  , ,  wL    wL  �  w�  �  w�    wL        B  , ,  y�    y�  �  zD  �  zD    y�        B  , ,  {�    {�  �  |�  �  |�    {�        B  , ,  ~6    ~6  �  ~�  �  ~�    ~6        B  , ,  ��    ��  �  �.  �  �.    ��        B  , ,  ��    ��  �  �|  �  �|    ��        B  , ,  �G  	�  �G  
�  ��  
�  ��  	�  �G  	�      B  , ,  �     �   �  ��  �  ��    �         B  , ,  �n    �n  �  �  �  �    �n        B  , ,  ��  	�  ��  
�  �?  
�  �?  	�  ��  	�      B  , ,  t�  �  t�  a  u�  a  u�  �  t�  �      B  , ,  wL  �  wL  a  w�  a  w�  �  wL  �      B  , ,  y�  �  y�  a  zD  a  zD  �  y�  �      B  , ,  {�  �  {�  a  |�  a  |�  �  {�  �      B  , ,  ~6  �  ~6  a  ~�  a  ~�  �  ~6  �      B  , ,  ��  �  ��  a  �.  a  �.  �  ��  �      B  , ,  y�  c  y�    zD    zD  c  y�  c      B  , ,  ��  �  ��  a  �|  a  �|  �  ��  �      B  , ,  �   �  �   a  ��  a  ��  �  �   �      B  , ,  {�  c  {�    |�    |�  c  {�  c      B  , ,  ~6  c  ~6    ~�    ~�  c  ~6  c      B  , ,  t�  �  t�  ]  u�  ]  u�  �  t�  �      B  , ,  wL  �  wL  ]  w�  ]  w�  �  wL  �      B  , ,  y�  �  y�  ]  zD  ]  zD  �  y�  �      B  , ,  {�  �  {�  ]  |�  ]  |�  �  {�  �      B  , ,  ~6  �  ~6  ]  ~�  ]  ~�  �  ~6  �      B  , ,  ��  �  ��  ]  �.  ]  �.  �  ��  �      B  , ,  ��  �  ��  ]  �|  ]  �|  �  ��  �      B  , ,  ��  c  ��    �.    �.  c  ��  c      B  , ,  �   �  �   ]  ��  ]  ��  �  �   �      B  , ,  �n  �  �n  ]  �  ]  �  �  �n  �      B  , ,  ��  c  ��    �|    �|  c  ��  c      B  , ,  �   c  �     ��    ��  c  �   c      B  , ,  �n  c  �n    �    �  c  �n  c      B  , ,  t�  �  t�  e  u�  e  u�  �  t�  �      B  , ,  wL  �  wL  e  w�  e  w�  �  wL  �      B  , ,  y�  �  y�  e  zD  e  zD  �  y�  �      B  , ,  {�  �  {�  e  |�  e  |�  �  {�  �      B  , ,  ~6  �  ~6  e  ~�  e  ~�  �  ~6  �      B  , ,  ��  �  ��  e  �.  e  �.  �  ��  �      B  , ,  ��  �  ��  e  �|  e  �|  �  ��  �      B  , ,  �   �  �   e  ��  e  ��  �  �   �      B  , ,  �n  �  �n  e  �  e  �  �  �n  �      B  , ,  �n  �  �n  a  �  a  �  �  �n  �      B  , ,  y�    y�  �  zD  �  zD    y�        B  , ,  �     �   �  ��  �  ��    �         B  , ,  {�    {�  �  |�  �  |�    {�        B  , ,  �n    �n  �  �  �  �    �n        B  , ,  t�  _  t�  	  u�  	  u�  _  t�  _      B  , ,  wL  _  wL  	  w�  	  w�  _  wL  _      B  , ,  y�  _  y�  	  zD  	  zD  _  y�  _      B  , ,  {�  _  {�  	  |�  	  |�  _  {�  _      B  , ,  ~6  _  ~6  	  ~�  	  ~�  _  ~6  _      B  , ,  ��  _  ��  	  �.  	  �.  _  ��  _      B  , ,  ��  _  ��  	  �|  	  �|  _  ��  _      B  , ,  �   _  �   	  ��  	  ��  _  �   _      B  , ,  �n  _  �n  	  �  	  �  _  �n  _      B  , ,  ~6    ~6  �  ~�  �  ~�    ~6        B  , ,  [�  5  [�  �  \b  �  \b  5  [�  5      B  , ,  ]�  g  ]�    ^�    ^�  g  ]�  g      B  , ,  `@  g  `@    `�    `�  g  `@  g      B  , ,  b�  g  b�    c8    c8  g  b�  g      B  , ,  d�  g  d�    e�    e�  g  d�  g      B  , ,  g*    g*  �  g�  �  g�    g*        B  , ,  [�  1  [�  �  \b  �  \b  1  [�  1      B  , ,  ]�  c  ]�    ^�    ^�  c  ]�  c      B  , ,  ix  �  ix  a  j"  a  j"  �  ix  �      B  , ,  k�  �  k�  a  lp  a  lp  �  k�  �      B  , ,  n  �  n  a  n�  a  n�  �  n  �      B  , ,  pb  �  pb  a  q  a  q  �  pb  �      B  , ,  `@  c  `@    `�    `�  c  `@  c      B  , ,  b�  c  b�    c8    c8  c  b�  c      B  , ,  ix    ix  �  j"  �  j"    ix        B  , ,  k�    k�  �  lp  �  lp    k�        B  , ,  n    n  �  n�  �  n�    n        B  , ,  pb    pb  �  q  �  q    pb        B  , ,  d�  c  d�    e�    e�  c  d�  c      B  , ,  g*  c  g*    g�    g�  c  g*  c      B  , ,  ix  c  ix    j"    j"  c  ix  c      B  , ,  k�  c  k�    lp    lp  c  k�  c      B  , ,  [�  �  [�  3  \b  3  \b  �  [�  �      B  , ,  ]�  �  ]�  e  ^�  e  ^�  �  ]�  �      B  , ,  `@  �  `@  e  `�  e  `�  �  `@  �      B  , ,  b�  �  b�  e  c8  e  c8  �  b�  �      B  , ,  d�  �  d�  e  e�  e  e�  �  d�  �      B  , ,  [�  �  [�  +  \b  +  \b  �  [�  �      B  , ,  ]�  �  ]�  ]  ^�  ]  ^�  �  ]�  �      B  , ,  `@  �  `@  ]  `�  ]  `�  �  `@  �      B  , ,  b�  �  b�  ]  c8  ]  c8  �  b�  �      B  , ,  d�  �  d�  ]  e�  ]  e�  �  d�  �      B  , ,  g*  �  g*  ]  g�  ]  g�  �  g*  �      B  , ,  n  c  n    n�    n�  c  n  c      B  , ,  g*  �  g*  e  g�  e  g�  �  g*  �      B  , ,  ix  �  ix  ]  j"  ]  j"  �  ix  �      B  , ,  k�  �  k�  ]  lp  ]  lp  �  k�  �      B  , ,  n  �  n  ]  n�  ]  n�  �  n  �      B  , ,  pb  �  pb  ]  q  ]  q  �  pb  �      B  , ,  pb  c  pb    q    q  c  pb  c      B  , ,  g*  g  g*    g�    g�  g  g*  g      B  , ,  ix  g  ix    j"    j"  g  ix  g      B  , ,  [�  
�  [�  �  \b  �  \b  
�  [�  
�      B  , ,  k�  g  k�    lp    lp  g  k�  g      B  , ,  [�  	�  [�  
7  \b  
7  \b  	�  [�  	�      B  , ,  _  	�  _  
�  _�  
�  _�  	�  _  	�      B  , ,  ag  	�  ag  
�  b  
�  b  	�  ag  	�      B  , ,  c�  	�  c�  
�  d_  
�  d_  	�  c�  	�      B  , ,  ix  �  ix  e  j"  e  j"  �  ix  �      B  , ,  f  	�  f  
�  f�  
�  f�  	�  f  	�      B  , ,  hQ  	�  hQ  
�  h�  
�  h�  	�  hQ  	�      B  , ,  k�  �  k�  e  lp  e  lp  �  k�  �      B  , ,  j�  	�  j�  
�  kI  
�  kI  	�  j�  	�      B  , ,  n  �  n  e  n�  e  n�  �  n  �      B  , ,  pb  �  pb  e  q  e  q  �  pb  �      B  , ,  l�  	�  l�  
�  m�  
�  m�  	�  l�  	�      B  , ,  o;  	�  o;  
�  o�  
�  o�  	�  o;  	�      B  , ,  q�  	�  q�  
�  r3  
�  r3  	�  q�  	�      B  , ,  n  g  n    n�    n�  g  n  g      B  , ,  pb  g  pb    q    q  g  pb  g      B  , ,  [�  �  [�  �  \b  �  \b  �  [�  �      B  , ,  [�  �  [�  /  \b  /  \b  �  [�  �      B  , ,  ]�  �  ]�  a  ^�  a  ^�  �  ]�  �      B  , ,  `@  �  `@  a  `�  a  `�  �  `@  �      B  , ,  b�  �  b�  a  c8  a  c8  �  b�  �      B  , ,  d�  �  d�  a  e�  a  e�  �  d�  �      B  , ,  g*  �  g*  a  g�  a  g�  �  g*  �      B  , ,  [�  �  [�  �  \b  �  \b  �  [�  �      B  , ,  [�  -  [�  �  \b  �  \b  -  [�  -      B  , ,  ]�    ]�  �  ^�  �  ^�    ]�        B  , ,  `@    `@  �  `�  �  `�    `@        B  , ,  ]�  _  ]�  	  ^�  	  ^�  _  ]�  _      B  , ,  `@  _  `@  	  `�  	  `�  _  `@  _      B  , ,  b�  _  b�  	  c8  	  c8  _  b�  _      B  , ,  d�  _  d�  	  e�  	  e�  _  d�  _      B  , ,  g*  _  g*  	  g�  	  g�  _  g*  _      B  , ,  ix  _  ix  	  j"  	  j"  _  ix  _      B  , ,  k�  _  k�  	  lp  	  lp  _  k�  _      B  , ,  n  _  n  	  n�  	  n�  _  n  _      B  , ,  pb  _  pb  	  q  	  q  _  pb  _      B  , ,  b�    b�  �  c8  �  c8    b�        B  , ,  d�    d�  �  e�  �  e�    d�        B  , ,  ]�    ]�  �  ^�  �  ^�    ]�        B  , ,  g*    g*  �  g�  �  g�    g*        B  , ,  ix    ix  �  j"  �  j"    ix        B  , ,  k�    k�  �  lp  �  lp    k�        B  , ,  n    n  �  n�  �  n�    n        B  , ,  pb    pb  �  q  �  q    pb        B  , ,  `@    `@  �  `�  �  `�    `@        B  , ,  b�    b�  �  c8  �  c8    b�        B  , ,  d�    d�  �  e�  �  e�    d�        B  , ,  b�     b�   �  c8   �  c8     b�         B  , ,  d�     d�   �  e�   �  e�     d�         B  , ,  g*     g*   �  g�   �  g�     g*         B  , ,  ix     ix   �  j"   �  j"     ix         B  , ,  k�     k�   �  lp   �  lp     k�         B  , ,  n     n   �  n�   �  n�     n         B  , ,  pb     pb   �  q   �  q     pb         B  , ,  k�  �  k�  a  lp  a  lp  �  k�  �      B  , ,  n  �  n  a  n�  a  n�  �  n  �      B  , ,  pb  �  pb  a  q  a  q  �  pb  �      B  , ,  b�    b�  �  c8  �  c8    b�        B  , ,  d�    d�  �  e�  �  e�    d�        B  , ,  [�����  [�����  \b����  \b����  [�����      B  , ,  ]�����  ]����e  ^����e  ^�����  ]�����      B  , ,  `@����  `@���e  `����e  `�����  `@����      B  , ,  b�����  b����e  c8���e  c8����  b�����      B  , ,  d�����  d����e  e����e  e�����  d�����      B  , ,  g*����  g*���e  g����e  g�����  g*����      B  , ,  ix����  ix���e  j"���e  j"����  ix����      B  , ,  k�����  k����e  lp���e  lp����  k�����      B  , ,  n����  n���e  n����e  n�����  n����      B  , ,  pb����  pb���e  q���e  q����  pb����      B  , ,  g*    g*  �  g�  �  g�    g*        B  , ,  ix    ix  �  j"  �  j"    ix        B  , ,  k�    k�  �  lp  �  lp    k�        B  , ,  [�����  [����C  \b���C  \b����  [�����      B  , ,  ]����g  ]����  ^����  ^����g  ]����g      B  , ,  `@���g  `@���  `����  `����g  `@���g      B  , ,  b����g  b����  c8���  c8���g  b����g      B  , ,  d����g  d����  e����  e����g  d����g      B  , ,  g*���g  g*���  g����  g����g  g*���g      B  , ,  ix���g  ix���  j"���  j"���g  ix���g      B  , ,  k����g  k����  lp���  lp���g  k����g      B  , ,  n���g  n���  n����  n����g  n���g      B  , ,  pb���g  pb���  q���  q���g  pb���g      B  , ,  n    n  �  n�  �  n�    n        B  , ,  pb    pb  �  q  �  q    pb        B  , ,  `@  _  `@  	  `�  	  `�  _  `@  _      B  , ,  b�  _  b�  	  c8  	  c8  _  b�  _      B  , ,  d�  _  d�  	  e�  	  e�  _  d�  _      B  , ,  g*  _  g*  	  g�  	  g�  _  g*  _      B  , ,  ix  _  ix  	  j"  	  j"  _  ix  _      B  , ,  k�  _  k�  	  lp  	  lp  _  k�  _      B  , ,  n  _  n  	  n�  	  n�  _  n  _      B  , ,  [�  �  [�  ?  \b  ?  \b  �  [�  �      B  , ,  ]�  c  ]�    ^�    ^�  c  ]�  c      B  , ,  `@  c  `@    `�    `�  c  `@  c      B  , ,  b�  c  b�    c8    c8  c  b�  c      B  , ,  d�  c  d�    e�    e�  c  d�  c      B  , ,  [����E  [�����  \b����  \b���E  [����E      B  , ,  ]����  ]�����  ^�����  ^����  ]����      B  , ,  `@���  `@����  `�����  `����  `@���      B  , ,  b����  b�����  c8����  c8���  b����      B  , ,  d����  d�����  e�����  e����  d����      B  , ,  g*���  g*����  g�����  g����  g*���      B  , ,  ix���  ix����  j"����  j"���  ix���      B  , ,  k����  k�����  lp����  lp���  k����      B  , ,  n���  n����  n�����  n����  n���      B  , ,  pb���  pb����  q����  q���  pb���      B  , ,  g*  c  g*    g�    g�  c  g*  c      B  , ,  ix  c  ix    j"    j"  c  ix  c      B  , ,  k�  c  k�    lp    lp  c  k�  c      B  , ,  n  c  n    n�    n�  c  n  c      B  , ,  pb  c  pb    q    q  c  pb  c      B  , ,  pb  _  pb  	  q  	  q  _  pb  _      B  , ,  [�  �  [�  �  \b  �  \b  �  [�  �      B  , ,  [�  �  [�  ;  \b  ;  \b  �  [�  �      B  , ,  ]�  _  ]�  	  ^�  	  ^�  _  ]�  _      B  , ,  [�  =  [�  �  \b  �  \b  =  [�  =      B  , ,  ]�    ]�  �  ^�  �  ^�    ]�        B  , ,  `@    `@  �  `�  �  `�    `@        B  , ,  [�  �  [�  �  \b  �  \b  �  [�  �      B  , ,  ]�  �  ]�  a  ^�  a  ^�  �  ]�  �      B  , ,  [�����  [�����  \b����  \b����  [�����      B  , ,  `@  �  `@  a  `�  a  `�  �  `@  �      B  , ,  b�  �  b�  a  c8  a  c8  �  b�  �      B  , ,  d�  �  d�  a  e�  a  e�  �  d�  �      B  , ,  g*  �  g*  a  g�  a  g�  �  g*  �      B  , ,  ix  �  ix  a  j"  a  j"  �  ix  �      B  , ,  [�   A  [�   �  \b   �  \b   A  [�   A      B  , ,  ]�     ]�   �  ^�   �  ^�     ]�         B  , ,  `@     `@   �  `�   �  `�     `@         B  , ,  y�    y�  �  zD  �  zD    y�        B  , ,  {�    {�  �  |�  �  |�    {�        B  , ,  ~6    ~6  �  ~�  �  ~�    ~6        B  , ,  ��    ��  �  �.  �  �.    ��        B  , ,  ��    ��  �  �|  �  �|    ��        B  , ,  �     �   �  ��  �  ��    �         B  , ,  �n    �n  �  �  �  �    �n        B  , ,  ��  _  ��  	  �|  	  �|  _  ��  _      B  , ,  t����g  t����  u����  u����g  t����g      B  , ,  wL���g  wL���  w����  w����g  wL���g      B  , ,  y����g  y����  zD���  zD���g  y����g      B  , ,  {����g  {����  |����  |����g  {����g      B  , ,  ~6���g  ~6���  ~����  ~����g  ~6���g      B  , ,  �����g  �����  �.���  �.���g  �����g      B  , ,  �����g  �����  �|���  �|���g  �����g      B  , ,  � ���g  � ���  �����  �����g  � ���g      B  , ,  �n���g  �n���  ����  ����g  �n���g      B  , ,  �   _  �   	  ��  	  ��  _  �   _      B  , ,  �n  _  �n  	  �  	  �  _  �n  _      B  , ,  t�  _  t�  	  u�  	  u�  _  t�  _      B  , ,  wL  _  wL  	  w�  	  w�  _  wL  _      B  , ,  y�  _  y�  	  zD  	  zD  _  y�  _      B  , ,  t�  �  t�  a  u�  a  u�  �  t�  �      B  , ,  wL  �  wL  a  w�  a  w�  �  wL  �      B  , ,  y�  �  y�  a  zD  a  zD  �  y�  �      B  , ,  t�     t�   �  u�   �  u�     t�         B  , ,  wL     wL   �  w�   �  w�     wL         B  , ,  y�     y�   �  zD   �  zD     y�         B  , ,  {�     {�   �  |�   �  |�     {�         B  , ,  ~6     ~6   �  ~�   �  ~�     ~6         B  , ,  ��     ��   �  �.   �  �.     ��         B  , ,  ��     ��   �  �|   �  �|     ��         B  , ,  �      �    �  ��   �  ��     �          B  , ,  �n     �n   �  �   �  �     �n         B  , ,  {�  �  {�  a  |�  a  |�  �  {�  �      B  , ,  ~6  �  ~6  a  ~�  a  ~�  �  ~6  �      B  , ,  ��  �  ��  a  �.  a  �.  �  ��  �      B  , ,  t�  c  t�    u�    u�  c  t�  c      B  , ,  wL  c  wL    w�    w�  c  wL  c      B  , ,  y�  c  y�    zD    zD  c  y�  c      B  , ,  {�  c  {�    |�    |�  c  {�  c      B  , ,  t����  t�����  u�����  u����  t����      B  , ,  wL���  wL����  w�����  w����  wL���      B  , ,  y����  y�����  zD����  zD���  y����      B  , ,  {����  {�����  |�����  |����  {����      B  , ,  ~6���  ~6����  ~�����  ~����  ~6���      B  , ,  �����  ������  �.����  �.���  �����      B  , ,  �����  ������  �|����  �|���  �����      B  , ,  � ���  � ����  ������  �����  � ���      B  , ,  �n���  �n����  �����  ����  �n���      B  , ,  ~6  c  ~6    ~�    ~�  c  ~6  c      B  , ,  ��  c  ��    �.    �.  c  ��  c      B  , ,  ��  c  ��    �|    �|  c  ��  c      B  , ,  �   c  �     ��    ��  c  �   c      B  , ,  �n  c  �n    �    �  c  �n  c      B  , ,  ��  �  ��  a  �|  a  �|  �  ��  �      B  , ,  �   �  �   a  ��  a  ��  �  �   �      B  , ,  �n  �  �n  a  �  a  �  �  �n  �      B  , ,  t�����  t����e  u����e  u�����  t�����      B  , ,  wL����  wL���e  w����e  w�����  wL����      B  , ,  y�����  y����e  zD���e  zD����  y�����      B  , ,  {�����  {����e  |����e  |�����  {�����      B  , ,  ~6����  ~6���e  ~����e  ~�����  ~6����      B  , ,  ������  �����e  �.���e  �.����  ������      B  , ,  ������  �����e  �|���e  �|����  ������      B  , ,  � ����  � ���e  �����e  ������  � ����      B  , ,  �n����  �n���e  ����e  �����  �n����      B  , ,  {�  _  {�  	  |�  	  |�  _  {�  _      B  , ,  ~6  _  ~6  	  ~�  	  ~�  _  ~6  _      B  , ,  ��  _  ��  	  �.  	  �.  _  ��  _      B  , ,  t�    t�  �  u�  �  u�    t�        B  , ,  wL    wL  �  w�  �  w�    wL        B  , ,  ��    ��  �  �r  �  �r    ��        B  , ,  ��    ��  �  �r  �  �r    ��        B  , ,  ��  �  ��  a  �r  a  �r  �  ��  �      B  , ,  ��  _  ��  	  �r  	  �r  _  ��  _      B  , ,  ��  c  ��    �r    �r  c  ��  c      B  , ,  ��    ��  �  �r  �  �r    ��        B  , ,  ��  �  ��    ��    ��  �  ��  �      B  , ,  �1  �  �1    ��    ��  �  �1  �      B  , ,  �  �  �    �)    �)  �  �  �      B  , ,  ��  �  ��    �w    �w  �  ��  �      B  , ,  �  �  �    ��    ��  �  �  �      B  , ,  �i  �  �i    �    �  �  �i  �      B  , ,  ��  �  ��    �a    �a  �  ��  �      B  , ,  �  �  �    ��    ��  �  �  �      B  , ,  �S  �  �S    ��    ��  �  �S  �      B  , ,  ��  �  ��    �K    �K  �  ��  �      B  , ,  ��     ��   �  �r   �  �r     ��         B  , ,  ��  �  ��    ��    ��  �  ��  �      B  , ,  �=  �  �=    ��    ��  �  �=  �      B  , ,  ��  �  ��    �5    �5  �  ��  �      B  , ,  ��  �  ��    ��    ��  �  ��  �      B  , ,  �'  �  �'    ��    ��  �  �'  �      B  , ,  �u  �  �u    �    �  �  �u  �      B  , ,  ��  �  ��    �m    �m  �  ��  �      B  , ,  �  �  �    ��    ��  �  �  �      B  , ,  �_  �  �_    �	    �	  �  �_  �      B  , ,  ��  �  ��    �W    �W  �  ��  �      B  , ,  ��  �  ��  e  �r  e  �r  �  ��  �      B  , ,  ������  �����e  �r���e  �r����  ������      B  , ,  ��  �  ��  ]  �r  ]  �r  �  ��  �      B  , ,  ��  c  ��    �r    �r  c  ��  c      B  , ,  �����g  �����  �r���  �r���g  �����g      B  , ,  ��  _  ��  	  �r  	  �r  _  ��  _      B  , ,  ��  �  ��  a  �r  a  �r  �  ��  �      B  , ,  �����  ������  �r����  �r���  �����      B  , ,  ��  g  ��    �r    �r  g  ��  g      B  , ,  ��  _  ��  	  �\  	  �\  _  ��  _      B  , ,  �   _  �   	  ��  	  ��  _  �   _      B  , ,  �N  _  �N  	  ��  	  ��  _  �N  _      B  , ,  ��  _  ��  	  �F  	  �F  _  ��  _      B  , ,  ��  _  ��  	  ��  	  ��  _  ��  _      B  , ,  �8  _  �8  	  ��  	  ��  _  �8  _      B  , ,  ��  _  ��  	  �0  	  �0  _  ��  _      B  , ,  ��  �  ��  a  �0  a  �0  �  ��  �      B  , ,  ��  �  ��  a  �~  a  �~  �  ��  �      B  , ,  �    �  �  ��  �  ��    �        B  , ,  �d    �d  �  �  �  �    �d        B  , ,  ��    ��  �  ��  �  ��    ��        B  , ,  �8    �8  �  ��  �  ��    �8        B  , ,  ��    ��  �  �0  �  �0    ��        B  , ,  ��    ��  �  �~  �  �~    ��        B  , ,  ��  _  ��  	  �~  	  �~  _  ��  _      B  , ,  �8  g  �8    ��    ��  g  �8  g      B  , ,  �    �  �  ��  �  ��    �        B  , ,  �d    �d  �  �  �  �    �d        B  , ,  ��    ��  �  �\  �  �\    ��        B  , ,  �     �   �  ��  �  ��    �         B  , ,  �N    �N  �  ��  �  ��    �N        B  , ,  ��    ��  �  �F  �  �F    ��        B  , ,  ��    ��  �  ��  �  ��    ��        B  , ,  �8    �8  �  ��  �  ��    �8        B  , ,  ��    ��  �  �0  �  �0    ��        B  , ,  ��  g  ��    �0    �0  g  ��  g      B  , ,  ��    ��  �  �~  �  �~    ��        B  , ,  ��  g  ��    �~    �~  g  ��  g      B  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      B  , ,  �=  	�  �=  
�  ��  
�  ��  	�  �=  	�      B  , ,  ��  	�  ��  
�  �5  
�  �5  	�  ��  	�      B  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      B  , ,  �  �  �  e  ��  e  ��  �  �  �      B  , ,  �d  �  �d  e  �  e  �  �  �d  �      B  , ,  ��  �  ��  e  �\  e  �\  �  ��  �      B  , ,  �   �  �   e  ��  e  ��  �  �   �      B  , ,  �N  �  �N  e  ��  e  ��  �  �N  �      B  , ,  ��  �  ��  e  �F  e  �F  �  ��  �      B  , ,  �'  	�  �'  
�  ��  
�  ��  	�  �'  	�      B  , ,  �u  	�  �u  
�  �  
�  �  	�  �u  	�      B  , ,  �  �  �  ]  ��  ]  ��  �  �  �      B  , ,  �d  �  �d  ]  �  ]  �  �  �d  �      B  , ,  ��  �  ��  ]  �\  ]  �\  �  ��  �      B  , ,  �   �  �   ]  ��  ]  ��  �  �   �      B  , ,  �N  �  �N  ]  ��  ]  ��  �  �N  �      B  , ,  ��  �  ��  ]  �F  ]  �F  �  ��  �      B  , ,  ��  �  ��  ]  ��  ]  ��  �  ��  �      B  , ,  �8  �  �8  ]  ��  ]  ��  �  �8  �      B  , ,  ��  �  ��  ]  �0  ]  �0  �  ��  �      B  , ,  ��  �  ��  ]  �~  ]  �~  �  ��  �      B  , ,  ��  �  ��  e  ��  e  ��  �  ��  �      B  , ,  �8  �  �8  e  ��  e  ��  �  �8  �      B  , ,  ��  �  ��  e  �0  e  �0  �  ��  �      B  , ,  ��  �  ��  e  �~  e  �~  �  ��  �      B  , ,  ��  	�  ��  
�  �m  
�  �m  	�  ��  	�      B  , ,  �  c  �    ��    ��  c  �  c      B  , ,  �d  c  �d    �    �  c  �d  c      B  , ,  ��  c  ��    �\    �\  c  ��  c      B  , ,  �   c  �     ��    ��  c  �   c      B  , ,  �N  c  �N    ��    ��  c  �N  c      B  , ,  ��  c  ��    �F    �F  c  ��  c      B  , ,  ��  c  ��    ��    ��  c  ��  c      B  , ,  �8  c  �8    ��    ��  c  �8  c      B  , ,  ��  c  ��    �0    �0  c  ��  c      B  , ,  ��  c  ��    �~    �~  c  ��  c      B  , ,  ��    ��  �  �\  �  �\    ��        B  , ,  �     �   �  ��  �  ��    �         B  , ,  �N    �N  �  ��  �  ��    �N        B  , ,  ��    ��  �  �F  �  �F    ��        B  , ,  �  	�  �  
�  ��  
�  ��  	�  �  	�      B  , ,  �_  	�  �_  
�  �	  
�  �	  	�  �_  	�      B  , ,  ��  	�  ��  
�  �W  
�  �W  	�  ��  	�      B  , ,  �  �  �  a  ��  a  ��  �  �  �      B  , ,  �d  �  �d  a  �  a  �  �  �d  �      B  , ,  ��  �  ��  a  �\  a  �\  �  ��  �      B  , ,  �   �  �   a  ��  a  ��  �  �   �      B  , ,  �N  �  �N  a  ��  a  ��  �  �N  �      B  , ,  ��  �  ��  a  �F  a  �F  �  ��  �      B  , ,  �  _  �  	  ��  	  ��  _  �  _      B  , ,  ��  �  ��  a  ��  a  ��  �  ��  �      B  , ,  �8  �  �8  a  ��  a  ��  �  �8  �      B  , ,  �d  _  �d  	  �  	  �  _  �d  _      B  , ,  �  g  �    ��    ��  g  �  g      B  , ,  �d  g  �d    �    �  g  �d  g      B  , ,  ��  g  ��    �\    �\  g  ��  g      B  , ,  �   g  �     ��    ��  g  �   g      B  , ,  �N  g  �N    ��    ��  g  �N  g      B  , ,  ��  g  ��    �F    �F  g  ��  g      B  , ,  ��  g  ��    ��    ��  g  ��  g      B  , ,  ��  �  ��  e  ��  e  ��  �  ��  �      B  , ,  �,  �  �,  e  ��  e  ��  �  �,  �      B  , ,  �z  �  �z  e  �$  e  �$  �  �z  �      B  , ,  �  	�  �  
�  ��  
�  ��  	�  �  	�      B  , ,  �
    �
  �  ��  �  ��    �
        B  , ,  �X    �X  �  �  �  �    �X        B  , ,  ��    ��  �  �P  �  �P    ��        B  , ,  ��    ��  �  ��  �  ��    ��        B  , ,  �B    �B  �  ��  �  ��    �B        B  , ,  ��    ��  �  �:  �  �:    ��        B  , ,  ��    ��  �  ��  �  ��    ��        B  , ,  �,    �,  �  ��  �  ��    �,        B  , ,  �z    �z  �  �$  �  �$    �z        B  , ,  �i  	�  �i  
�  �  
�  �  	�  �i  	�      B  , ,  ��  	�  ��  
�  �a  
�  �a  	�  ��  	�      B  , ,  �  	�  �  
�  ��  
�  ��  	�  �  	�      B  , ,  �
  c  �
    ��    ��  c  �
  c      B  , ,  �X  c  �X    �    �  c  �X  c      B  , ,  ��  c  ��    �P    �P  c  ��  c      B  , ,  ��  c  ��    ��    ��  c  ��  c      B  , ,  �B  c  �B    ��    ��  c  �B  c      B  , ,  ��  c  ��    �:    �:  c  ��  c      B  , ,  ��  c  ��    ��    ��  c  ��  c      B  , ,  �,  c  �,    ��    ��  c  �,  c      B  , ,  �z  c  �z    �$    �$  c  �z  c      B  , ,  �
  �  �
  e  ��  e  ��  �  �
  �      B  , ,  �X  �  �X  e  �  e  �  �  �X  �      B  , ,  �S  	�  �S  
�  ��  
�  ��  	�  �S  	�      B  , ,  ��  	�  ��  
�  �K  
�  �K  	�  ��  	�      B  , ,  ��  _  ��  	  ��  	  ��  _  ��  _      B  , ,  �B  _  �B  	  ��  	  ��  _  �B  _      B  , ,  ��  _  ��  	  �:  	  �:  _  ��  _      B  , ,  ��  _  ��  	  ��  	  ��  _  ��  _      B  , ,  �
    �
  �  ��  �  ��    �
        B  , ,  �X    �X  �  �  �  �    �X        B  , ,  ��    ��  �  �P  �  �P    ��        B  , ,  ��    ��  �  ��  �  ��    ��        B  , ,  �B    �B  �  ��  �  ��    �B        B  , ,  ��    ��  �  �:  �  �:    ��        B  , ,  ��    ��  �  ��  �  ��    ��        B  , ,  �,    �,  �  ��  �  ��    �,        B  , ,  �
  �  �
  a  ��  a  ��  �  �
  �      B  , ,  �X  �  �X  a  �  a  �  �  �X  �      B  , ,  �
  �  �
  ]  ��  ]  ��  �  �
  �      B  , ,  �X  �  �X  ]  �  ]  �  �  �X  �      B  , ,  ��  �  ��  a  �P  a  �P  �  ��  �      B  , ,  ��  �  ��  a  ��  a  ��  �  ��  �      B  , ,  �B  �  �B  a  ��  a  ��  �  �B  �      B  , ,  ��  �  ��  a  �:  a  �:  �  ��  �      B  , ,  ��  �  ��  a  ��  a  ��  �  ��  �      B  , ,  �,  �  �,  a  ��  a  ��  �  �,  �      B  , ,  �z  �  �z  a  �$  a  �$  �  �z  �      B  , ,  ��  �  ��  ]  �P  ]  �P  �  ��  �      B  , ,  ��  �  ��  ]  ��  ]  ��  �  ��  �      B  , ,  �B  �  �B  ]  ��  ]  ��  �  �B  �      B  , ,  ��  �  ��  ]  �:  ]  �:  �  ��  �      B  , ,  ��  �  ��  ]  ��  ]  ��  �  ��  �      B  , ,  �,  �  �,  ]  ��  ]  ��  �  �,  �      B  , ,  �z  �  �z  ]  �$  ]  �$  �  �z  �      B  , ,  �,  _  �,  	  ��  	  ��  _  �,  _      B  , ,  �z  _  �z  	  �$  	  �$  _  �z  _      B  , ,  �z    �z  �  �$  �  �$    �z        B  , ,  �
  g  �
    ��    ��  g  �
  g      B  , ,  �X  g  �X    �    �  g  �X  g      B  , ,  ��  g  ��    �P    �P  g  ��  g      B  , ,  ��  g  ��    ��    ��  g  ��  g      B  , ,  �B  g  �B    ��    ��  g  �B  g      B  , ,  ��  g  ��    �:    �:  g  ��  g      B  , ,  ��  g  ��    ��    ��  g  ��  g      B  , ,  �,  g  �,    ��    ��  g  �,  g      B  , ,  �z  g  �z    �$    �$  g  �z  g      B  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      B  , ,  �1  	�  �1  
�  ��  
�  ��  	�  �1  	�      B  , ,  �  	�  �  
�  �)  
�  �)  	�  �  	�      B  , ,  ��  	�  ��  
�  �w  
�  �w  	�  ��  	�      B  , ,  ��  �  ��  e  �P  e  �P  �  ��  �      B  , ,  ��  �  ��  e  ��  e  ��  �  ��  �      B  , ,  �B  �  �B  e  ��  e  ��  �  �B  �      B  , ,  ��  �  ��  e  �:  e  �:  �  ��  �      B  , ,  �
  _  �
  	  ��  	  ��  _  �
  _      B  , ,  �X  _  �X  	  �  	  �  _  �X  _      B  , ,  ��  _  ��  	  �P  	  �P  _  ��  _      B  , ,  �B     �B   �  ��   �  ��     �B         B  , ,  ��     ��   �  �:   �  �:     ��         B  , ,  ��     ��   �  ��   �  ��     ��         B  , ,  �,     �,   �  ��   �  ��     �,         B  , ,  �
  _  �
  	  ��  	  ��  _  �
  _      B  , ,  �
���g  �
���  �����  �����g  �
���g      B  , ,  �X���g  �X���  ����  ����g  �X���g      B  , ,  �����g  �����  �P���  �P���g  �����g      B  , ,  �����g  �����  �����  �����g  �����g      B  , ,  �B���g  �B���  �����  �����g  �B���g      B  , ,  �����g  �����  �:���  �:���g  �����g      B  , ,  �����g  �����  �����  �����g  �����g      B  , ,  �,���g  �,���  �����  �����g  �,���g      B  , ,  �z���g  �z���  �$���  �$���g  �z���g      B  , ,  �z     �z   �  �$   �  �$     �z         B  , ,  �X  _  �X  	  �  	  �  _  �X  _      B  , ,  ��  _  ��  	  �P  	  �P  _  ��  _      B  , ,  ��  _  ��  	  ��  	  ��  _  ��  _      B  , ,  �B  _  �B  	  ��  	  ��  _  �B  _      B  , ,  ��  _  ��  	  �:  	  �:  _  ��  _      B  , ,  ��  _  ��  	  ��  	  ��  _  ��  _      B  , ,  �,  _  �,  	  ��  	  ��  _  �,  _      B  , ,  �z  _  �z  	  �$  	  �$  _  �z  _      B  , ,  �
����  �
���e  �����e  ������  �
����      B  , ,  �X����  �X���e  ����e  �����  �X����      B  , ,  ������  �����e  �P���e  �P����  ������      B  , ,  ������  �����e  �����e  ������  ������      B  , ,  �B����  �B���e  �����e  ������  �B����      B  , ,  ������  �����e  �:���e  �:����  ������      B  , ,  ������  �����e  �����e  ������  ������      B  , ,  �,����  �,���e  �����e  ������  �,����      B  , ,  �z����  �z���e  �$���e  �$����  �z����      B  , ,  �B  �  �B  a  ��  a  ��  �  �B  �      B  , ,  ��  �  ��  a  �:  a  �:  �  ��  �      B  , ,  ��  �  ��  a  ��  a  ��  �  ��  �      B  , ,  �,  �  �,  a  ��  a  ��  �  �,  �      B  , ,  �z  �  �z  a  �$  a  �$  �  �z  �      B  , ,  �z    �z  �  �$  �  �$    �z        B  , ,  �
���  �
����  ������  �����  �
���      B  , ,  �X���  �X����  �����  ����  �X���      B  , ,  �����  ������  �P����  �P���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �B���  �B����  ������  �����  �B���      B  , ,  �����  ������  �:����  �:���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �,���  �,����  ������  �����  �,���      B  , ,  �z���  �z����  �$����  �$���  �z���      B  , ,  ��    ��  �  �P  �  �P    ��        B  , ,  �
  c  �
    ��    ��  c  �
  c      B  , ,  �X  c  �X    �    �  c  �X  c      B  , ,  ��  c  ��    �P    �P  c  ��  c      B  , ,  ��  c  ��    ��    ��  c  ��  c      B  , ,  �B  c  �B    ��    ��  c  �B  c      B  , ,  ��  c  ��    �:    �:  c  ��  c      B  , ,  ��  c  ��    ��    ��  c  ��  c      B  , ,  �,  c  �,    ��    ��  c  �,  c      B  , ,  �z  c  �z    �$    �$  c  �z  c      B  , ,  ��    ��  �  ��  �  ��    ��        B  , ,  �B    �B  �  ��  �  ��    �B        B  , ,  ��    ��  �  �:  �  �:    ��        B  , ,  ��    ��  �  ��  �  ��    ��        B  , ,  �,    �,  �  ��  �  ��    �,        B  , ,  �
  �  �
  a  ��  a  ��  �  �
  �      B  , ,  �X  �  �X  a  �  a  �  �  �X  �      B  , ,  ��  �  ��  a  �P  a  �P  �  ��  �      B  , ,  ��  �  ��  a  ��  a  ��  �  ��  �      B  , ,  �
     �
   �  ��   �  ��     �
         B  , ,  �
    �
  �  ��  �  ��    �
        B  , ,  �X    �X  �  �  �  �    �X        B  , ,  �X     �X   �  �   �  �     �X         B  , ,  ��     ��   �  �P   �  �P     ��         B  , ,  ��     ��   �  ��   �  ��     ��         B  , ,  �8���g  �8���  �����  �����g  �8���g      B  , ,  �����g  �����  �0���  �0���g  �����g      B  , ,  �����g  �����  �~���  �~���g  �����g      B  , ,  � ����  � ���e  �����e  ������  � ����      B  , ,  �N����  �N���e  �����e  ������  �N����      B  , ,  ������  �����e  �F���e  �F����  ������      B  , ,  ������  �����e  �����e  ������  ������      B  , ,  �8����  �8���e  �����e  ������  �8����      B  , ,  ������  �����e  �0���e  �0����  ������      B  , ,  ������  �����e  �~���e  �~����  ������      B  , ,  ��  �  ��  a  �~  a  �~  �  ��  �      B  , ,  �     �   �  ��  �  ��    �         B  , ,  �  _  �  	  ��  	  ��  _  �  _      B  , ,  �d  _  �d  	  �  	  �  _  �d  _      B  , ,  ��  _  ��  	  �\  	  �\  _  ��  _      B  , ,  �   _  �   	  ��  	  ��  _  �   _      B  , ,  �N  _  �N  	  ��  	  ��  _  �N  _      B  , ,  ��  _  ��  	  �F  	  �F  _  ��  _      B  , ,  ��  _  ��  	  ��  	  ��  _  ��  _      B  , ,  �8  _  �8  	  ��  	  ��  _  �8  _      B  , ,  ��  _  ��  	  �0  	  �0  _  ��  _      B  , ,  ��  _  ��  	  �~  	  �~  _  ��  _      B  , ,  �N    �N  �  ��  �  ��    �N        B  , ,  ��    ��  �  �F  �  �F    ��        B  , ,  �  c  �    ��    ��  c  �  c      B  , ,  �d  c  �d    �    �  c  �d  c      B  , ,  ��  c  ��    �\    �\  c  ��  c      B  , ,  �   c  �     ��    ��  c  �   c      B  , ,  �N  c  �N    ��    ��  c  �N  c      B  , ,  ��  c  ��    �F    �F  c  ��  c      B  , ,  ��  c  ��    ��    ��  c  ��  c      B  , ,  �8  c  �8    ��    ��  c  �8  c      B  , ,  ��  c  ��    �0    �0  c  ��  c      B  , ,  ��  c  ��    �~    �~  c  ��  c      B  , ,  ��    ��  �  ��  �  ��    ��        B  , ,  �8    �8  �  ��  �  ��    �8        B  , ,  ��    ��  �  �0  �  �0    ��        B  , ,  ��    ��  �  �~  �  �~    ��        B  , ,  �    �  �  ��  �  ��    �        B  , ,  �d    �d  �  �  �  �    �d        B  , ,  ��    ��  �  �\  �  �\    ��        B  , ,  �  �  �  a  ��  a  ��  �  �  �      B  , ,  �d  �  �d  a  �  a  �  �  �d  �      B  , ,  ��  �  ��  a  �\  a  �\  �  ��  �      B  , ,  �   �  �   a  ��  a  ��  �  �   �      B  , ,  �N  �  �N  a  ��  a  ��  �  �N  �      B  , ,  ����  �����  ������  �����  ����      B  , ,  �d���  �d����  �����  ����  �d���      B  , ,  �����  ������  �\����  �\���  �����      B  , ,  � ���  � ����  ������  �����  � ���      B  , ,  �N���  �N����  ������  �����  �N���      B  , ,  �����  ������  �F����  �F���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �8���  �8����  ������  �����  �8���      B  , ,  �����  ������  �0����  �0���  �����      B  , ,  �����  ������  �~����  �~���  �����      B  , ,  ��  �  ��  a  �F  a  �F  �  ��  �      B  , ,  �     �   �  ��   �  ��     �         B  , ,  �d     �d   �  �   �  �     �d         B  , ,  ��     ��   �  �\   �  �\     ��         B  , ,  �      �    �  ��   �  ��     �          B  , ,  �N     �N   �  ��   �  ��     �N         B  , ,  ��     ��   �  �F   �  �F     ��         B  , ,  ��     ��   �  ��   �  ��     ��         B  , ,  �8     �8   �  ��   �  ��     �8         B  , ,  ��     ��   �  �0   �  �0     ��         B  , ,  ��     ��   �  �~   �  �~     ��         B  , ,  ��  �  ��  a  ��  a  ��  �  ��  �      B  , ,  �8  �  �8  a  ��  a  ��  �  �8  �      B  , ,  ��  �  ��  a  �0  a  �0  �  ��  �      B  , ,  �����  ����e  �����e  ������  �����      B  , ,  �d����  �d���e  ����e  �����  �d����      B  , ,  ������  �����e  �\���e  �\����  ������      B  , ,  ����g  ����  �����  �����g  ����g      B  , ,  �d���g  �d���  ����  ����g  �d���g      B  , ,  �����g  �����  �\���  �\���g  �����g      B  , ,  � ���g  � ���  �����  �����g  � ���g      B  , ,  �N���g  �N���  �����  �����g  �N���g      B  , ,  �����g  �����  �F���  �F���g  �����g      B  , ,  �����g  �����  �����  �����g  �����g      B  , ,  ������  �����I  �H���I  �H����  ������      B  , ,  ������  ������  �H����  �H����  ������      B  , ,  �����/  ������  �H����  �H���/  �����/      B  , ,  �����  ������  �H����  �H���  �����      B  , ,  �����  �����S  �f���S  �f���  �����      B  , ,  �����U  ������  �f����  �f���U  �����U      B  , ,  �����  �����  �f���  �f���  �����      B  , ,  �����  �����W  �f���W  �f���  �����      B  , ,  �����Y  �����  �f���  �f���Y  �����Y      B  , ,  �����  �����  �f���  �f���  �����      B  , ,  �����  �����[  �f���[  �f���  �����      B  , ,  �����]  �����  �f���  �f���]  �����]      B  , ,  �����U  ������  �f����  �f���U  �����U      B  , ,  �����  ����ܫ  �f��ܫ  �f���  �����      B  , ,  ����ڭ  �����W  �f���W  �f��ڭ  ����ڭ      B  , ,  �����Y  �����  �f���  �f���Y  �����Y      B  , ,  �����  ����د  �f��د  �f���  �����      B  , ,  ����ֱ  �����[  �f���[  �f��ֱ  ����ֱ      B  , ,  �����]  �����  �f���  �f���]  �����]      B  , ,  �����	  ����Գ  �f��Գ  �f���	  �����	      B  , ,  ����ϕ  �����?  �H���?  �H��ϕ  ����ϕ      B  , ,  ������  ����·  �H��·  �H����  ������      B  , ,  �����%  ������  �H����  �H���%  �����%      B  , ,  �����  ����ʽ  �H��ʽ  �H���  �����      B  , ,  ����ş  �����I  �f���I  �f��ş  ����ş      B  , ,  �����K  ������  �f����  �f���K  �����K      B  , ,  ������  ����á  �f��á  �f����  ������      B  , ,  ������  �����M  �f���M  �f����  ������      B  , ,  �����O  ������  �f����  �f���O  �����O      B  , ,  �����  �����S  �r���S  �r���  �����      B  , ,  �����U  ������  �r����  �r���U  �����U      B  , ,  �
���  �
���  �����  �����  �
���      B  , ,  �X���  �X���  ����  ����  �X���      B  , ,  �����  �����  �P���  �P���  �����      B  , ,  �����  �����  �����  �����  �����      B  , ,  �B���  �B���  �����  �����  �B���      B  , ,  �����  �����  �:���  �:���  �����      B  , ,  �����  �����  �����  �����  �����      B  , ,  �,���  �,���  �����  �����  �,���      B  , ,  �z���  �z���  �$���  �$���  �z���      B  , ,  �����  �����  �r���  �r���  �����      B  , ,  ����  ����  �����  �����  ����      B  , ,  �d���  �d���  ����  ����  �d���      B  , ,  �����  �����  �\���  �\���  �����      B  , ,  � ���  � ���  �����  �����  � ���      B  , ,  �N���  �N���  �����  �����  �N���      B  , ,  �����  �����  �F���  �F���  �����      B  , ,  �����  �����  �����  �����  �����      B  , ,  �8���  �8���  �����  �����  �8���      B  , ,  �����  �����  �0���  �0���  �����      B  , ,  �����  �����  �~���  �~���  �����      B  , ,  �����  �����W  �r���W  �r���  �����      B  , ,  �����Y  �����  �r���  �r���Y  �����Y      B  , ,  �����  �����  �r���  �r���  �����      B  , ,  �����  �����[  �r���[  �r���  �����      B  , ,  �����]  �����  �r���  �r���]  �����]      B  , ,  �����U  ������  �r����  �r���U  �����U      B  , ,  �*���/  �*����  ������  �����/  �*���/      B  , ,  �~���/  �~����  �(����  �(���/  �~���/      B  , ,  �����/  ������  �|����  �|���/  �����/      B  , ,  �&���/  �&����  ������  �����/  �&���/      B  , ,  �z���/  �z����  �$����  �$���/  �z���/      B  , ,  �����/  ������  �x����  �x���/  �����/      B  , ,  �"���/  �"����  ������  �����/  �"���/      B  , ,  �v���/  �v����  � ����  � ���/  �v���/      B  , ,  �����/  ������  �t����  �t���/  �����/      B  , ,  ����/  �����  ������  �����/  ����/      B  , ,  �r���/  �r����  �����  ����/  �r���/      B  , ,  �����/  ������  �p����  �p���/  �����/      B  , ,  �����  ������  �0����  �0���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �.���  �.����  ������  �����  �.���      B  , ,  �����  ������  �,����  �,���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �*���  �*����  ������  �����  �*���      B  , ,  �~���  �~����  �(����  �(���  �~���      B  , ,  �����  ������  �|����  �|���  �����      B  , ,  �&���  �&����  ������  �����  �&���      B  , ,  �z���  �z����  �$����  �$���  �z���      B  , ,  �����  ������  �x����  �x���  �����      B  , ,  �"���  �"����  ������  �����  �"���      B  , ,  �v���  �v����  � ����  � ���  �v���      B  , ,  �����  ������  �t����  �t���  �����      B  , ,  ����  �����  ������  �����  ����      B  , ,  �r���  �r����  �����  ����  �r���      B  , ,  �����  ������  �p����  �p���  �����      B  , ,  �"����  �"���I  �����I  ������  �"����      B  , ,  ����  ����S  �����S  �����  ����      B  , ,  �d���  �d���S  ����S  ����  �d���      B  , ,  �����  �����S  �\���S  �\���  �����      B  , ,  � ���  � ���S  �����S  �����  � ���      B  , ,  �N���  �N���S  �����S  �����  �N���      B  , ,  �����  �����S  �F���S  �F���  �����      B  , ,  �����  �����S  �����S  �����  �����      B  , ,  �8���  �8���S  �����S  �����  �8���      B  , ,  �����  �����S  �0���S  �0���  �����      B  , ,  �����  �����S  �~���S  �~���  �����      B  , ,  �v����  �v���I  � ���I  � ����  �v����      B  , ,  ����U  �����  ������  �����U  ����U      B  , ,  �d���U  �d����  �����  ����U  �d���U      B  , ,  �����U  ������  �\����  �\���U  �����U      B  , ,  � ���U  � ����  ������  �����U  � ���U      B  , ,  �N���U  �N����  ������  �����U  �N���U      B  , ,  �����U  ������  �F����  �F���U  �����U      B  , ,  �����U  ������  ������  �����U  �����U      B  , ,  �8���U  �8����  ������  �����U  �8���U      B  , ,  �����U  ������  �0����  �0���U  �����U      B  , ,  �����U  ������  �~����  �~���U  �����U      B  , ,  ������  �����I  �t���I  �t����  ������      B  , ,  �����  ����I  �����I  ������  �����      B  , ,  �r����  �r���I  ����I  �����  �r����      B  , ,  ������  �����I  �p���I  �p����  ������      B  , ,  ������  ������  �0����  �0����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �.����  �.����  ������  ������  �.����      B  , ,  ������  ������  �,����  �,����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �*����  �*����  ������  ������  �*����      B  , ,  �~����  �~����  �(����  �(����  �~����      B  , ,  ������  ������  �|����  �|����  ������      B  , ,  �&����  �&����  ������  ������  �&����      B  , ,  �z����  �z����  �$����  �$����  �z����      B  , ,  ������  ������  �x����  �x����  ������      B  , ,  �"����  �"����  ������  ������  �"����      B  , ,  �v����  �v����  � ����  � ����  �v����      B  , ,  ������  ������  �t����  �t����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �r����  �r����  �����  �����  �r����      B  , ,  ������  ������  �p����  �p����  ������      B  , ,  �����/  ������  �0����  �0���/  �����/      B  , ,  �����/  ������  ������  �����/  �����/      B  , ,  �.���/  �.����  ������  �����/  �.���/      B  , ,  �����/  ������  �,����  �,���/  �����/      B  , ,  �����/  ������  ������  �����/  �����/      B  , ,  ������  �����I  �0���I  �0����  ������      B  , ,  ������  �����I  �����I  ������  ������      B  , ,  �.����  �.���I  �����I  ������  �.����      B  , ,  ������  �����I  �,���I  �,����  ������      B  , ,  ������  �����I  �����I  ������  ������      B  , ,  �*����  �*���I  �����I  ������  �*����      B  , ,  �~����  �~���I  �(���I  �(����  �~����      B  , ,  ������  �����I  �|���I  �|����  ������      B  , ,  �&����  �&���I  �����I  ������  �&����      B  , ,  �z����  �z���I  �$���I  �$����  �z����      B  , ,  ������  �����I  �x���I  �x����  ������      B  , ,  �B���  �B���S  �����S  �����  �B���      B  , ,  �����  �����S  �:���S  �:���  �����      B  , ,  �����  �����S  �����S  �����  �����      B  , ,  �,���  �,���S  �����S  �����  �,���      B  , ,  �z���  �z���S  �$���S  �$���  �z���      B  , ,  �����/  ������  ������  �����/  �����/      B  , ,  �2���/  �2����  ������  �����/  �2���/      B  , ,  �2����  �2����  ������  ������  �2����      B  , ,  ������  �����I  �����I  ������  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �F����  �F����  ������  ������  �F����      B  , ,  ������  ������  �D����  �D����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �B����  �B����  ������  ������  �B����      B  , ,  ������  ������  �@����  �@����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �B����  �B���I  �����I  ������  �B����      B  , ,  �
���U  �
����  ������  �����U  �
���U      B  , ,  �X���U  �X����  �����  ����U  �X���U      B  , ,  �����U  ������  �P����  �P���U  �����U      B  , ,  �����U  ������  ������  �����U  �����U      B  , ,  �B���U  �B����  ������  �����U  �B���U      B  , ,  �����U  ������  �:����  �:���U  �����U      B  , ,  �����U  ������  ������  �����U  �����U      B  , ,  �,���U  �,����  ������  �����U  �,���U      B  , ,  �z���U  �z����  �$����  �$���U  �z���U      B  , ,  �>����  �>����  ������  ������  �>����      B  , ,  ������  ������  �<����  �<����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �:����  �:����  ������  ������  �:����      B  , ,  ������  ������  �8����  �8����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �6����  �6����  ������  ������  �6����      B  , ,  ������  ������  �4����  �4����  ������      B  , ,  ������  �����I  �D���I  �D����  ������      B  , ,  �����  ������  ������  �����  �����      B  , ,  �F���  �F����  ������  �����  �F���      B  , ,  ������  �����I  �@���I  �@����  ������      B  , ,  �����  ������  �D����  �D���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �B���  �B����  ������  �����  �B���      B  , ,  �����  ������  �@����  �@���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �>���  �>����  ������  �����  �>���      B  , ,  �����  ������  �<����  �<���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �:���  �:����  ������  �����  �:���      B  , ,  �����  ������  �8����  �8���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �6���  �6����  ������  �����  �6���      B  , ,  �����  ������  �4����  �4���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �2���  �2����  ������  �����  �2���      B  , ,  ������  ������  ������  ������  ������      B  , ,  �F����  �F���I  �����I  ������  �F����      B  , ,  �����/  ������  ������  �����/  �����/      B  , ,  �F���/  �F����  ������  �����/  �F���/      B  , ,  �����/  ������  �D����  �D���/  �����/      B  , ,  ������  �����I  �����I  ������  ������      B  , ,  �����/  ������  ������  �����/  �����/      B  , ,  �>����  �>���I  �����I  ������  �>����      B  , ,  �B���/  �B����  ������  �����/  �B���/      B  , ,  ������  �����I  �<���I  �<����  ������      B  , ,  �����/  ������  �@����  �@���/  �����/      B  , ,  ������  �����I  �����I  ������  ������      B  , ,  �����/  ������  ������  �����/  �����/      B  , ,  �:����  �:���I  �����I  ������  �:����      B  , ,  �>���/  �>����  ������  �����/  �>���/      B  , ,  ������  �����I  �8���I  �8����  ������      B  , ,  �����/  ������  �<����  �<���/  �����/      B  , ,  ������  �����I  �����I  ������  ������      B  , ,  �6����  �6���I  �����I  ������  �6����      B  , ,  ������  �����I  �4���I  �4����  ������      B  , ,  ������  �����I  �����I  ������  ������      B  , ,  �2����  �2���I  �����I  ������  �2����      B  , ,  �����/  ������  ������  �����/  �����/      B  , ,  �:���/  �:����  ������  �����/  �:���/      B  , ,  �����/  ������  �8����  �8���/  �����/      B  , ,  �����/  ������  ������  �����/  �����/      B  , ,  �6���/  �6����  ������  �����/  �6���/      B  , ,  �����/  ������  �4����  �4���/  �����/      B  , ,  ������  �����I  �����I  ������  ������      B  , ,  �
���  �
���S  �����S  �����  �
���      B  , ,  �X���  �X���S  ����S  ����  �X���      B  , ,  �����  �����S  �P���S  �P���  �����      B  , ,  �����  �����S  �����S  �����  �����      B  , ,  �����  �����  �:���  �:���  �����      B  , ,  �����  �����  �����  �����  �����      B  , ,  �,���  �,���  �����  �����  �,���      B  , ,  �z���  �z���  �$���  �$���  �z���      B  , ,  �B���  �B���W  �����W  �����  �B���      B  , ,  �����  �����W  �:���W  �:���  �����      B  , ,  �
���  �
���[  �����[  �����  �
���      B  , ,  �X���  �X���[  ����[  ����  �X���      B  , ,  �����  �����[  �P���[  �P���  �����      B  , ,  �����  �����[  �����[  �����  �����      B  , ,  �B���  �B���[  �����[  �����  �B���      B  , ,  �����  �����[  �:���[  �:���  �����      B  , ,  �����  �����[  �����[  �����  �����      B  , ,  �,���  �,���[  �����[  �����  �,���      B  , ,  �z���  �z���[  �$���[  �$���  �z���      B  , ,  �����  �����W  �����W  �����  �����      B  , ,  �,���  �,���W  �����W  �����  �,���      B  , ,  �
���]  �
���  �����  �����]  �
���]      B  , ,  �X���]  �X���  ����  ����]  �X���]      B  , ,  �����]  �����  �P���  �P���]  �����]      B  , ,  �����]  �����  �����  �����]  �����]      B  , ,  �B���]  �B���  �����  �����]  �B���]      B  , ,  �����]  �����  �:���  �:���]  �����]      B  , ,  �����]  �����  �����  �����]  �����]      B  , ,  �,���]  �,���  �����  �����]  �,���]      B  , ,  �z���]  �z���  �$���  �$���]  �z���]      B  , ,  �z���  �z���W  �$���W  �$���  �z���      B  , ,  ������  �����  �����  ������  ������      B  , ,  �1����  �1���  �����  ������  �1����      B  , ,  �����  ����  �)���  �)����  �����      B  , ,  ������  �����  �w���  �w����  ������      B  , ,  �����  ����  �����  ������  �����      B  , ,  �i����  �i���  ����  �����  �i����      B  , ,  ������  �����  �a���  �a����  ������      B  , ,  �����  ����  �����  ������  �����      B  , ,  �S����  �S���  �����  ������  �S����      B  , ,  ������  �����  �K���  �K����  ������      B  , ,  ������  �����u  �����u  ������  ������      B  , ,  �1����  �1���u  �����u  ������  �1����      B  , ,  �����  ����u  �)���u  �)����  �����      B  , ,  ������  �����u  �w���u  �w����  ������      B  , ,  �����  ����u  �����u  ������  �����      B  , ,  �i����  �i���u  ����u  �����  �i����      B  , ,  ������  �����u  �a���u  �a����  ������      B  , ,  �����  ����u  �����u  ������  �����      B  , ,  �S����  �S���u  �����u  ������  �S����      B  , ,  ������  �����u  �K���u  �K����  ������      B  , ,  �
���  �
���W  �����W  �����  �
���      B  , ,  �
���U  �
����  ������  �����U  �
���U      B  , ,  �X���U  �X����  �����  ����U  �X���U      B  , ,  �����U  ������  �P����  �P���U  �����U      B  , ,  �����U  ������  ������  �����U  �����U      B  , ,  �B���U  �B����  ������  �����U  �B���U      B  , ,  �����U  ������  �:����  �:���U  �����U      B  , ,  �����U  ������  ������  �����U  �����U      B  , ,  �,���U  �,����  ������  �����U  �,���U      B  , ,  �z���U  �z����  �$����  �$���U  �z���U      B  , ,  �X���  �X���W  ����W  ����  �X���      B  , ,  �
���Y  �
���  �����  �����Y  �
���Y      B  , ,  �X���Y  �X���  ����  ����Y  �X���Y      B  , ,  �����Y  �����  �P���  �P���Y  �����Y      B  , ,  �����Y  �����  �����  �����Y  �����Y      B  , ,  �B���Y  �B���  �����  �����Y  �B���Y      B  , ,  �����Y  �����  �:���  �:���Y  �����Y      B  , ,  �����Y  �����  �����  �����Y  �����Y      B  , ,  �,���Y  �,���  �����  �����Y  �,���Y      B  , ,  �z���Y  �z���  �$���  �$���Y  �z���Y      B  , ,  �����  �����W  �P���W  �P���  �����      B  , ,  �����  �����W  �����W  �����  �����      B  , ,  �
���  �
���  �����  �����  �
���      B  , ,  �X���  �X���  ����  ����  �X���      B  , ,  �����  �����  �P���  �P���  �����      B  , ,  �����  �����  �����  �����  �����      B  , ,  �B���  �B���  �����  �����  �B���      B  , ,  �8���]  �8���  �����  �����]  �8���]      B  , ,  �����]  �����  �0���  �0���]  �����]      B  , ,  �����]  �����  �~���  �~���]  �����]      B  , ,  �����  �����  �\���  �\���  �����      B  , ,  � ���  � ���  �����  �����  � ���      B  , ,  �N���  �N���  �����  �����  �N���      B  , ,  �����  �����  �F���  �F���  �����      B  , ,  �����  �����  �����  �����  �����      B  , ,  �8���  �8���  �����  �����  �8���      B  , ,  �����  �����  �0���  �0���  �����      B  , ,  �����  �����  �~���  �~���  �����      B  , ,  �d���Y  �d���  ����  ����Y  �d���Y      B  , ,  �����Y  �����  �\���  �\���Y  �����Y      B  , ,  ������  �����  �����  ������  ������      B  , ,  �=����  �=���  �����  ������  �=����      B  , ,  ������  �����  �5���  �5����  ������      B  , ,  ������  �����  �����  ������  ������      B  , ,  �'����  �'���  �����  ������  �'����      B  , ,  �u����  �u���  ����  �����  �u����      B  , ,  ������  �����  �m���  �m����  ������      B  , ,  �����  ����  �����  ������  �����      B  , ,  �_����  �_���  �	���  �	����  �_����      B  , ,  ������  �����  �W���  �W����  ������      B  , ,  � ���Y  � ���  �����  �����Y  � ���Y      B  , ,  �N���Y  �N���  �����  �����Y  �N���Y      B  , ,  �����Y  �����  �F���  �F���Y  �����Y      B  , ,  �����Y  �����  �����  �����Y  �����Y      B  , ,  �8���Y  �8���  �����  �����Y  �8���Y      B  , ,  �����Y  �����  �0���  �0���Y  �����Y      B  , ,  �����Y  �����  �~���  �~���Y  �����Y      B  , ,  �d���  �d���W  ����W  ����  �d���      B  , ,  �����  �����W  �\���W  �\���  �����      B  , ,  ����  ����[  �����[  �����  ����      B  , ,  ������  �����u  �����u  ������  ������      B  , ,  �=����  �=���u  �����u  ������  �=����      B  , ,  ������  �����u  �5���u  �5����  ������      B  , ,  ������  �����u  �����u  ������  ������      B  , ,  �'����  �'���u  �����u  ������  �'����      B  , ,  �u����  �u���u  ����u  �����  �u����      B  , ,  ������  �����u  �m���u  �m����  ������      B  , ,  �����  ����u  �����u  ������  �����      B  , ,  �_����  �_���u  �	���u  �	����  �_����      B  , ,  ������  �����u  �W���u  �W����  ������      B  , ,  �d���  �d���[  ����[  ����  �d���      B  , ,  �����  �����[  �\���[  �\���  �����      B  , ,  � ���  � ���[  �����[  �����  � ���      B  , ,  �N���  �N���[  �����[  �����  �N���      B  , ,  �����  �����[  �F���[  �F���  �����      B  , ,  �����  �����[  �����[  �����  �����      B  , ,  �8���  �8���[  �����[  �����  �8���      B  , ,  �����  �����[  �0���[  �0���  �����      B  , ,  �����  �����[  �~���[  �~���  �����      B  , ,  � ���  � ���W  �����W  �����  � ���      B  , ,  �N���  �N���W  �����W  �����  �N���      B  , ,  ����U  �����  ������  �����U  ����U      B  , ,  �d���U  �d����  �����  ����U  �d���U      B  , ,  �����U  ������  �\����  �\���U  �����U      B  , ,  � ���U  � ����  ������  �����U  � ���U      B  , ,  �N���U  �N����  ������  �����U  �N���U      B  , ,  �����U  ������  �F����  �F���U  �����U      B  , ,  �����U  ������  ������  �����U  �����U      B  , ,  �8���U  �8����  ������  �����U  �8���U      B  , ,  �����U  ������  �0����  �0���U  �����U      B  , ,  �����U  ������  �~����  �~���U  �����U      B  , ,  �����  �����W  �F���W  �F���  �����      B  , ,  �����  �����W  �����W  �����  �����      B  , ,  �8���  �8���W  �����W  �����  �8���      B  , ,  �����  �����W  �0���W  �0���  �����      B  , ,  �����  �����W  �~���W  �~���  �����      B  , ,  ����  ����W  �����W  �����  ����      B  , ,  ����Y  ����  �����  �����Y  ����Y      B  , ,  ����  ����  �����  �����  ����      B  , ,  �d���  �d���  ����  ����  �d���      B  , ,  ����]  ����  �����  �����]  ����]      B  , ,  �d���]  �d���  ����  ����]  �d���]      B  , ,  �����]  �����  �\���  �\���]  �����]      B  , ,  � ���]  � ���  �����  �����]  � ���]      B  , ,  �N���]  �N���  �����  �����]  �N���]      B  , ,  �����]  �����  �F���  �F���]  �����]      B  , ,  �����]  �����  �����  �����]  �����]      B  , ,  r����  r����W  sZ���W  sZ���  r����      B  , ,  r����Y  r����  sZ���  sZ���Y  r����Y      B  , ,  r����  r����  sZ���  sZ���  r����      B  , ,  r����  r����[  sZ���[  sZ���  r����      B  , ,  r����  r����S  sZ���S  sZ���  r����      B  , ,  r����]  r����  sZ���  sZ���]  r����]      B  , ,  r����U  r�����  sZ����  sZ���U  r����U      B  , ,  r����U  r�����  sZ����  sZ���U  r����U      B  , ,  [�����  [����y  \b���y  \b����  [�����      B  , ,  ]����  ]����  ^����  ^����  ]����      B  , ,  `@���  `@���  `����  `����  `@���      B  , ,  b����  b����  c8���  c8���  b����      B  , ,  d����  d����  e����  e����  d����      B  , ,  g*���  g*���  g����  g����  g*���      B  , ,  ix���  ix���  j"���  j"���  ix���      B  , ,  k����  k����  lp���  lp���  k����      B  , ,  n���  n���  n����  n����  n���      B  , ,  pb���  pb���  q���  q���  pb���      B  , ,  r����  r����  sZ���  sZ���  r����      B  , ,  t����  t����  u����  u����  t����      B  , ,  wL���  wL���  w����  w����  wL���      B  , ,  y����  y����  zD���  zD���  y����      B  , ,  {����  {����  |����  |����  {����      B  , ,  ~6���  ~6���  ~����  ~����  ~6���      B  , ,  �����  �����  �.���  �.���  �����      B  , ,  �����  �����  �|���  �|���  �����      B  , ,  � ���  � ���  �����  �����  � ���      B  , ,  �n���  �n���  ����  ����  �n���      B  , ,  t^����  t^���I  u���I  u����  t^����      B  , ,  �R����  �R���I  �����I  ������  �R����      B  , ,  s
���  s
����  s�����  s����  s
���      B  , ,  t����  t����S  u����S  u����  t����      B  , ,  wL���  wL���S  w����S  w����  wL���      B  , ,  y����  y����S  zD���S  zD���  y����      B  , ,  {����  {����S  |����S  |����  {����      B  , ,  ~6���  ~6���S  ~����S  ~����  ~6���      B  , ,  �����  �����S  �.���S  �.���  �����      B  , ,  t^���  t^����  u����  u���  t^���      B  , ,  �����  �����S  �|���S  �|���  �����      B  , ,  � ���  � ���S  �����S  �����  � ���      B  , ,  �n���  �n���S  ����S  ����  �n���      B  , ,  s
���/  s
����  s�����  s����/  s
���/      B  , ,  t^���/  t^����  u����  u���/  t^���/      B  , ,  u����/  u�����  v\����  v\���/  u����/      B  , ,  w���/  w����  w�����  w����/  w���/      B  , ,  xZ���/  xZ����  y����  y���/  xZ���/      B  , ,  y����/  y�����  zX����  zX���/  y����/      B  , ,  {���/  {����  {�����  {����/  {���/      B  , ,  |V���/  |V����  } ����  } ���/  |V���/      B  , ,  }����/  }�����  ~T����  ~T���/  }����/      B  , ,  ~����/  ~�����  �����  ����/  ~����/      B  , ,  �R���/  �R����  ������  �����/  �R���/      B  , ,  �����/  ������  �P����  �P���/  �����/      B  , ,  �����/  ������  ������  �����/  �����/      B  , ,  �N���/  �N����  ������  �����/  �N���/      B  , ,  �����/  ������  �L����  �L���/  �����/      B  , ,  u����  u�����  v\����  v\���  u����      B  , ,  t����U  t�����  u�����  u����U  t����U      B  , ,  wL���U  wL����  w�����  w����U  wL���U      B  , ,  y����U  y�����  zD����  zD���U  y����U      B  , ,  {����U  {�����  |�����  |����U  {����U      B  , ,  ~6���U  ~6����  ~�����  ~����U  ~6���U      B  , ,  �����U  ������  �.����  �.���U  �����U      B  , ,  �����U  ������  �|����  �|���U  �����U      B  , ,  � ���U  � ����  ������  �����U  � ���U      B  , ,  �n���U  �n����  �����  ����U  �n���U      B  , ,  �����/  ������  ������  �����/  �����/      B  , ,  �J���/  �J����  ������  �����/  �J���/      B  , ,  s
����  s
����  s�����  s�����  s
����      B  , ,  t^����  t^����  u����  u����  t^����      B  , ,  u�����  u�����  v\����  v\����  u�����      B  , ,  w����  w����  w�����  w�����  w����      B  , ,  xZ����  xZ����  y����  y����  xZ����      B  , ,  y�����  y�����  zX����  zX����  y�����      B  , ,  {����  {����  {�����  {�����  {����      B  , ,  |V����  |V����  } ����  } ����  |V����      B  , ,  w���  w����  w�����  w����  w���      B  , ,  }�����  }�����  ~T����  ~T����  }�����      B  , ,  ~�����  ~�����  �����  �����  ~�����      B  , ,  �R����  �R����  ������  ������  �R����      B  , ,  ������  ������  �P����  �P����  ������      B  , ,  xZ���  xZ����  y����  y���  xZ���      B  , ,  y����  y�����  zX����  zX���  y����      B  , ,  {���  {����  {�����  {����  {���      B  , ,  |V���  |V����  } ����  } ���  |V���      B  , ,  }����  }�����  ~T����  ~T���  }����      B  , ,  ������  �����I  �P���I  �P����  ������      B  , ,  ~����  ~�����  �����  ����  ~����      B  , ,  �R���  �R����  ������  �����  �R���      B  , ,  �����  ������  �P����  �P���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �N���  �N����  ������  �����  �N���      B  , ,  �����  ������  �L����  �L���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �J���  �J����  ������  �����  �J���      B  , ,  �N����  �N���I  �����I  ������  �N����      B  , ,  ������  �����I  �L���I  �L����  ������      B  , ,  ������  �����I  �����I  ������  ������      B  , ,  �J����  �J���I  �����I  ������  �J����      B  , ,  s
����  s
���I  s����I  s�����  s
����      B  , ,  ������  �����I  �����I  ������  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �N����  �N����  ������  ������  �N����      B  , ,  ������  ������  �L����  �L����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �J����  �J����  ������  ������  �J����      B  , ,  u�����  u����I  v\���I  v\����  u�����      B  , ,  w����  w���I  w����I  w�����  w����      B  , ,  xZ����  xZ���I  y���I  y����  xZ����      B  , ,  y�����  y����I  zX���I  zX����  y�����      B  , ,  {����  {���I  {����I  {�����  {����      B  , ,  |V����  |V���I  } ���I  } ����  |V����      B  , ,  }�����  }����I  ~T���I  ~T����  }�����      B  , ,  ~�����  ~����I  ����I  �����  ~�����      B  , ,  pb����  pb���I  q���I  q����  pb����      B  , ,  q�����  q����I  r`���I  r`����  q�����      B  , ,  c���  c����  c�����  c����  c���      B  , ,  dn���  dn����  e����  e���  dn���      B  , ,  e����  e�����  fl����  fl���  e����      B  , ,  ]�����  ]����I  ^t���I  ^t����  ]�����      B  , ,  ]�����  ]�����  ^t����  ^t����  ]�����      B  , ,  [����#  [�����  \b����  \b���#  [����#      B  , ,  ]����U  ]�����  ^�����  ^����U  ]����U      B  , ,  `@���U  `@����  `�����  `����U  `@���U      B  , ,  b����U  b�����  c8����  c8���U  b����U      B  , ,  d����U  d�����  e�����  e����U  d����U      B  , ,  g*���U  g*����  g�����  g����U  g*���U      B  , ,  ix���U  ix����  j"����  j"���U  ix���U      B  , ,  k����U  k�����  lp����  lp���U  k����U      B  , ,  n���U  n����  n�����  n����U  n���U      B  , ,  pb���U  pb����  q����  q���U  pb���U      B  , ,  _����  _����  _�����  _�����  _����      B  , ,  `r����  `r����  a����  a����  `r����      B  , ,  a�����  a�����  bp����  bp����  a�����      B  , ,  c����  c����  c�����  c�����  c����      B  , ,  dn����  dn����  e����  e����  dn����      B  , ,  e�����  e�����  fl����  fl����  e�����      B  , ,  g����  g����  g�����  g�����  g����      B  , ,  hj����  hj����  i����  i����  hj����      B  , ,  _����  _���I  _����I  _�����  _����      B  , ,  ]����/  ]�����  ^t����  ^t���/  ]����/      B  , ,  _���/  _����  _�����  _����/  _���/      B  , ,  `r���/  `r����  a����  a���/  `r���/      B  , ,  i�����  i�����  jh����  jh����  i�����      B  , ,  k����  k����  k�����  k�����  k����      B  , ,  lf����  lf����  m����  m����  lf����      B  , ,  m�����  m�����  nd����  nd����  m�����      B  , ,  o����  o����  o�����  o�����  o����      B  , ,  pb����  pb����  q����  q����  pb����      B  , ,  q�����  q�����  r`����  r`����  q�����      B  , ,  a����/  a�����  bp����  bp���/  a����/      B  , ,  c���/  c����  c�����  c����/  c���/      B  , ,  dn���/  dn����  e����  e���/  dn���/      B  , ,  e����/  e�����  fl����  fl���/  e����/      B  , ,  g���/  g����  g�����  g����/  g���/      B  , ,  hj���/  hj����  i����  i���/  hj���/      B  , ,  g���  g����  g�����  g����  g���      B  , ,  i����/  i�����  jh����  jh���/  i����/      B  , ,  a�����  a����I  bp���I  bp����  a�����      B  , ,  [����  [�����  \b����  \b���  [����      B  , ,  [�����  [����u  \b���u  \b����  [�����      B  , ,  [����w  [����!  \b���!  \b���w  [����w      B  , ,  ]����  ]����S  ^����S  ^����  ]����      B  , ,  `@���  `@���S  `����S  `����  `@���      B  , ,  b����  b����S  c8���S  c8���  b����      B  , ,  d����  d����S  e����S  e����  d����      B  , ,  g*���  g*���S  g����S  g����  g*���      B  , ,  ix���  ix���S  j"���S  j"���  ix���      B  , ,  k����  k����S  lp���S  lp���  k����      B  , ,  n���  n���S  n����S  n����  n���      B  , ,  pb���  pb���S  q���S  q���  pb���      B  , ,  hj���  hj����  i����  i���  hj���      B  , ,  i����  i�����  jh����  jh���  i����      B  , ,  k���  k����  k�����  k����  k���      B  , ,  lf���  lf����  m����  m���  lf���      B  , ,  m����  m�����  nd����  nd���  m����      B  , ,  o���  o����  o�����  o����  o���      B  , ,  pb���  pb����  q����  q���  pb���      B  , ,  q����  q�����  r`����  r`���  q����      B  , ,  ]����  ]�����  ^t����  ^t���  ]����      B  , ,  _���  _����  _�����  _����  _���      B  , ,  `r���  `r����  a����  a���  `r���      B  , ,  k���/  k����  k�����  k����/  k���/      B  , ,  lf���/  lf����  m����  m���/  lf���/      B  , ,  m����/  m�����  nd����  nd���/  m����/      B  , ,  o���/  o����  o�����  o����/  o���/      B  , ,  pb���/  pb����  q����  q���/  pb���/      B  , ,  q����/  q�����  r`����  r`���/  q����/      B  , ,  c����  c���I  c����I  c�����  c����      B  , ,  a����  a�����  bp����  bp���  a����      B  , ,  dn����  dn���I  e���I  e����  dn����      B  , ,  `r����  `r���I  a���I  a����  `r����      B  , ,  e�����  e����I  fl���I  fl����  e�����      B  , ,  hj����  hj���I  i���I  i����  hj����      B  , ,  g����  g���I  g����I  g�����  g����      B  , ,  i�����  i����I  jh���I  jh����  i�����      B  , ,  k����  k���I  k����I  k�����  k����      B  , ,  lf����  lf���I  m���I  m����  lf����      B  , ,  m�����  m����I  nd���I  nd����  m�����      B  , ,  o����  o���I  o����I  o�����  o����      B  , ,  _����  _���u  _����u  _�����  _����      B  , ,  ag����  ag���u  b���u  b����  ag����      B  , ,  c�����  c����u  d_���u  d_����  c�����      B  , ,  f����  f���u  f����u  f�����  f����      B  , ,  hQ����  hQ���u  h����u  h�����  hQ����      B  , ,  j�����  j����u  kI���u  kI����  j�����      B  , ,  l�����  l����u  m����u  m�����  l�����      B  , ,  o;����  o;���u  o����u  o�����  o;����      B  , ,  q�����  q����u  r3���u  r3����  q�����      B  , ,  `@���]  `@���  `����  `����]  `@���]      B  , ,  b����]  b����  c8���  c8���]  b����]      B  , ,  d����]  d����  e����  e����]  d����]      B  , ,  g*���]  g*���  g����  g����]  g*���]      B  , ,  ix���]  ix���  j"���  j"���]  ix���]      B  , ,  k����]  k����  lp���  lp���]  k����]      B  , ,  n���]  n���  n����  n����]  n���]      B  , ,  pb���]  pb���  q���  q���]  pb���]      B  , ,  ix���Y  ix���  j"���  j"���Y  ix���Y      B  , ,  k����Y  k����  lp���  lp���Y  k����Y      B  , ,  n���Y  n���  n����  n����Y  n���Y      B  , ,  pb���Y  pb���  q���  q���Y  pb���Y      B  , ,  `@���  `@���W  `����W  `����  `@���      B  , ,  b����  b����W  c8���W  c8���  b����      B  , ,  [�����  [����}  \b���}  \b����  [�����      B  , ,  ]����  ]����  ^����  ^����  ]����      B  , ,  [����  [����)  \b���)  \b���  [����      B  , ,  ]����  ]����[  ^����[  ^����  ]����      B  , ,  `@���  `@���[  `����[  `����  `@���      B  , ,  b����  b����[  c8���[  c8���  b����      B  , ,  [�����  [���߅  \b��߅  \b����  [�����      B  , ,  [���݇  [����1  \b���1  \b��݇  [���݇      B  , ,  ]����U  ]�����  ^�����  ^����U  ]����U      B  , ,  `@���U  `@����  `�����  `����U  `@���U      B  , ,  b����U  b�����  c8����  c8���U  b����U      B  , ,  d����U  d�����  e�����  e����U  d����U      B  , ,  g*���U  g*����  g�����  g����U  g*���U      B  , ,  ix���U  ix����  j"����  j"���U  ix���U      B  , ,  k����U  k�����  lp����  lp���U  k����U      B  , ,  n���U  n����  n�����  n����U  n���U      B  , ,  pb���U  pb����  q����  q���U  pb���U      B  , ,  d����  d����[  e����[  e����  d����      B  , ,  g*���  g*���[  g����[  g����  g*���      B  , ,  ix���  ix���[  j"���[  j"���  ix���      B  , ,  k����  k����[  lp���[  lp���  k����      B  , ,  n���  n���[  n����[  n����  n���      B  , ,  pb���  pb���[  q���[  q���  pb���      B  , ,  `@���  `@���  `����  `����  `@���      B  , ,  b����  b����  c8���  c8���  b����      B  , ,  d����  d����  e����  e����  d����      B  , ,  g*���  g*���  g����  g����  g*���      B  , ,  [�����  [����  \b���  \b����  [�����      B  , ,  [����  [����-  \b���-  \b���  [����      B  , ,  _����  _���  _����  _�����  _����      B  , ,  ag����  ag���  b���  b����  ag����      B  , ,  c�����  c����  d_���  d_����  c�����      B  , ,  f����  f���  f����  f�����  f����      B  , ,  hQ����  hQ���  h����  h�����  hQ����      B  , ,  j�����  j����  kI���  kI����  j�����      B  , ,  l�����  l����  m����  m�����  l�����      B  , ,  o;����  o;���  o����  o�����  o;����      B  , ,  q�����  q����  r3���  r3����  q�����      B  , ,  ix���  ix���  j"���  j"���  ix���      B  , ,  k����  k����  lp���  lp���  k����      B  , ,  n���  n���  n����  n����  n���      B  , ,  pb���  pb���  q���  q���  pb���      B  , ,  d����  d����W  e����W  e����  d����      B  , ,  g*���  g*���W  g����W  g����  g*���      B  , ,  ix���  ix���W  j"���W  j"���  ix���      B  , ,  k����  k����W  lp���W  lp���  k����      B  , ,  n���  n���W  n����W  n����  n���      B  , ,  pb���  pb���W  q���W  q���  pb���      B  , ,  [����{  [����%  \b���%  \b���{  [����{      B  , ,  ]����  ]����W  ^����W  ^����  ]����      B  , ,  [����'  [�����  \b����  \b���'  [����'      B  , ,  ]����Y  ]����  ^����  ^����Y  ]����Y      B  , ,  `@���Y  `@���  `����  `����Y  `@���Y      B  , ,  b����Y  b����  c8���  c8���Y  b����Y      B  , ,  d����Y  d����  e����  e����Y  d����Y      B  , ,  g*���Y  g*���  g����  g����Y  g*���Y      B  , ,  [����+  [�����  \b����  \b���+  [����+      B  , ,  ]����]  ]����  ^����  ^����]  ]����]      B  , ,  [����/  [�����  \b����  \b���/  [����/      B  , ,  �n���  �n���  ����  ����  �n���      B  , ,  �����Y  �����  �.���  �.���Y  �����Y      B  , ,  �����Y  �����  �|���  �|���Y  �����Y      B  , ,  � ���Y  � ���  �����  �����Y  � ���Y      B  , ,  �n���Y  �n���  ����  ����Y  �n���Y      B  , ,  �����  �����W  �.���W  �.���  �����      B  , ,  t����  t����[  u����[  u����  t����      B  , ,  s�����  s����  t����  t�����  s�����      B  , ,  v%����  v%���  v����  v�����  v%����      B  , ,  xs����  xs���  y���  y����  xs����      B  , ,  z�����  z����  {k���  {k����  z�����      B  , ,  }����  }���  }����  }�����  }����      B  , ,  ]����  ]���  ����  �����  ]����      B  , ,  ������  �����  �U���  �U����  ������      B  , ,  ������  �����  �����  ������  ������      B  , ,  �G����  �G���  �����  ������  �G����      B  , ,  ������  �����  �?���  �?����  ������      B  , ,  wL���  wL���[  w����[  w����  wL���      B  , ,  y����  y����[  zD���[  zD���  y����      B  , ,  {����  {����[  |����[  |����  {����      B  , ,  ~6���  ~6���[  ~����[  ~����  ~6���      B  , ,  t����]  t����  u����  u����]  t����]      B  , ,  wL���]  wL���  w����  w����]  wL���]      B  , ,  y����]  y����  zD���  zD���]  y����]      B  , ,  t����U  t�����  u�����  u����U  t����U      B  , ,  wL���U  wL����  w�����  w����U  wL���U      B  , ,  y����U  y�����  zD����  zD���U  y����U      B  , ,  {����U  {�����  |�����  |����U  {����U      B  , ,  ~6���U  ~6����  ~�����  ~����U  ~6���U      B  , ,  �����U  ������  �.����  �.���U  �����U      B  , ,  �����U  ������  �|����  �|���U  �����U      B  , ,  � ���U  � ����  ������  �����U  � ���U      B  , ,  �n���U  �n����  �����  ����U  �n���U      B  , ,  {����]  {����  |����  |����]  {����]      B  , ,  ~6���]  ~6���  ~����  ~����]  ~6���]      B  , ,  �����]  �����  �.���  �.���]  �����]      B  , ,  �����]  �����  �|���  �|���]  �����]      B  , ,  � ���]  � ���  �����  �����]  � ���]      B  , ,  �n���]  �n���  ����  ����]  �n���]      B  , ,  �����  �����[  �.���[  �.���  �����      B  , ,  �����  �����[  �|���[  �|���  �����      B  , ,  � ���  � ���[  �����[  �����  � ���      B  , ,  �n���  �n���[  ����[  ����  �n���      B  , ,  �����  �����W  �|���W  �|���  �����      B  , ,  � ���  � ���W  �����W  �����  � ���      B  , ,  �n���  �n���W  ����W  ����  �n���      B  , ,  t����  t����W  u����W  u����  t����      B  , ,  wL���  wL���W  w����W  w����  wL���      B  , ,  y����  y����W  zD���W  zD���  y����      B  , ,  {����  {����W  |����W  |����  {����      B  , ,  ~6���  ~6���W  ~����W  ~����  ~6���      B  , ,  t����Y  t����  u����  u����Y  t����Y      B  , ,  wL���Y  wL���  w����  w����Y  wL���Y      B  , ,  y����Y  y����  zD���  zD���Y  y����Y      B  , ,  {����Y  {����  |����  |����Y  {����Y      B  , ,  ~6���Y  ~6���  ~����  ~����Y  ~6���Y      B  , ,  s�����  s����u  t����u  t�����  s�����      B  , ,  v%����  v%���u  v����u  v�����  v%����      B  , ,  xs����  xs���u  y���u  y����  xs����      B  , ,  z�����  z����u  {k���u  {k����  z�����      B  , ,  }����  }���u  }����u  }�����  }����      B  , ,  ]����  ]���u  ����u  �����  ]����      B  , ,  ������  �����u  �U���u  �U����  ������      B  , ,  ������  �����u  �����u  ������  ������      B  , ,  �G����  �G���u  �����u  ������  �G����      B  , ,  ������  �����u  �?���u  �?����  ������      B  , ,  t����  t����  u����  u����  t����      B  , ,  wL���  wL���  w����  w����  wL���      B  , ,  y����  y����  zD���  zD���  y����      B  , ,  {����  {����  |����  |����  {����      B  , ,  ~6���  ~6���  ~����  ~����  ~6���      B  , ,  �����  �����  �.���  �.���  �����      B  , ,  �����  �����  �|���  �|���  �����      B  , ,  � ���  � ���  �����  �����  � ���      B  , ,  r���ڭ  r����W  sZ���W  sZ��ڭ  r���ڭ      B  , ,  r����Y  r����  sZ���  sZ���Y  r����Y      B  , ,  r����  r���د  sZ��د  sZ���  r����      B  , ,  r���ֱ  r����[  sZ���[  sZ��ֱ  r���ֱ      B  , ,  r����]  r����  sZ���  sZ���]  r����]      B  , ,  r����	  r���Գ  sZ��Գ  sZ���	  r����	      B  , ,  ]�����  ]���·  ^t��·  ^t����  ]�����      B  , ,  _����  _��·  _���·  _�����  _����      B  , ,  `r����  `r��·  a��·  a����  `r����      B  , ,  a�����  a���·  bp��·  bp����  a�����      B  , ,  c����  c��·  c���·  c�����  c����      B  , ,  dn����  dn��·  e��·  e����  dn����      B  , ,  e�����  e���·  fl��·  fl����  e�����      B  , ,  g����  g��·  g���·  g�����  g����      B  , ,  hj����  hj��·  i��·  i����  hj����      B  , ,  i�����  i���·  jh��·  jh����  i�����      B  , ,  k����  k��·  k���·  k�����  k����      B  , ,  lf����  lf��·  m��·  m����  lf����      B  , ,  m�����  m���·  nd��·  nd����  m�����      B  , ,  o����  o��·  o���·  o�����  o����      B  , ,  pb����  pb��·  q��·  q����  pb����      B  , ,  q�����  q���·  r`��·  r`����  q�����      B  , ,  s
����  s
��·  s���·  s�����  s
����      B  , ,  t^����  t^��·  u��·  u����  t^����      B  , ,  u�����  u���·  v\��·  v\����  u�����      B  , ,  w����  w��·  w���·  w�����  w����      B  , ,  xZ����  xZ��·  y��·  y����  xZ����      B  , ,  y�����  y���·  zX��·  zX����  y�����      B  , ,  {����  {��·  {���·  {�����  {����      B  , ,  |V����  |V��·  } ��·  } ����  |V����      B  , ,  }�����  }���·  ~T��·  ~T����  }�����      B  , ,  ~�����  ~���·  ���·  �����  ~�����      B  , ,  �R����  �R��·  ����·  ������  �R����      B  , ,  ������  ����·  �P��·  �P����  ������      B  , ,  ������  ����·  ����·  ������  ������      B  , ,  �N����  �N��·  ����·  ������  �N����      B  , ,  ������  ����·  �L��·  �L����  ������      B  , ,  ������  ����·  ����·  ������  ������      B  , ,  �J����  �J��·  ����·  ������  �J����      B  , ,  r����  r���ܫ  sZ��ܫ  sZ���  r����      B  , ,  r���ş  r����I  sZ���I  sZ��ş  r���ş      B  , ,  r����K  r�����  sZ����  sZ���K  r����K      B  , ,  r�����  r���á  sZ��á  sZ����  r�����      B  , ,  r�����  r����M  sZ���M  sZ����  r�����      B  , ,  r����O  r�����  sZ����  sZ���O  r����O      B  , ,  ~6���]  ~6���  ~����  ~����]  ~6���]      B  , ,  �����]  �����  �.���  �.���]  �����]      B  , ,  �����]  �����  �|���  �|���]  �����]      B  , ,  � ���]  � ���  �����  �����]  � ���]      B  , ,  �n���]  �n���  ����  ����]  �n���]      B  , ,  ~6��ڭ  ~6���W  ~����W  ~���ڭ  ~6��ڭ      B  , ,  t����	  t���Գ  u���Գ  u����	  t����	      B  , ,  wL���	  wL��Գ  w���Գ  w����	  wL���	      B  , ,  y����	  y���Գ  zD��Գ  zD���	  y����	      B  , ,  {����	  {���Գ  |���Գ  |����	  {����	      B  , ,  ~6���	  ~6��Գ  ~���Գ  ~����	  ~6���	      B  , ,  �����	  ����Գ  �.��Գ  �.���	  �����	      B  , ,  �����	  ����Գ  �|��Գ  �|���	  �����	      B  , ,  � ���	  � ��Գ  ����Գ  �����	  � ���	      B  , ,  �n���	  �n��Գ  ���Գ  ����	  �n���	      B  , ,  s
��ϕ  s
���?  s����?  s���ϕ  s
��ϕ      B  , ,  t^��ϕ  t^���?  u���?  u��ϕ  t^��ϕ      B  , ,  u���ϕ  u����?  v\���?  v\��ϕ  u���ϕ      B  , ,  w��ϕ  w���?  w����?  w���ϕ  w��ϕ      B  , ,  xZ��ϕ  xZ���?  y���?  y��ϕ  xZ��ϕ      B  , ,  y���ϕ  y����?  zX���?  zX��ϕ  y���ϕ      B  , ,  {��ϕ  {���?  {����?  {���ϕ  {��ϕ      B  , ,  |V��ϕ  |V���?  } ���?  } ��ϕ  |V��ϕ      B  , ,  }���ϕ  }����?  ~T���?  ~T��ϕ  }���ϕ      B  , ,  ~���ϕ  ~����?  ����?  ���ϕ  ~���ϕ      B  , ,  �R��ϕ  �R���?  �����?  ����ϕ  �R��ϕ      B  , ,  ����ϕ  �����?  �P���?  �P��ϕ  ����ϕ      B  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      B  , ,  �N��ϕ  �N���?  �����?  ����ϕ  �N��ϕ      B  , ,  ����ϕ  �����?  �L���?  �L��ϕ  ����ϕ      B  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      B  , ,  �J��ϕ  �J���?  �����?  ����ϕ  �J��ϕ      B  , ,  ����ڭ  �����W  �.���W  �.��ڭ  ����ڭ      B  , ,  ����ڭ  �����W  �|���W  �|��ڭ  ����ڭ      B  , ,  � ��ڭ  � ���W  �����W  ����ڭ  � ��ڭ      B  , ,  �n��ڭ  �n���W  ����W  ���ڭ  �n��ڭ      B  , ,  t���ڭ  t����W  u����W  u���ڭ  t���ڭ      B  , ,  t����Y  t����  u����  u����Y  t����Y      B  , ,  wL���Y  wL���  w����  w����Y  wL���Y      B  , ,  y����Y  y����  zD���  zD���Y  y����Y      B  , ,  {����Y  {����  |����  |����Y  {����Y      B  , ,  ~6���Y  ~6���  ~����  ~����Y  ~6���Y      B  , ,  �����Y  �����  �.���  �.���Y  �����Y      B  , ,  �����Y  �����  �|���  �|���Y  �����Y      B  , ,  � ���Y  � ���  �����  �����Y  � ���Y      B  , ,  �n���Y  �n���  ����  ����Y  �n���Y      B  , ,  wL��ڭ  wL���W  w����W  w���ڭ  wL��ڭ      B  , ,  t����  t���د  u���د  u����  t����      B  , ,  wL���  wL��د  w���د  w����  wL���      B  , ,  y����  y���د  zD��د  zD���  y����      B  , ,  {����  {���د  |���د  |����  {����      B  , ,  ~6���  ~6��د  ~���د  ~����  ~6���      B  , ,  �����  ����د  �.��د  �.���  �����      B  , ,  �����  ����د  �|��د  �|���  �����      B  , ,  � ���  � ��د  ����د  �����  � ���      B  , ,  �n���  �n��د  ���د  ����  �n���      B  , ,  y���ڭ  y����W  zD���W  zD��ڭ  y���ڭ      B  , ,  t���ֱ  t����[  u����[  u���ֱ  t���ֱ      B  , ,  wL��ֱ  wL���[  w����[  w���ֱ  wL��ֱ      B  , ,  y���ֱ  y����[  zD���[  zD��ֱ  y���ֱ      B  , ,  {���ֱ  {����[  |����[  |���ֱ  {���ֱ      B  , ,  ~6��ֱ  ~6���[  ~����[  ~���ֱ  ~6��ֱ      B  , ,  ����ֱ  �����[  �.���[  �.��ֱ  ����ֱ      B  , ,  ����ֱ  �����[  �|���[  �|��ֱ  ����ֱ      B  , ,  � ��ֱ  � ���[  �����[  ����ֱ  � ��ֱ      B  , ,  �n��ֱ  �n���[  ����[  ���ֱ  �n��ֱ      B  , ,  t����  t���ܫ  u���ܫ  u����  t����      B  , ,  wL���  wL��ܫ  w���ܫ  w����  wL���      B  , ,  y����  y���ܫ  zD��ܫ  zD���  y����      B  , ,  {����  {���ܫ  |���ܫ  |����  {����      B  , ,  {���ڭ  {����W  |����W  |���ڭ  {���ڭ      B  , ,  ~6���  ~6��ܫ  ~���ܫ  ~����  ~6���      B  , ,  t����]  t����  u����  u����]  t����]      B  , ,  �����  ����ܫ  �.��ܫ  �.���  �����      B  , ,  wL���]  wL���  w����  w����]  wL���]      B  , ,  �����  ����ܫ  �|��ܫ  �|���  �����      B  , ,  y����]  y����  zD���  zD���]  y����]      B  , ,  � ���  � ��ܫ  ����ܫ  �����  � ���      B  , ,  {����]  {����  |����  |����]  {����]      B  , ,  �n���  �n��ܫ  ���ܫ  ����  �n���      B  , ,  d����Y  d����  e����  e����Y  d����Y      B  , ,  ix���  ix��ܫ  j"��ܫ  j"���  ix���      B  , ,  [�����  [���ӑ  \b��ӑ  \b����  [�����      B  , ,  [���ѓ  [����=  \b���=  \b��ѓ  [���ѓ      B  , ,  ]���ϕ  ]����?  ^t���?  ^t��ϕ  ]���ϕ      B  , ,  _��ϕ  _���?  _����?  _���ϕ  _��ϕ      B  , ,  `r��ϕ  `r���?  a���?  a��ϕ  `r��ϕ      B  , ,  a���ϕ  a����?  bp���?  bp��ϕ  a���ϕ      B  , ,  c��ϕ  c���?  c����?  c���ϕ  c��ϕ      B  , ,  dn��ϕ  dn���?  e���?  e��ϕ  dn��ϕ      B  , ,  e���ϕ  e����?  fl���?  fl��ϕ  e���ϕ      B  , ,  g��ϕ  g���?  g����?  g���ϕ  g��ϕ      B  , ,  hj��ϕ  hj���?  i���?  i��ϕ  hj��ϕ      B  , ,  i���ϕ  i����?  jh���?  jh��ϕ  i���ϕ      B  , ,  k��ϕ  k���?  k����?  k���ϕ  k��ϕ      B  , ,  lf��ϕ  lf���?  m���?  m��ϕ  lf��ϕ      B  , ,  m���ϕ  m����?  nd���?  nd��ϕ  m���ϕ      B  , ,  o��ϕ  o���?  o����?  o���ϕ  o��ϕ      B  , ,  pb��ϕ  pb���?  q���?  q��ϕ  pb��ϕ      B  , ,  q���ϕ  q����?  r`���?  r`��ϕ  q���ϕ      B  , ,  g*���Y  g*���  g����  g����Y  g*���Y      B  , ,  ix���Y  ix���  j"���  j"���Y  ix���Y      B  , ,  k����Y  k����  lp���  lp���Y  k����Y      B  , ,  b����  b���ܫ  c8��ܫ  c8���  b����      B  , ,  [�����  [���׍  \b��׍  \b����  [�����      B  , ,  ]���ֱ  ]����[  ^����[  ^���ֱ  ]���ֱ      B  , ,  `@��ֱ  `@���[  `����[  `���ֱ  `@��ֱ      B  , ,  b���ֱ  b����[  c8���[  c8��ֱ  b���ֱ      B  , ,  d���ֱ  d����[  e����[  e���ֱ  d���ֱ      B  , ,  g*��ֱ  g*���[  g����[  g���ֱ  g*��ֱ      B  , ,  ix��ֱ  ix���[  j"���[  j"��ֱ  ix��ֱ      B  , ,  k���ֱ  k����[  lp���[  lp��ֱ  k���ֱ      B  , ,  n��ֱ  n���[  n����[  n���ֱ  n��ֱ      B  , ,  pb��ֱ  pb���[  q���[  q��ֱ  pb��ֱ      B  , ,  n���Y  n���  n����  n����Y  n���Y      B  , ,  pb���Y  pb���  q���  q���Y  pb���Y      B  , ,  pb��ڭ  pb���W  q���W  q��ڭ  pb��ڭ      B  , ,  k����  k���ܫ  lp��ܫ  lp���  k����      B  , ,  n���  n��ܫ  n���ܫ  n����  n���      B  , ,  [����3  [�����  \b����  \b���3  [����3      B  , ,  [�����  [���ۉ  \b��ۉ  \b����  [�����      B  , ,  ]���ڭ  ]����W  ^����W  ^���ڭ  ]���ڭ      B  , ,  `@��ڭ  `@���W  `����W  `���ڭ  `@��ڭ      B  , ,  b���ڭ  b����W  c8���W  c8��ڭ  b���ڭ      B  , ,  d���ڭ  d����W  e����W  e���ڭ  d���ڭ      B  , ,  g*��ڭ  g*���W  g����W  g���ڭ  g*��ڭ      B  , ,  d����  d���ܫ  e���ܫ  e����  d����      B  , ,  [���Տ  [����9  \b���9  \b��Տ  [���Տ      B  , ,  ]����]  ]����  ^����  ^����]  ]����]      B  , ,  `@���]  `@���  `����  `����]  `@���]      B  , ,  b����]  b����  c8���  c8���]  b����]      B  , ,  d����]  d����  e����  e����]  d����]      B  , ,  g*���]  g*���  g����  g����]  g*���]      B  , ,  ix���]  ix���  j"���  j"���]  ix���]      B  , ,  k����]  k����  lp���  lp���]  k����]      B  , ,  n���]  n���  n����  n����]  n���]      B  , ,  pb���]  pb���  q���  q���]  pb���]      B  , ,  ix��ڭ  ix���W  j"���W  j"��ڭ  ix��ڭ      B  , ,  k���ڭ  k����W  lp���W  lp��ڭ  k���ڭ      B  , ,  `@���  `@��ܫ  `���ܫ  `����  `@���      B  , ,  [����7  [�����  \b����  \b���7  [����7      B  , ,  ]����  ]���د  ^���د  ^����  ]����      B  , ,  `@���  `@��د  `���د  `����  `@���      B  , ,  b����  b���د  c8��د  c8���  b����      B  , ,  d����  d���د  e���د  e����  d����      B  , ,  g*���  g*��د  g���د  g����  g*���      B  , ,  ix���  ix��د  j"��د  j"���  ix���      B  , ,  g*���  g*��ܫ  g���ܫ  g����  g*���      B  , ,  [����;  [�����  \b����  \b���;  [����;      B  , ,  ]����	  ]���Գ  ^���Գ  ^����	  ]����	      B  , ,  `@���	  `@��Գ  `���Գ  `����	  `@���	      B  , ,  b����	  b���Գ  c8��Գ  c8���	  b����	      B  , ,  pb���  pb��ܫ  q��ܫ  q���  pb���      B  , ,  d����	  d���Գ  e���Գ  e����	  d����	      B  , ,  g*���	  g*��Գ  g���Գ  g����	  g*���	      B  , ,  ix���	  ix��Գ  j"��Գ  j"���	  ix���	      B  , ,  k����	  k���Գ  lp��Գ  lp���	  k����	      B  , ,  n���	  n��Գ  n���Գ  n����	  n���	      B  , ,  pb���	  pb��Գ  q��Գ  q���	  pb���	      B  , ,  k����  k���د  lp��د  lp���  k����      B  , ,  n���  n��د  n���د  n����  n���      B  , ,  pb���  pb��د  q��د  q���  pb���      B  , ,  n��ڭ  n���W  n����W  n���ڭ  n��ڭ      B  , ,  ]����  ]���ܫ  ^���ܫ  ^����  ]����      B  , ,  [���ً  [����5  \b���5  \b��ً  [���ً      B  , ,  ]����Y  ]����  ^����  ^����Y  ]����Y      B  , ,  `@���Y  `@���  `����  `����Y  `@���Y      B  , ,  b����Y  b����  c8���  c8���Y  b����Y      B  , ,  pb���%  pb����  q����  q���%  pb���%      B  , ,  q����%  q�����  r`����  r`���%  q����%      B  , ,  ]����%  ]�����  ^t����  ^t���%  ]����%      B  , ,  _���%  _����  _�����  _����%  _���%      B  , ,  ]����  ]���ʽ  ^t��ʽ  ^t���  ]����      B  , ,  _���  _��ʽ  _���ʽ  _����  _���      B  , ,  `r���  `r��ʽ  a��ʽ  a���  `r���      B  , ,  a����  a���ʽ  bp��ʽ  bp���  a����      B  , ,  c���  c��ʽ  c���ʽ  c����  c���      B  , ,  dn���  dn��ʽ  e��ʽ  e���  dn���      B  , ,  e����  e���ʽ  fl��ʽ  fl���  e����      B  , ,  g���  g��ʽ  g���ʽ  g����  g���      B  , ,  hj���  hj��ʽ  i��ʽ  i���  hj���      B  , ,  i����  i���ʽ  jh��ʽ  jh���  i����      B  , ,  k���  k��ʽ  k���ʽ  k����  k���      B  , ,  lf���  lf��ʽ  m��ʽ  m���  lf���      B  , ,  m����  m���ʽ  nd��ʽ  nd���  m����      B  , ,  o���  o��ʽ  o���ʽ  o����  o���      B  , ,  pb���  pb��ʽ  q��ʽ  q���  pb���      B  , ,  q����  q���ʽ  r`��ʽ  r`���  q����      B  , ,  `r���%  `r����  a����  a���%  `r���%      B  , ,  a����%  a�����  bp����  bp���%  a����%      B  , ,  [����  [���ȿ  \b��ȿ  \b���  [����      B  , ,  [�����  [����k  \b���k  \b����  [�����      B  , ,  [����m  [����  \b���  \b���m  [����m      B  , ,  ]���ş  ]����I  ^����I  ^���ş  ]���ş      B  , ,  `@��ş  `@���I  `����I  `���ş  `@��ş      B  , ,  b���ş  b����I  c8���I  c8��ş  b���ş      B  , ,  d���ş  d����I  e����I  e���ş  d���ş      B  , ,  g*��ş  g*���I  g����I  g���ş  g*��ş      B  , ,  ix��ş  ix���I  j"���I  j"��ş  ix��ş      B  , ,  k���ş  k����I  lp���I  lp��ş  k���ş      B  , ,  n��ş  n���I  n����I  n���ş  n��ş      B  , ,  pb��ş  pb���I  q���I  q��ş  pb��ş      B  , ,  c���%  c����  c�����  c����%  c���%      B  , ,  dn���%  dn����  e����  e���%  dn���%      B  , ,  [����  [�����  \b����  \b���  [����      B  , ,  ]����K  ]�����  ^�����  ^����K  ]����K      B  , ,  `@���K  `@����  `�����  `����K  `@���K      B  , ,  b����K  b�����  c8����  c8���K  b����K      B  , ,  d����K  d�����  e�����  e����K  d����K      B  , ,  g*���K  g*����  g�����  g����K  g*���K      B  , ,  ix���K  ix����  j"����  j"���K  ix���K      B  , ,  k����K  k�����  lp����  lp���K  k����K      B  , ,  n���K  n����  n�����  n����K  n���K      B  , ,  pb���K  pb����  q����  q���K  pb���K      B  , ,  e����%  e�����  fl����  fl���%  e����%      B  , ,  g���%  g����  g�����  g����%  g���%      B  , ,  [�����  [����o  \b���o  \b����  [�����      B  , ,  ]�����  ]���á  ^���á  ^�����  ]�����      B  , ,  `@����  `@��á  `���á  `�����  `@����      B  , ,  b�����  b���á  c8��á  c8����  b�����      B  , ,  d�����  d���á  e���á  e�����  d�����      B  , ,  g*����  g*��á  g���á  g�����  g*����      B  , ,  ix����  ix��á  j"��á  j"����  ix����      B  , ,  k�����  k���á  lp��á  lp����  k�����      B  , ,  n����  n��á  n���á  n�����  n����      B  , ,  pb����  pb��á  q��á  q����  pb����      B  , ,  hj���%  hj����  i����  i���%  hj���%      B  , ,  i����%  i�����  jh����  jh���%  i����%      B  , ,  [����q  [����  \b���  \b���q  [����q      B  , ,  ]�����  ]����M  ^����M  ^�����  ]�����      B  , ,  `@����  `@���M  `����M  `�����  `@����      B  , ,  b�����  b����M  c8���M  c8����  b�����      B  , ,  d�����  d����M  e����M  e�����  d�����      B  , ,  g*����  g*���M  g����M  g�����  g*����      B  , ,  ix����  ix���M  j"���M  j"����  ix����      B  , ,  k�����  k����M  lp���M  lp����  k�����      B  , ,  n����  n���M  n����M  n�����  n����      B  , ,  pb����  pb���M  q���M  q����  pb����      B  , ,  k���%  k����  k�����  k����%  k���%      B  , ,  lf���%  lf����  m����  m���%  lf���%      B  , ,  [����  [�����  \b����  \b���  [����      B  , ,  ]����O  ]�����  ^�����  ^����O  ]����O      B  , ,  `@���O  `@����  `�����  `����O  `@���O      B  , ,  b����O  b�����  c8����  c8���O  b����O      B  , ,  d����O  d�����  e�����  e����O  d����O      B  , ,  g*���O  g*����  g�����  g����O  g*���O      B  , ,  ix���O  ix����  j"����  j"���O  ix���O      B  , ,  k����O  k�����  lp����  lp���O  k����O      B  , ,  n���O  n����  n�����  n����O  n���O      B  , ,  pb���O  pb����  q����  q���O  pb���O      B  , ,  m����%  m�����  nd����  nd���%  m����%      B  , ,  o���%  o����  o�����  o����%  o���%      B  , ,  xZ���  xZ��ʽ  y��ʽ  y���  xZ���      B  , ,  y����  y���ʽ  zX��ʽ  zX���  y����      B  , ,  {���  {��ʽ  {���ʽ  {����  {���      B  , ,  |V���  |V��ʽ  } ��ʽ  } ���  |V���      B  , ,  }����  }���ʽ  ~T��ʽ  ~T���  }����      B  , ,  ~����  ~���ʽ  ���ʽ  ����  ~����      B  , ,  t����K  t�����  u�����  u����K  t����K      B  , ,  wL���K  wL����  w�����  w����K  wL���K      B  , ,  y����K  y�����  zD����  zD���K  y����K      B  , ,  {����K  {�����  |�����  |����K  {����K      B  , ,  ~6���K  ~6����  ~�����  ~����K  ~6���K      B  , ,  �����K  ������  �.����  �.���K  �����K      B  , ,  �����K  ������  �|����  �|���K  �����K      B  , ,  � ���K  � ����  ������  �����K  � ���K      B  , ,  �n���K  �n����  �����  ����K  �n���K      B  , ,  �R���  �R��ʽ  ����ʽ  �����  �R���      B  , ,  �����  ����ʽ  �P��ʽ  �P���  �����      B  , ,  �����  ����ʽ  ����ʽ  �����  �����      B  , ,  �N���  �N��ʽ  ����ʽ  �����  �N���      B  , ,  �����  ����ʽ  �L��ʽ  �L���  �����      B  , ,  �����  ����ʽ  ����ʽ  �����  �����      B  , ,  �J���  �J��ʽ  ����ʽ  �����  �J���      B  , ,  t^���%  t^����  u����  u���%  t^���%      B  , ,  u����%  u�����  v\����  v\���%  u����%      B  , ,  w���%  w����  w�����  w����%  w���%      B  , ,  xZ���%  xZ����  y����  y���%  xZ���%      B  , ,  y����%  y�����  zX����  zX���%  y����%      B  , ,  t�����  t���á  u���á  u�����  t�����      B  , ,  wL����  wL��á  w���á  w�����  wL����      B  , ,  y�����  y���á  zD��á  zD����  y�����      B  , ,  {�����  {���á  |���á  |�����  {�����      B  , ,  ~6����  ~6��á  ~���á  ~�����  ~6����      B  , ,  ������  ����á  �.��á  �.����  ������      B  , ,  ������  ����á  �|��á  �|����  ������      B  , ,  � ����  � ��á  ����á  ������  � ����      B  , ,  �n����  �n��á  ���á  �����  �n����      B  , ,  {���%  {����  {�����  {����%  {���%      B  , ,  |V���%  |V����  } ����  } ���%  |V���%      B  , ,  }����%  }�����  ~T����  ~T���%  }����%      B  , ,  ~����%  ~�����  �����  ����%  ~����%      B  , ,  �R���%  �R����  ������  �����%  �R���%      B  , ,  �����%  ������  �P����  �P���%  �����%      B  , ,  �����%  ������  ������  �����%  �����%      B  , ,  �N���%  �N����  ������  �����%  �N���%      B  , ,  �����%  ������  �L����  �L���%  �����%      B  , ,  �����%  ������  ������  �����%  �����%      B  , ,  t���ş  t����I  u����I  u���ş  t���ş      B  , ,  wL��ş  wL���I  w����I  w���ş  wL��ş      B  , ,  t�����  t����M  u����M  u�����  t�����      B  , ,  wL����  wL���M  w����M  w�����  wL����      B  , ,  y�����  y����M  zD���M  zD����  y�����      B  , ,  {�����  {����M  |����M  |�����  {�����      B  , ,  ~6����  ~6���M  ~����M  ~�����  ~6����      B  , ,  ������  �����M  �.���M  �.����  ������      B  , ,  ������  �����M  �|���M  �|����  ������      B  , ,  � ����  � ���M  �����M  ������  � ����      B  , ,  �n����  �n���M  ����M  �����  �n����      B  , ,  y���ş  y����I  zD���I  zD��ş  y���ş      B  , ,  {���ş  {����I  |����I  |���ş  {���ş      B  , ,  ~6��ş  ~6���I  ~����I  ~���ş  ~6��ş      B  , ,  ����ş  �����I  �.���I  �.��ş  ����ş      B  , ,  ����ş  �����I  �|���I  �|��ş  ����ş      B  , ,  � ��ş  � ���I  �����I  ����ş  � ��ş      B  , ,  �n��ş  �n���I  ����I  ���ş  �n��ş      B  , ,  �J���%  �J����  ������  �����%  �J���%      B  , ,  s
���%  s
����  s�����  s����%  s
���%      B  , ,  s
���  s
��ʽ  s���ʽ  s����  s
���      B  , ,  t^���  t^��ʽ  u��ʽ  u���  t^���      B  , ,  u����  u���ʽ  v\��ʽ  v\���  u����      B  , ,  t����O  t�����  u�����  u����O  t����O      B  , ,  wL���O  wL����  w�����  w����O  wL���O      B  , ,  y����O  y�����  zD����  zD���O  y����O      B  , ,  {����O  {�����  |�����  |����O  {����O      B  , ,  ~6���O  ~6����  ~�����  ~����O  ~6���O      B  , ,  �����O  ������  �.����  �.���O  �����O      B  , ,  �����O  ������  �|����  �|���O  �����O      B  , ,  � ���O  � ����  ������  �����O  � ���O      B  , ,  �n���O  �n����  �����  ����O  �n���O      B  , ,  w���  w��ʽ  w���ʽ  w����  w���      B  , ,  �B����  �B��·  ����·  ������  �B����      B  , ,  ������  ����·  �@��·  �@����  ������      B  , ,  ������  ����·  ����·  ������  ������      B  , ,  �>����  �>��·  ����·  ������  �>����      B  , ,  ������  ����·  �<��·  �<����  ������      B  , ,  ������  ����·  ����·  ������  ������      B  , ,  �:����  �:��·  ����·  ������  �:����      B  , ,  ������  ����·  �8��·  �8����  ������      B  , ,  ������  ����·  ����·  ������  ������      B  , ,  �6����  �6��·  ����·  ������  �6����      B  , ,  ������  ����·  �4��·  �4����  ������      B  , ,  ������  ����·  ����·  ������  ������      B  , ,  �2����  �2��·  ����·  ������  �2����      B  , ,  ������  ����·  �0��·  �0����  ������      B  , ,  ������  ����·  ����·  ������  ������      B  , ,  �.����  �.��·  ����·  ������  �.����      B  , ,  ������  ����·  �,��·  �,����  ������      B  , ,  ������  ����·  ����·  ������  ������      B  , ,  �*����  �*��·  ����·  ������  �*����      B  , ,  �~����  �~��·  �(��·  �(����  �~����      B  , ,  ������  ����·  �|��·  �|����  ������      B  , ,  �&����  �&��·  ����·  ������  �&����      B  , ,  �z����  �z��·  �$��·  �$����  �z����      B  , ,  ������  ����·  �x��·  �x����  ������      B  , ,  �"����  �"��·  ����·  ������  �"����      B  , ,  �v����  �v��·  � ��·  � ����  �v����      B  , ,  ������  ����·  �t��·  �t����  ������      B  , ,  �����  ���·  ����·  ������  �����      B  , ,  �r����  �r��·  ���·  �����  �r����      B  , ,  ������  ����·  �p��·  �p����  ������      B  , ,  �����]  �����  �r���  �r���]  �����]      B  , ,  ����ڭ  �����W  �r���W  �r��ڭ  ����ڭ      B  , ,  �����	  ����Գ  �r��Գ  �r���	  �����	      B  , ,  �����  ����د  �r��د  �r���  �����      B  , ,  �����  ����ܫ  �r��ܫ  �r���  �����      B  , ,  ����ş  �����I  �r���I  �r��ş  ����ş      B  , ,  �����K  ������  �r����  �r���K  �����K      B  , ,  ������  ����á  �r��á  �r����  ������      B  , ,  ����ֱ  �����[  �r���[  �r��ֱ  ����ֱ      B  , ,  ������  �����M  �r���M  �r����  ������      B  , ,  �����Y  �����  �r���  �r���Y  �����Y      B  , ,  ������  ����·  ����·  ������  ������      B  , ,  �F����  �F��·  ����·  ������  �F����      B  , ,  ������  ����·  �D��·  �D����  ������      B  , ,  ������  ����·  ����·  ������  ������      B  , ,  �����O  ������  �r����  �r���O  �����O      B  , ,  �����Y  �����  �����  �����Y  �����Y      B  , ,  ���ڭ  ����W  �����W  ����ڭ  ���ڭ      B  , ,  �d��ڭ  �d���W  ����W  ���ڭ  �d��ڭ      B  , ,  ����ڭ  �����W  �\���W  �\��ڭ  ����ڭ      B  , ,  � ��ڭ  � ���W  �����W  ����ڭ  � ��ڭ      B  , ,  �N��ڭ  �N���W  �����W  ����ڭ  �N��ڭ      B  , ,  ����ڭ  �����W  �F���W  �F��ڭ  ����ڭ      B  , ,  ����ڭ  �����W  �����W  ����ڭ  ����ڭ      B  , ,  �8��ڭ  �8���W  �����W  ����ڭ  �8��ڭ      B  , ,  ����ڭ  �����W  �0���W  �0��ڭ  ����ڭ      B  , ,  ����ڭ  �����W  �~���W  �~��ڭ  ����ڭ      B  , ,  �8���Y  �8���  �����  �����Y  �8���Y      B  , ,  ����	  ���Գ  ����Գ  �����	  ����	      B  , ,  �d���	  �d��Գ  ���Գ  ����	  �d���	      B  , ,  �����	  ����Գ  �\��Գ  �\���	  �����	      B  , ,  � ���	  � ��Գ  ����Գ  �����	  � ���	      B  , ,  �N���	  �N��Գ  ����Գ  �����	  �N���	      B  , ,  �����	  ����Գ  �F��Գ  �F���	  �����	      B  , ,  �����	  ����Գ  ����Գ  �����	  �����	      B  , ,  �8���	  �8��Գ  ����Գ  �����	  �8���	      B  , ,  �����	  ����Գ  �0��Գ  �0���	  �����	      B  , ,  �����	  ����Գ  �~��Գ  �~���	  �����	      B  , ,  �����Y  �����  �0���  �0���Y  �����Y      B  , ,  ����  ���د  ����د  �����  ����      B  , ,  �d���  �d��د  ���د  ����  �d���      B  , ,  �����  ����د  �\��د  �\���  �����      B  , ,  � ���  � ��د  ����د  �����  � ���      B  , ,  �N���  �N��د  ����د  �����  �N���      B  , ,  �����  ����د  �F��د  �F���  �����      B  , ,  �����  ����د  ����د  �����  �����      B  , ,  �8���  �8��د  ����د  �����  �8���      B  , ,  �����  ����د  �0��د  �0���  �����      B  , ,  �����  ����د  �~��د  �~���  �����      B  , ,  �����Y  �����  �~���  �~���Y  �����Y      B  , ,  ����  ���ܫ  ����ܫ  �����  ����      B  , ,  �����Y  �����  �F���  �F���Y  �����Y      B  , ,  �d���  �d��ܫ  ���ܫ  ����  �d���      B  , ,  �����  ����ܫ  �\��ܫ  �\���  �����      B  , ,  � ���  � ��ܫ  ����ܫ  �����  � ���      B  , ,  �N���  �N��ܫ  ����ܫ  �����  �N���      B  , ,  �����  ����ܫ  �F��ܫ  �F���  �����      B  , ,  �����  ����ܫ  ����ܫ  �����  �����      B  , ,  �8���  �8��ܫ  ����ܫ  �����  �8���      B  , ,  �����  ����ܫ  �0��ܫ  �0���  �����      B  , ,  �����  ����ܫ  �~��ܫ  �~���  �����      B  , ,  ����]  ����  �����  �����]  ����]      B  , ,  ����ϕ  �����?  �0���?  �0��ϕ  ����ϕ      B  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      B  , ,  �.��ϕ  �.���?  �����?  ����ϕ  �.��ϕ      B  , ,  ����ϕ  �����?  �,���?  �,��ϕ  ����ϕ      B  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      B  , ,  �*��ϕ  �*���?  �����?  ����ϕ  �*��ϕ      B  , ,  �~��ϕ  �~���?  �(���?  �(��ϕ  �~��ϕ      B  , ,  ����ϕ  �����?  �|���?  �|��ϕ  ����ϕ      B  , ,  �&��ϕ  �&���?  �����?  ����ϕ  �&��ϕ      B  , ,  �z��ϕ  �z���?  �$���?  �$��ϕ  �z��ϕ      B  , ,  ����ϕ  �����?  �x���?  �x��ϕ  ����ϕ      B  , ,  �"��ϕ  �"���?  �����?  ����ϕ  �"��ϕ      B  , ,  �v��ϕ  �v���?  � ���?  � ��ϕ  �v��ϕ      B  , ,  ����ϕ  �����?  �t���?  �t��ϕ  ����ϕ      B  , ,  �d���]  �d���  ����  ����]  �d���]      B  , ,  ���ϕ  ����?  �����?  ����ϕ  ���ϕ      B  , ,  �r��ϕ  �r���?  ����?  ���ϕ  �r��ϕ      B  , ,  ����ϕ  �����?  �p���?  �p��ϕ  ����ϕ      B  , ,  �����]  �����  �\���  �\���]  �����]      B  , ,  ���ֱ  ����[  �����[  ����ֱ  ���ֱ      B  , ,  �d��ֱ  �d���[  ����[  ���ֱ  �d��ֱ      B  , ,  ����ֱ  �����[  �\���[  �\��ֱ  ����ֱ      B  , ,  � ��ֱ  � ���[  �����[  ����ֱ  � ��ֱ      B  , ,  �N��ֱ  �N���[  �����[  ����ֱ  �N��ֱ      B  , ,  ����ֱ  �����[  �F���[  �F��ֱ  ����ֱ      B  , ,  � ���]  � ���  �����  �����]  � ���]      B  , ,  ����ֱ  �����[  �����[  ����ֱ  ����ֱ      B  , ,  �8��ֱ  �8���[  �����[  ����ֱ  �8��ֱ      B  , ,  ����ֱ  �����[  �0���[  �0��ֱ  ����ֱ      B  , ,  ����ֱ  �����[  �~���[  �~��ֱ  ����ֱ      B  , ,  �N���]  �N���  �����  �����]  �N���]      B  , ,  ����Y  ����  �����  �����Y  ����Y      B  , ,  �d���Y  �d���  ����  ����Y  �d���Y      B  , ,  �����Y  �����  �\���  �\���Y  �����Y      B  , ,  � ���Y  � ���  �����  �����Y  � ���Y      B  , ,  �N���Y  �N���  �����  �����Y  �N���Y      B  , ,  �����]  �����  �F���  �F���]  �����]      B  , ,  �����]  �����  �����  �����]  �����]      B  , ,  �8���]  �8���  �����  �����]  �8���]      B  , ,  �����]  �����  �0���  �0���]  �����]      B  , ,  �����]  �����  �~���  �~���]  �����]      B  , ,  ����ڭ  �����W  �:���W  �:��ڭ  ����ڭ      B  , ,  �
���  �
��ܫ  ����ܫ  �����  �
���      B  , ,  �
��ڭ  �
���W  �����W  ����ڭ  �
��ڭ      B  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      B  , ,  �F��ϕ  �F���?  �����?  ����ϕ  �F��ϕ      B  , ,  ����ϕ  �����?  �D���?  �D��ϕ  ����ϕ      B  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      B  , ,  �B��ϕ  �B���?  �����?  ����ϕ  �B��ϕ      B  , ,  ����ϕ  �����?  �@���?  �@��ϕ  ����ϕ      B  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      B  , ,  �>��ϕ  �>���?  �����?  ����ϕ  �>��ϕ      B  , ,  ����ϕ  �����?  �<���?  �<��ϕ  ����ϕ      B  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      B  , ,  ����ڭ  �����W  �����W  ����ڭ  ����ڭ      B  , ,  �:��ϕ  �:���?  �����?  ����ϕ  �:��ϕ      B  , ,  ����ϕ  �����?  �8���?  �8��ϕ  ����ϕ      B  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      B  , ,  �6��ϕ  �6���?  �����?  ����ϕ  �6��ϕ      B  , ,  ����ϕ  �����?  �4���?  �4��ϕ  ����ϕ      B  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      B  , ,  �2��ϕ  �2���?  �����?  ����ϕ  �2��ϕ      B  , ,  �,��ڭ  �,���W  �����W  ����ڭ  �,��ڭ      B  , ,  �z��ڭ  �z���W  �$���W  �$��ڭ  �z��ڭ      B  , ,  �z���]  �z���  �$���  �$���]  �z���]      B  , ,  �X��ڭ  �X���W  ����W  ���ڭ  �X��ڭ      B  , ,  ����ڭ  �����W  �P���W  �P��ڭ  ����ڭ      B  , ,  ����ڭ  �����W  �����W  ����ڭ  ����ڭ      B  , ,  �
���]  �
���  �����  �����]  �
���]      B  , ,  �����  ����د  ����د  �����  �����      B  , ,  �B���  �B��د  ����د  �����  �B���      B  , ,  �����  ����د  �:��د  �:���  �����      B  , ,  �����  ����د  ����د  �����  �����      B  , ,  �,���  �,��د  ����د  �����  �,���      B  , ,  �z���  �z��د  �$��د  �$���  �z���      B  , ,  �X���]  �X���  ����  ����]  �X���]      B  , ,  �����]  �����  �P���  �P���]  �����]      B  , ,  �����]  �����  �����  �����]  �����]      B  , ,  �B���]  �B���  �����  �����]  �B���]      B  , ,  �����]  �����  �:���  �:���]  �����]      B  , ,  �
���Y  �
���  �����  �����Y  �
���Y      B  , ,  �X���Y  �X���  ����  ����Y  �X���Y      B  , ,  �
��ֱ  �
���[  �����[  ����ֱ  �
��ֱ      B  , ,  �X��ֱ  �X���[  ����[  ���ֱ  �X��ֱ      B  , ,  ����ֱ  �����[  �P���[  �P��ֱ  ����ֱ      B  , ,  ����ֱ  �����[  �����[  ����ֱ  ����ֱ      B  , ,  �B��ֱ  �B���[  �����[  ����ֱ  �B��ֱ      B  , ,  ����ֱ  �����[  �:���[  �:��ֱ  ����ֱ      B  , ,  ����ֱ  �����[  �����[  ����ֱ  ����ֱ      B  , ,  �,��ֱ  �,���[  �����[  ����ֱ  �,��ֱ      B  , ,  �z��ֱ  �z���[  �$���[  �$��ֱ  �z��ֱ      B  , ,  �����]  �����  �����  �����]  �����]      B  , ,  �X���  �X��ܫ  ���ܫ  ����  �X���      B  , ,  �����  ����ܫ  �P��ܫ  �P���  �����      B  , ,  �
���  �
��د  ����د  �����  �
���      B  , ,  �X���  �X��د  ���د  ����  �X���      B  , ,  �����  ����د  �P��د  �P���  �����      B  , ,  �����  ����ܫ  ����ܫ  �����  �����      B  , ,  �B���  �B��ܫ  ����ܫ  �����  �B���      B  , ,  �����  ����ܫ  �:��ܫ  �:���  �����      B  , ,  �����  ����ܫ  ����ܫ  �����  �����      B  , ,  �,���  �,��ܫ  ����ܫ  �����  �,���      B  , ,  �z���  �z��ܫ  �$��ܫ  �$���  �z���      B  , ,  �����Y  �����  �P���  �P���Y  �����Y      B  , ,  �����Y  �����  �����  �����Y  �����Y      B  , ,  �B���Y  �B���  �����  �����Y  �B���Y      B  , ,  �����Y  �����  �:���  �:���Y  �����Y      B  , ,  �����Y  �����  �����  �����Y  �����Y      B  , ,  �,���Y  �,���  �����  �����Y  �,���Y      B  , ,  �z���Y  �z���  �$���  �$���Y  �z���Y      B  , ,  �
���	  �
��Գ  ����Գ  �����	  �
���	      B  , ,  �X���	  �X��Գ  ���Գ  ����	  �X���	      B  , ,  �����	  ����Գ  �P��Գ  �P���	  �����	      B  , ,  �����	  ����Գ  ����Գ  �����	  �����	      B  , ,  �B���	  �B��Գ  ����Գ  �����	  �B���	      B  , ,  �����	  ����Գ  �:��Գ  �:���	  �����	      B  , ,  �����	  ����Գ  ����Գ  �����	  �����	      B  , ,  �,���	  �,��Գ  ����Գ  �����	  �,���	      B  , ,  �z���	  �z��Գ  �$��Գ  �$���	  �z���	      B  , ,  �,���]  �,���  �����  �����]  �,���]      B  , ,  �B��ڭ  �B���W  �����W  ����ڭ  �B��ڭ      B  , ,  ����ş  �����I  �����I  ����ş  ����ş      B  , ,  �B��ş  �B���I  �����I  ����ş  �B��ş      B  , ,  ����ş  �����I  �:���I  �:��ş  ����ş      B  , ,  ����ş  �����I  �����I  ����ş  ����ş      B  , ,  �,��ş  �,���I  �����I  ����ş  �,��ş      B  , ,  �z��ş  �z���I  �$���I  �$��ş  �z��ş      B  , ,  �>���  �>��ʽ  ����ʽ  �����  �>���      B  , ,  �
����  �
��á  ����á  ������  �
����      B  , ,  �X����  �X��á  ���á  �����  �X����      B  , ,  ������  ����á  �P��á  �P����  ������      B  , ,  ������  ����á  ����á  ������  ������      B  , ,  �B����  �B��á  ����á  ������  �B����      B  , ,  ������  ����á  �:��á  �:����  ������      B  , ,  ������  ����á  ����á  ������  ������      B  , ,  �,����  �,��á  ����á  ������  �,����      B  , ,  �z����  �z��á  �$��á  �$����  �z����      B  , ,  �����  ����ʽ  �<��ʽ  �<���  �����      B  , ,  �����  ����ʽ  ����ʽ  �����  �����      B  , ,  �:���  �:��ʽ  ����ʽ  �����  �:���      B  , ,  �����  ����ʽ  �8��ʽ  �8���  �����      B  , ,  �����  ����ʽ  ����ʽ  �����  �����      B  , ,  �6���  �6��ʽ  ����ʽ  �����  �6���      B  , ,  �����  ����ʽ  �4��ʽ  �4���  �����      B  , ,  �����  ����ʽ  ����ʽ  �����  �����      B  , ,  �2���  �2��ʽ  ����ʽ  �����  �2���      B  , ,  �F���%  �F����  ������  �����%  �F���%      B  , ,  �����%  ������  �D����  �D���%  �����%      B  , ,  �����%  ������  ������  �����%  �����%      B  , ,  �B���%  �B����  ������  �����%  �B���%      B  , ,  �����%  ������  �@����  �@���%  �����%      B  , ,  �����%  ������  ������  �����%  �����%      B  , ,  �>���%  �>����  ������  �����%  �>���%      B  , ,  �����%  ������  �<����  �<���%  �����%      B  , ,  �����%  ������  ������  �����%  �����%      B  , ,  �:���%  �:����  ������  �����%  �:���%      B  , ,  �����%  ������  �8����  �8���%  �����%      B  , ,  �����%  ������  ������  �����%  �����%      B  , ,  �
���K  �
����  ������  �����K  �
���K      B  , ,  �
����  �
���M  �����M  ������  �
����      B  , ,  �X����  �X���M  ����M  �����  �X����      B  , ,  ������  �����M  �P���M  �P����  ������      B  , ,  ������  �����M  �����M  ������  ������      B  , ,  �B����  �B���M  �����M  ������  �B����      B  , ,  ������  �����M  �:���M  �:����  ������      B  , ,  ������  �����M  �����M  ������  ������      B  , ,  �,����  �,���M  �����M  ������  �,����      B  , ,  �z����  �z���M  �$���M  �$����  �z����      B  , ,  �X���K  �X����  �����  ����K  �X���K      B  , ,  �����K  ������  �P����  �P���K  �����K      B  , ,  �����K  ������  ������  �����K  �����K      B  , ,  �B���K  �B����  ������  �����K  �B���K      B  , ,  �����K  ������  �:����  �:���K  �����K      B  , ,  �����K  ������  ������  �����K  �����K      B  , ,  �,���K  �,����  ������  �����K  �,���K      B  , ,  �z���K  �z����  �$����  �$���K  �z���K      B  , ,  �6���%  �6����  ������  �����%  �6���%      B  , ,  �����%  ������  �4����  �4���%  �����%      B  , ,  �����%  ������  ������  �����%  �����%      B  , ,  �2���%  �2����  ������  �����%  �2���%      B  , ,  �����%  ������  ������  �����%  �����%      B  , ,  �����  ����ʽ  ����ʽ  �����  �����      B  , ,  �F���  �F��ʽ  ����ʽ  �����  �F���      B  , ,  �����  ����ʽ  �D��ʽ  �D���  �����      B  , ,  �����  ����ʽ  ����ʽ  �����  �����      B  , ,  �B���  �B��ʽ  ����ʽ  �����  �B���      B  , ,  �����  ����ʽ  �@��ʽ  �@���  �����      B  , ,  �����  ����ʽ  ����ʽ  �����  �����      B  , ,  �
��ş  �
���I  �����I  ����ş  �
��ş      B  , ,  �X��ş  �X���I  ����I  ���ş  �X��ş      B  , ,  �
���O  �
����  ������  �����O  �
���O      B  , ,  �X���O  �X����  �����  ����O  �X���O      B  , ,  �����O  ������  �P����  �P���O  �����O      B  , ,  �����O  ������  ������  �����O  �����O      B  , ,  �B���O  �B����  ������  �����O  �B���O      B  , ,  �����O  ������  �:����  �:���O  �����O      B  , ,  �����O  ������  ������  �����O  �����O      B  , ,  �,���O  �,����  ������  �����O  �,���O      B  , ,  �z���O  �z����  �$����  �$���O  �z���O      B  , ,  ����ş  �����I  �P���I  �P��ş  ����ş      B  , ,  ������  ����á  �0��á  �0����  ������      B  , ,  ������  ����á  �~��á  �~����  ������      B  , ,  �����  ����ʽ  ����ʽ  �����  �����      B  , ,  �.���  �.��ʽ  ����ʽ  �����  �.���      B  , ,  �����  ����ʽ  �,��ʽ  �,���  �����      B  , ,  �����  ����ʽ  ����ʽ  �����  �����      B  , ,  �*���  �*��ʽ  ����ʽ  �����  �*���      B  , ,  �~���  �~��ʽ  �(��ʽ  �(���  �~���      B  , ,  �����  ����ʽ  �|��ʽ  �|���  �����      B  , ,  �&���  �&��ʽ  ����ʽ  �����  �&���      B  , ,  �z���  �z��ʽ  �$��ʽ  �$���  �z���      B  , ,  �����  ����ʽ  �x��ʽ  �x���  �����      B  , ,  �"���  �"��ʽ  ����ʽ  �����  �"���      B  , ,  �v���  �v��ʽ  � ��ʽ  � ���  �v���      B  , ,  �����  ����ʽ  �t��ʽ  �t���  �����      B  , ,  ����K  �����  ������  �����K  ����K      B  , ,  �d���K  �d����  �����  ����K  �d���K      B  , ,  �����K  ������  �\����  �\���K  �����K      B  , ,  � ���K  � ����  ������  �����K  � ���K      B  , ,  �N���K  �N����  ������  �����K  �N���K      B  , ,  �����K  ������  �F����  �F���K  �����K      B  , ,  �����K  ������  ������  �����K  �����K      B  , ,  �8���K  �8����  ������  �����K  �8���K      B  , ,  �����K  ������  �0����  �0���K  �����K      B  , ,  �����K  ������  �~����  �~���K  �����K      B  , ,  ����  ���ʽ  ����ʽ  �����  ����      B  , ,  �r���  �r��ʽ  ���ʽ  ����  �r���      B  , ,  �����  ����ʽ  �p��ʽ  �p���  �����      B  , ,  ���ş  ����I  �����I  ����ş  ���ş      B  , ,  �d��ş  �d���I  ����I  ���ş  �d��ş      B  , ,  ����ş  �����I  �\���I  �\��ş  ����ş      B  , ,  � ��ş  � ���I  �����I  ����ş  � ��ş      B  , ,  �N��ş  �N���I  �����I  ����ş  �N��ş      B  , ,  �����  ����M  �����M  ������  �����      B  , ,  �d����  �d���M  ����M  �����  �d����      B  , ,  ������  �����M  �\���M  �\����  ������      B  , ,  � ����  � ���M  �����M  ������  � ����      B  , ,  �N����  �N���M  �����M  ������  �N����      B  , ,  ������  �����M  �F���M  �F����  ������      B  , ,  ������  �����M  �����M  ������  ������      B  , ,  �8����  �8���M  �����M  ������  �8����      B  , ,  ������  �����M  �0���M  �0����  ������      B  , ,  ������  �����M  �~���M  �~����  ������      B  , ,  ����ş  �����I  �F���I  �F��ş  ����ş      B  , ,  ����ş  �����I  �����I  ����ş  ����ş      B  , ,  �8��ş  �8���I  �����I  ����ş  �8��ş      B  , ,  ����ş  �����I  �0���I  �0��ş  ����ş      B  , ,  ����ş  �����I  �~���I  �~��ş  ����ş      B  , ,  �����%  ������  ������  �����%  �����%      B  , ,  �.���%  �.����  ������  �����%  �.���%      B  , ,  �����%  ������  �,����  �,���%  �����%      B  , ,  �����%  ������  ������  �����%  �����%      B  , ,  �*���%  �*����  ������  �����%  �*���%      B  , ,  �~���%  �~����  �(����  �(���%  �~���%      B  , ,  �����%  ������  �|����  �|���%  �����%      B  , ,  �&���%  �&����  ������  �����%  �&���%      B  , ,  �z���%  �z����  �$����  �$���%  �z���%      B  , ,  �����%  ������  �x����  �x���%  �����%      B  , ,  �"���%  �"����  ������  �����%  �"���%      B  , ,  �v���%  �v����  � ����  � ���%  �v���%      B  , ,  �����%  ������  �t����  �t���%  �����%      B  , ,  ����%  �����  ������  �����%  ����%      B  , ,  �r���%  �r����  �����  ����%  �r���%      B  , ,  �����%  ������  �p����  �p���%  �����%      B  , ,  �����%  ������  �0����  �0���%  �����%      B  , ,  �����  ����ʽ  �0��ʽ  �0���  �����      B  , ,  �����  ���á  ����á  ������  �����      B  , ,  �d����  �d��á  ���á  �����  �d����      B  , ,  ������  ����á  �\��á  �\����  ������      B  , ,  � ����  � ��á  ����á  ������  � ����      B  , ,  �N����  �N��á  ����á  ������  �N����      B  , ,  ������  ����á  �F��á  �F����  ������      B  , ,  ������  ����á  ����á  ������  ������      B  , ,  �8����  �8��á  ����á  ������  �8����      B  , ,  ����O  �����  ������  �����O  ����O      B  , ,  �d���O  �d����  �����  ����O  �d���O      B  , ,  �����O  ������  �\����  �\���O  �����O      B  , ,  � ���O  � ����  ������  �����O  � ���O      B  , ,  �N���O  �N����  ������  �����O  �N���O      B  , ,  �����O  ������  �F����  �F���O  �����O      B  , ,  �����O  ������  ������  �����O  �����O      B  , ,  �8���O  �8����  ������  �����O  �8���O      B  , ,  �����O  ������  �0����  �0���O  �����O      B  , ,  �����O  ������  �~����  �~���O  �����O      B  , ,  �"���  �"���  �����  �����  �"���      B  , ,  �p���  �p���  ����  ����  �p���      B  , ,  �����  �����  �h���  �h���  �����      B  , ,  ����  ����  �����  �����  ����      B  , ,  �Z���  �Z���  ����  ����  �Z���      B  , ,  Ũ���  Ũ���  �R���  �R���  Ũ���      B  , ,  �����  �����  Ƞ���  Ƞ���  �����      B  , ,  �D���  �D���  �����  �����  �D���      B  , ,  ̒���  ̒���  �<���  �<���  ̒���      B  , ,  �����  �����  ϊ���  ϊ���  �����      B  , ,  �.���  �.���  �����  �����  �.���      B  , ,  �h����  �h���y  ����y  �����  �h����      B  , ,  �.���U  �.����  ������  �����U  �.���U      B  , ,  �h���#  �h����  �����  ����#  �h���#      B  , ,  �V���  �V����  � ����  � ���  �V���      B  , ,  �����  ����I  Ь���I  Ь����  �����      B  , ,  �h���  �h����  �����  ����  �h���      B  , ,  �V����  �V���I  � ���I  � ����  �V����      B  , ,  �h����  �h���u  ����u  �����  �h����      B  , ,  �.���  �.���S  �����S  �����  �.���      B  , ,  �h���w  �h���!  ����!  ����w  �h���w      B  , ,  ����/  �����  Ь����  Ь���/  ����/      B  , ,  �V���/  �V����  � ����  � ���/  �V���/      B  , ,  �����  �����  Ь����  Ь����  �����      B  , ,  �V����  �V����  � ����  � ����  �V����      B  , ,  ����  �����  Ь����  Ь���  ����      B  , ,  �b����  �b���I  ����I  �����  �b����      B  , ,  ƶ����  ƶ���I  �`���I  �`����  ƶ����      B  , ,  �
����  �
���I  ȴ���I  ȴ����  �
����      B  , ,  �n����  �n����  �����  �����  �n����      B  , ,  ������  ������  �l����  �l����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �j����  �j����  �����  �����  �j����      B  , ,  ������  ������  �h����  �h����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �f����  �f����  �����  �����  �f����      B  , ,  º����  º����  �d����  �d����  º����      B  , ,  �����  �����  ĸ����  ĸ����  �����      B  , ,  �b����  �b����  �����  �����  �b����      B  , ,  ƶ����  ƶ����  �`����  �`����  ƶ����      B  , ,  �
����  �
����  ȴ����  ȴ����  �
����      B  , ,  �n���/  �n����  �����  ����/  �n���/      B  , ,  �����/  ������  �l����  �l���/  �����/      B  , ,  ����/  �����  ������  �����/  ����/      B  , ,  �j���/  �j����  �����  ����/  �j���/      B  , ,  �����/  ������  �h����  �h���/  �����/      B  , ,  ����/  �����  ������  �����/  ����/      B  , ,  �f���/  �f����  �����  ����/  �f���/      B  , ,  º���/  º����  �d����  �d���/  º���/      B  , ,  ����/  �����  ĸ����  ĸ���/  ����/      B  , ,  �b���/  �b����  �����  ����/  �b���/      B  , ,  ƶ���/  ƶ����  �`����  �`���/  ƶ���/      B  , ,  �
���/  �
����  ȴ����  ȴ���/  �
���/      B  , ,  �^���/  �^����  �����  ����/  �^���/      B  , ,  ʲ���/  ʲ����  �\����  �\���/  ʲ���/      B  , ,  ����/  �����  ̰����  ̰���/  ����/      B  , ,  �Z���/  �Z����  �����  ����/  �Z���/      B  , ,  ή���/  ή����  �X����  �X���/  ή���/      B  , ,  �"���  �"���S  �����S  �����  �"���      B  , ,  �p���  �p���S  ����S  ����  �p���      B  , ,  �����  �����S  �h���S  �h���  �����      B  , ,  ����  ����S  �����S  �����  ����      B  , ,  �����  ����I  �����I  ������  �����      B  , ,  �j����  �j���I  ����I  �����  �j����      B  , ,  �"���U  �"����  ������  �����U  �"���U      B  , ,  �p���U  �p����  �����  ����U  �p���U      B  , ,  �����U  ������  �h����  �h���U  �����U      B  , ,  ����U  �����  ������  �����U  ����U      B  , ,  �Z���U  �Z����  �����  ����U  �Z���U      B  , ,  Ũ���U  Ũ����  �R����  �R���U  Ũ���U      B  , ,  �����U  ������  Ƞ����  Ƞ���U  �����U      B  , ,  �D���U  �D����  ������  �����U  �D���U      B  , ,  ̒���U  ̒����  �<����  �<���U  ̒���U      B  , ,  �����U  ������  ϊ����  ϊ���U  �����U      B  , ,  �Z���  �Z���S  ����S  ����  �Z���      B  , ,  Ũ���  Ũ���S  �R���S  �R���  Ũ���      B  , ,  �����  �����S  Ƞ���S  Ƞ���  �����      B  , ,  �D���  �D���S  �����S  �����  �D���      B  , ,  ̒���  ̒���S  �<���S  �<���  ̒���      B  , ,  �����  �����S  ϊ���S  ϊ���  �����      B  , ,  �n����  �n���I  ����I  �����  �n����      B  , ,  ������  �����I  �l���I  �l����  ������      B  , ,  ������  �����I  �h���I  �h����  ������      B  , ,  �����  ����I  �����I  ������  �����      B  , ,  �^����  �^����  �����  �����  �^����      B  , ,  ʲ����  ʲ����  �\����  �\����  ʲ����      B  , ,  �����  �����  ̰����  ̰����  �����      B  , ,  �Z����  �Z����  �����  �����  �Z����      B  , ,  ή����  ή����  �X����  �X����  ή����      B  , ,  �f����  �f���I  ����I  �����  �f����      B  , ,  º����  º���I  �d���I  �d����  º����      B  , ,  �^����  �^���I  ����I  �����  �^����      B  , ,  ʲ����  ʲ���I  �\���I  �\����  ʲ����      B  , ,  �����  ����I  ̰���I  ̰����  �����      B  , ,  �Z����  �Z���I  ����I  �����  �Z����      B  , ,  ή����  ή���I  �X���I  �X����  ή����      B  , ,  �n���  �n����  �����  ����  �n���      B  , ,  �����  ������  �l����  �l���  �����      B  , ,  ����  �����  ������  �����  ����      B  , ,  �j���  �j����  �����  ����  �j���      B  , ,  �����  ������  �h����  �h���  �����      B  , ,  ����  �����  ������  �����  ����      B  , ,  �f���  �f����  �����  ����  �f���      B  , ,  º���  º����  �d����  �d���  º���      B  , ,  ����  �����  ĸ����  ĸ���  ����      B  , ,  �b���  �b����  �����  ����  �b���      B  , ,  ƶ���  ƶ����  �`����  �`���  ƶ���      B  , ,  �
���  �
����  ȴ����  ȴ���  �
���      B  , ,  �^���  �^����  �����  ����  �^���      B  , ,  ʲ���  ʲ����  �\����  �\���  ʲ���      B  , ,  ����  �����  ̰����  ̰���  ����      B  , ,  �Z���  �Z����  �����  ����  �Z���      B  , ,  ή���  ή����  �X����  �X���  ή���      B  , ,  �����  ����I  ĸ���I  ĸ����  �����      B  , ,  ����  ����W  �����W  �����  ����      B  , ,  �Z���  �Z���W  ����W  ����  �Z���      B  , ,  Ũ���  Ũ���W  �R���W  �R���  Ũ���      B  , ,  �����  �����W  Ƞ���W  Ƞ���  �����      B  , ,  ������  �����  �����  ������  ������      B  , ,  �I����  �I���  �����  ������  �I����      B  , ,  ������  �����  �A���  �A����  ������      B  , ,  ������  �����  �����  ������  ������      B  , ,  �3����  �3���  �����  ������  �3����      B  , ,  ā����  ā���  �+���  �+����  ā����      B  , ,  ������  �����  �y���  �y����  ������      B  , ,  �����  ����  �����  ������  �����      B  , ,  �k����  �k���  ����  �����  �k����      B  , ,  ͹����  ͹���  �c���  �c����  ͹����      B  , ,  �D���  �D���W  �����W  �����  �D���      B  , ,  �"���]  �"���  �����  �����]  �"���]      B  , ,  �p���]  �p���  ����  ����]  �p���]      B  , ,  �����]  �����  �h���  �h���]  �����]      B  , ,  ����]  ����  �����  �����]  ����]      B  , ,  �Z���]  �Z���  ����  ����]  �Z���]      B  , ,  Ũ���]  Ũ���  �R���  �R���]  Ũ���]      B  , ,  �����]  �����  Ƞ���  Ƞ���]  �����]      B  , ,  �D���]  �D���  �����  �����]  �D���]      B  , ,  ̒���]  ̒���  �<���  �<���]  ̒���]      B  , ,  �����]  �����  ϊ���  ϊ���]  �����]      B  , ,  ̒���  ̒���W  �<���W  �<���  ̒���      B  , ,  �"���  �"���[  �����[  �����  �"���      B  , ,  �p���  �p���[  ����[  ����  �p���      B  , ,  �"���Y  �"���  �����  �����Y  �"���Y      B  , ,  �"���  �"���  �����  �����  �"���      B  , ,  �p���  �p���  ����  ����  �p���      B  , ,  �����  �����  �h���  �h���  �����      B  , ,  ����  ����  �����  �����  ����      B  , ,  �Z���  �Z���  ����  ����  �Z���      B  , ,  Ũ���  Ũ���  �R���  �R���  Ũ���      B  , ,  �����  �����  Ƞ���  Ƞ���  �����      B  , ,  �D���  �D���  �����  �����  �D���      B  , ,  ̒���  ̒���  �<���  �<���  ̒���      B  , ,  �����  �����  ϊ���  ϊ���  �����      B  , ,  �p���Y  �p���  ����  ����Y  �p���Y      B  , ,  �����Y  �����  �h���  �h���Y  �����Y      B  , ,  ����Y  ����  �����  �����Y  ����Y      B  , ,  �Z���Y  �Z���  ����  ����Y  �Z���Y      B  , ,  Ũ���Y  Ũ���  �R���  �R���Y  Ũ���Y      B  , ,  �����Y  �����  Ƞ���  Ƞ���Y  �����Y      B  , ,  �D���Y  �D���  �����  �����Y  �D���Y      B  , ,  ̒���Y  ̒���  �<���  �<���Y  ̒���Y      B  , ,  �����Y  �����  ϊ���  ϊ���Y  �����Y      B  , ,  �����  �����[  �h���[  �h���  �����      B  , ,  ����  ����[  �����[  �����  ����      B  , ,  �Z���  �Z���[  ����[  ����  �Z���      B  , ,  Ũ���  Ũ���[  �R���[  �R���  Ũ���      B  , ,  ������  �����u  �����u  ������  ������      B  , ,  �I����  �I���u  �����u  ������  �I����      B  , ,  ������  �����u  �A���u  �A����  ������      B  , ,  ������  �����u  �����u  ������  ������      B  , ,  �3����  �3���u  �����u  ������  �3����      B  , ,  ā����  ā���u  �+���u  �+����  ā����      B  , ,  ������  �����u  �y���u  �y����  ������      B  , ,  �����  ����u  �����u  ������  �����      B  , ,  �k����  �k���u  ����u  �����  �k����      B  , ,  ͹����  ͹���u  �c���u  �c����  ͹����      B  , ,  �����  �����[  Ƞ���[  Ƞ���  �����      B  , ,  �D���  �D���[  �����[  �����  �D���      B  , ,  ̒���  ̒���[  �<���[  �<���  ̒���      B  , ,  �����  �����[  ϊ���[  ϊ���  �����      B  , ,  �����  �����W  ϊ���W  ϊ���  �����      B  , ,  �"���U  �"����  ������  �����U  �"���U      B  , ,  �p���U  �p����  �����  ����U  �p���U      B  , ,  �����U  ������  �h����  �h���U  �����U      B  , ,  ����U  �����  ������  �����U  ����U      B  , ,  �Z���U  �Z����  �����  ����U  �Z���U      B  , ,  Ũ���U  Ũ����  �R����  �R���U  Ũ���U      B  , ,  �����U  ������  Ƞ����  Ƞ���U  �����U      B  , ,  �D���U  �D����  ������  �����U  �D���U      B  , ,  ̒���U  ̒����  �<����  �<���U  ̒���U      B  , ,  �����U  ������  ϊ����  ϊ���U  �����U      B  , ,  �"���  �"���W  �����W  �����  �"���      B  , ,  �p���  �p���W  ����W  ����  �p���      B  , ,  �����  �����W  �h���W  �h���  �����      B  , ,  �h����  �h��߅  ���߅  �����  �h����      B  , ,  �h��݇  �h���1  ����1  ���݇  �h��݇      B  , ,  �h���{  �h���%  ����%  ����{  �h���{      B  , ,  �.���]  �.���  �����  �����]  �.���]      B  , ,  �����  ����  б���  б����  �����      B  , ,  �.���  �.���  �����  �����  �.���      B  , ,  �h����  �h���}  ����}  �����  �h����      B  , ,  �h���  �h���-  ����-  ����  �h���      B  , ,  �h���+  �h����  �����  ����+  �h���+      B  , ,  �.���  �.���[  �����[  �����  �.���      B  , ,  �h����  �h���  ����  �����  �h����      B  , ,  �.���  �.���W  �����W  �����  �.���      B  , ,  �h���  �h���)  ����)  ����  �h���      B  , ,  �.���U  �.����  ������  �����U  �.���U      B  , ,  �.���Y  �.���  �����  �����Y  �.���Y      B  , ,  �����  ����u  б���u  б����  �����      B  , ,  �h���/  �h����  �����  ����/  �h���/      B  , ,  �h���'  �h����  �����  ����'  �h���'      B  , ,  �n����  �n��·  ���·  �����  �n����      B  , ,  ������  ����·  �l��·  �l����  ������      B  , ,  �����  ���·  ����·  ������  �����      B  , ,  �j����  �j��·  ���·  �����  �j����      B  , ,  ������  ����·  �h��·  �h����  ������      B  , ,  �����  ���·  ����·  ������  �����      B  , ,  �f����  �f��·  ���·  �����  �f����      B  , ,  º����  º��·  �d��·  �d����  º����      B  , ,  �����  ���·  ĸ��·  ĸ����  �����      B  , ,  �b����  �b��·  ���·  �����  �b����      B  , ,  ƶ����  ƶ��·  �`��·  �`����  ƶ����      B  , ,  �
����  �
��·  ȴ��·  ȴ����  �
����      B  , ,  �^����  �^��·  ���·  �����  �^����      B  , ,  ʲ����  ʲ��·  �\��·  �\����  ʲ����      B  , ,  �����  ���·  ̰��·  ̰����  �����      B  , ,  �Z����  �Z��·  ���·  �����  �Z����      B  , ,  ή����  ή��·  �X��·  �X����  ή����      B  , ,  �����  ���·  Ь��·  Ь����  �����      B  , ,  �V����  �V��·  � ��·  � ����  �V����      B  , ,  �h����  �h��ۉ  ���ۉ  �����  �h����      B  , ,  �.���  �.��ܫ  ����ܫ  �����  �.���      B  , ,  �h���3  �h����  �����  ����3  �h���3      B  , ,  �.��ֱ  �.���[  �����[  ����ֱ  �.��ֱ      B  , ,  �h����  �h��׍  ���׍  �����  �h����      B  , ,  ���ϕ  ����?  Ь���?  Ь��ϕ  ���ϕ      B  , ,  �V��ϕ  �V���?  � ���?  � ��ϕ  �V��ϕ      B  , ,  �.���Y  �.���  �����  �����Y  �.���Y      B  , ,  �h��ً  �h���5  ����5  ���ً  �h��ً      B  , ,  �.���	  �.��Գ  ����Գ  �����	  �.���	      B  , ,  �h���;  �h����  �����  ����;  �h���;      B  , ,  �h����  �h��ӑ  ���ӑ  �����  �h����      B  , ,  �h��ѓ  �h���=  ����=  ���ѓ  �h��ѓ      B  , ,  �.���  �.��د  ����د  �����  �.���      B  , ,  �h���7  �h����  �����  ����7  �h���7      B  , ,  �.���]  �.���  �����  �����]  �.���]      B  , ,  �h��Տ  �h���9  ����9  ���Տ  �h��Տ      B  , ,  �.��ڭ  �.���W  �����W  ����ڭ  �.��ڭ      B  , ,  ���ϕ  ����?  �����?  ����ϕ  ���ϕ      B  , ,  �f��ϕ  �f���?  ����?  ���ϕ  �f��ϕ      B  , ,  º��ϕ  º���?  �d���?  �d��ϕ  º��ϕ      B  , ,  ���ϕ  ����?  ĸ���?  ĸ��ϕ  ���ϕ      B  , ,  �b��ϕ  �b���?  ����?  ���ϕ  �b��ϕ      B  , ,  ƶ��ϕ  ƶ���?  �`���?  �`��ϕ  ƶ��ϕ      B  , ,  �
��ϕ  �
���?  ȴ���?  ȴ��ϕ  �
��ϕ      B  , ,  �^��ϕ  �^���?  ����?  ���ϕ  �^��ϕ      B  , ,  ʲ��ϕ  ʲ���?  �\���?  �\��ϕ  ʲ��ϕ      B  , ,  ���ϕ  ����?  ̰���?  ̰��ϕ  ���ϕ      B  , ,  �Z��ϕ  �Z���?  ����?  ���ϕ  �Z��ϕ      B  , ,  ή��ϕ  ή���?  �X���?  �X��ϕ  ή��ϕ      B  , ,  �Z��ڭ  �Z���W  ����W  ���ڭ  �Z��ڭ      B  , ,  Ũ��ڭ  Ũ���W  �R���W  �R��ڭ  Ũ��ڭ      B  , ,  �"���Y  �"���  �����  �����Y  �"���Y      B  , ,  �p���Y  �p���  ����  ����Y  �p���Y      B  , ,  �����Y  �����  �h���  �h���Y  �����Y      B  , ,  ����Y  ����  �����  �����Y  ����Y      B  , ,  �Z���Y  �Z���  ����  ����Y  �Z���Y      B  , ,  Ũ���Y  Ũ���  �R���  �R���Y  Ũ���Y      B  , ,  �����Y  �����  Ƞ���  Ƞ���Y  �����Y      B  , ,  �D���Y  �D���  �����  �����Y  �D���Y      B  , ,  ̒���Y  ̒���  �<���  �<���Y  ̒���Y      B  , ,  �����Y  �����  ϊ���  ϊ���Y  �����Y      B  , ,  �"���  �"��ܫ  ����ܫ  �����  �"���      B  , ,  �p���  �p��ܫ  ���ܫ  ����  �p���      B  , ,  �"���	  �"��Գ  ����Գ  �����	  �"���	      B  , ,  �p���	  �p��Գ  ���Գ  ����	  �p���	      B  , ,  �����	  ����Գ  �h��Գ  �h���	  �����	      B  , ,  ����	  ���Գ  ����Գ  �����	  ����	      B  , ,  �Z���	  �Z��Գ  ���Գ  ����	  �Z���	      B  , ,  Ũ���	  Ũ��Գ  �R��Գ  �R���	  Ũ���	      B  , ,  �����	  ����Գ  Ƞ��Գ  Ƞ���	  �����	      B  , ,  �D���	  �D��Գ  ����Գ  �����	  �D���	      B  , ,  ̒���	  ̒��Գ  �<��Գ  �<���	  ̒���	      B  , ,  �����	  ����Գ  ϊ��Գ  ϊ���	  �����	      B  , ,  �����  ����ܫ  �h��ܫ  �h���  �����      B  , ,  ����  ���ܫ  ����ܫ  �����  ����      B  , ,  �Z���  �Z��ܫ  ���ܫ  ����  �Z���      B  , ,  Ũ���  Ũ��ܫ  �R��ܫ  �R���  Ũ���      B  , ,  �"���]  �"���  �����  �����]  �"���]      B  , ,  �p���]  �p���  ����  ����]  �p���]      B  , ,  �����]  �����  �h���  �h���]  �����]      B  , ,  ����]  ����  �����  �����]  ����]      B  , ,  �Z���]  �Z���  ����  ����]  �Z���]      B  , ,  Ũ���]  Ũ���  �R���  �R���]  Ũ���]      B  , ,  �����]  �����  Ƞ���  Ƞ���]  �����]      B  , ,  �D���]  �D���  �����  �����]  �D���]      B  , ,  ̒���]  ̒���  �<���  �<���]  ̒���]      B  , ,  �"���  �"��د  ����د  �����  �"���      B  , ,  �p���  �p��د  ���د  ����  �p���      B  , ,  �����  ����د  �h��د  �h���  �����      B  , ,  ����  ���د  ����د  �����  ����      B  , ,  �Z���  �Z��د  ���د  ����  �Z���      B  , ,  Ũ���  Ũ��د  �R��د  �R���  Ũ���      B  , ,  �����  ����د  Ƞ��د  Ƞ���  �����      B  , ,  �D���  �D��د  ����د  �����  �D���      B  , ,  ̒���  ̒��د  �<��د  �<���  ̒���      B  , ,  �����  ����د  ϊ��د  ϊ���  �����      B  , ,  �����  ����ܫ  Ƞ��ܫ  Ƞ���  �����      B  , ,  �D���  �D��ܫ  ����ܫ  �����  �D���      B  , ,  �����]  �����  ϊ���  ϊ���]  �����]      B  , ,  ̒���  ̒��ܫ  �<��ܫ  �<���  ̒���      B  , ,  �����  ����ܫ  ϊ��ܫ  ϊ���  �����      B  , ,  ����ڭ  �����W  Ƞ���W  Ƞ��ڭ  ����ڭ      B  , ,  �D��ڭ  �D���W  �����W  ����ڭ  �D��ڭ      B  , ,  �D��ֱ  �D���[  �����[  ����ֱ  �D��ֱ      B  , ,  ̒��ֱ  ̒���[  �<���[  �<��ֱ  ̒��ֱ      B  , ,  ����ֱ  �����[  ϊ���[  ϊ��ֱ  ����ֱ      B  , ,  ̒��ڭ  ̒���W  �<���W  �<��ڭ  ̒��ڭ      B  , ,  ����ڭ  �����W  ϊ���W  ϊ��ڭ  ����ڭ      B  , ,  �"��ֱ  �"���[  �����[  ����ֱ  �"��ֱ      B  , ,  �p��ֱ  �p���[  ����[  ���ֱ  �p��ֱ      B  , ,  ����ֱ  �����[  �h���[  �h��ֱ  ����ֱ      B  , ,  ���ֱ  ����[  �����[  ����ֱ  ���ֱ      B  , ,  �Z��ֱ  �Z���[  ����[  ���ֱ  �Z��ֱ      B  , ,  Ũ��ֱ  Ũ���[  �R���[  �R��ֱ  Ũ��ֱ      B  , ,  ����ֱ  �����[  Ƞ���[  Ƞ��ֱ  ����ֱ      B  , ,  �n��ϕ  �n���?  ����?  ���ϕ  �n��ϕ      B  , ,  ����ϕ  �����?  �l���?  �l��ϕ  ����ϕ      B  , ,  ���ϕ  ����?  �����?  ����ϕ  ���ϕ      B  , ,  �j��ϕ  �j���?  ����?  ���ϕ  �j��ϕ      B  , ,  ����ϕ  �����?  �h���?  �h��ϕ  ����ϕ      B  , ,  �"��ڭ  �"���W  �����W  ����ڭ  �"��ڭ      B  , ,  �p��ڭ  �p���W  ����W  ���ڭ  �p��ڭ      B  , ,  ����ڭ  �����W  �h���W  �h��ڭ  ����ڭ      B  , ,  ���ڭ  ����W  �����W  ����ڭ  ���ڭ      B  , ,  ����ş  �����I  ϊ���I  ϊ��ş  ����ş      B  , ,  �"��ş  �"���I  �����I  ����ş  �"��ş      B  , ,  �p��ş  �p���I  ����I  ���ş  �p��ş      B  , ,  ����ş  �����I  �h���I  �h��ş  ����ş      B  , ,  ���ş  ����I  �����I  ����ş  ���ş      B  , ,  �Z��ş  �Z���I  ����I  ���ş  �Z��ş      B  , ,  Ũ��ş  Ũ���I  �R���I  �R��ş  Ũ��ş      B  , ,  ����ş  �����I  Ƞ���I  Ƞ��ş  ����ş      B  , ,  ����%  �����  ĸ����  ĸ���%  ����%      B  , ,  �D��ş  �D���I  �����I  ����ş  �D��ş      B  , ,  �b���%  �b����  �����  ����%  �b���%      B  , ,  �Z���%  �Z����  �����  ����%  �Z���%      B  , ,  ή���%  ή����  �X����  �X���%  ή���%      B  , ,  �n���%  �n����  �����  ����%  �n���%      B  , ,  �����%  ������  �l����  �l���%  �����%      B  , ,  �n���  �n��ʽ  ���ʽ  ����  �n���      B  , ,  �����  ����ʽ  �l��ʽ  �l���  �����      B  , ,  ����  ���ʽ  ����ʽ  �����  ����      B  , ,  �"���K  �"����  ������  �����K  �"���K      B  , ,  �p���K  �p����  �����  ����K  �p���K      B  , ,  ƶ���  ƶ��ʽ  �`��ʽ  �`���  ƶ���      B  , ,  �����K  ������  �h����  �h���K  �����K      B  , ,  ����K  �����  ������  �����K  ����K      B  , ,  �"����  �"���M  �����M  ������  �"����      B  , ,  �p����  �p���M  ����M  �����  �p����      B  , ,  ������  �����M  �h���M  �h����  ������      B  , ,  �����  ����M  �����M  ������  �����      B  , ,  �Z����  �Z���M  ����M  �����  �Z����      B  , ,  Ũ����  Ũ���M  �R���M  �R����  Ũ����      B  , ,  ������  �����M  Ƞ���M  Ƞ����  ������      B  , ,  �D����  �D���M  �����M  ������  �D����      B  , ,  ̒����  ̒���M  �<���M  �<����  ̒����      B  , ,  ������  �����M  ϊ���M  ϊ����  ������      B  , ,  �Z���K  �Z����  �����  ����K  �Z���K      B  , ,  Ũ���K  Ũ����  �R����  �R���K  Ũ���K      B  , ,  �����K  ������  Ƞ����  Ƞ���K  �����K      B  , ,  �D���K  �D����  ������  �����K  �D���K      B  , ,  ̒���K  ̒����  �<����  �<���K  ̒���K      B  , ,  �����K  ������  ϊ����  ϊ���K  �����K      B  , ,  �j���  �j��ʽ  ���ʽ  ����  �j���      B  , ,  �����  ����ʽ  �h��ʽ  �h���  �����      B  , ,  ����  ���ʽ  ����ʽ  �����  ����      B  , ,  �f���  �f��ʽ  ���ʽ  ����  �f���      B  , ,  �
���  �
��ʽ  ȴ��ʽ  ȴ���  �
���      B  , ,  �^���  �^��ʽ  ���ʽ  ����  �^���      B  , ,  �"����  �"��á  ����á  ������  �"����      B  , ,  �p����  �p��á  ���á  �����  �p����      B  , ,  ������  ����á  �h��á  �h����  ������      B  , ,  �����  ���á  ����á  ������  �����      B  , ,  �Z����  �Z��á  ���á  �����  �Z����      B  , ,  Ũ����  Ũ��á  �R��á  �R����  Ũ����      B  , ,  ������  ����á  Ƞ��á  Ƞ����  ������      B  , ,  �D����  �D��á  ����á  ������  �D����      B  , ,  ̒����  ̒��á  �<��á  �<����  ̒����      B  , ,  ������  ����á  ϊ��á  ϊ����  ������      B  , ,  ʲ���  ʲ��ʽ  �\��ʽ  �\���  ʲ���      B  , ,  ����  ���ʽ  ̰��ʽ  ̰���  ����      B  , ,  �Z���  �Z��ʽ  ���ʽ  ����  �Z���      B  , ,  ή���  ή��ʽ  �X��ʽ  �X���  ή���      B  , ,  ����%  �����  ������  �����%  ����%      B  , ,  �j���%  �j����  �����  ����%  �j���%      B  , ,  �����%  ������  �h����  �h���%  �����%      B  , ,  ����%  �����  ������  �����%  ����%      B  , ,  �f���%  �f����  �����  ����%  �f���%      B  , ,  º���%  º����  �d����  �d���%  º���%      B  , ,  ƶ���%  ƶ����  �`����  �`���%  ƶ���%      B  , ,  �
���%  �
����  ȴ����  ȴ���%  �
���%      B  , ,  �^���%  �^����  �����  ����%  �^���%      B  , ,  ʲ���%  ʲ����  �\����  �\���%  ʲ���%      B  , ,  ����%  �����  ̰����  ̰���%  ����%      B  , ,  º���  º��ʽ  �d��ʽ  �d���  º���      B  , ,  ����  ���ʽ  ĸ��ʽ  ĸ���  ����      B  , ,  �b���  �b��ʽ  ���ʽ  ����  �b���      B  , ,  ̒��ş  ̒���I  �<���I  �<��ş  ̒��ş      B  , ,  �"���O  �"����  ������  �����O  �"���O      B  , ,  �p���O  �p����  �����  ����O  �p���O      B  , ,  �����O  ������  �h����  �h���O  �����O      B  , ,  ����O  �����  ������  �����O  ����O      B  , ,  �Z���O  �Z����  �����  ����O  �Z���O      B  , ,  Ũ���O  Ũ����  �R����  �R���O  Ũ���O      B  , ,  �����O  ������  Ƞ����  Ƞ���O  �����O      B  , ,  �D���O  �D����  ������  �����O  �D���O      B  , ,  ̒���O  ̒����  �<����  �<���O  ̒���O      B  , ,  �����O  ������  ϊ����  ϊ���O  �����O      B  , ,  ����%  �����  Ь����  Ь���%  ����%      B  , ,  �.���K  �.����  ������  �����K  �.���K      B  , ,  �h���  �h����  �����  ����  �h���      B  , ,  �.����  �.���M  �����M  ������  �.����      B  , ,  �h���q  �h���  ����  ����q  �h���q      B  , ,  �V���%  �V����  � ����  � ���%  �V���%      B  , ,  ����  ���ʽ  Ь��ʽ  Ь���  ����      B  , ,  �V���  �V��ʽ  � ��ʽ  � ���  �V���      B  , ,  �.��ş  �.���I  �����I  ����ş  �.��ş      B  , ,  �h���  �h��ȿ  ���ȿ  ����  �h���      B  , ,  �h���m  �h���  ����  ����m  �h���m      B  , ,  �h����  �h���k  ����k  �����  �h����      B  , ,  �.����  �.��á  ����á  ������  �.����      B  , ,  �h����  �h���o  ����o  �����  �h����      B  , ,  �.���O  �.����  ������  �����O  �.���O      B  , ,  �h���  �h����  �����  ����  �h���      B  , ,  �����  ����5  �����5  ������  �����      B  , ,  �����  ����}  �����}  ������  �����      B  , ,  ����  �����  ������  �����  ����      B  , ,  ���}�  ���~s  ����~s  ����}�  ���}�      B  , ,  ���|  ���|�  ����|�  ����|  ���|      B  , ,  �"���O  �"����  ������  �����O  �"���O      B  , ,  �p���O  �p����  �����  ����O  �p���O      B  , ,  �����O  ������  �h����  �h���O  �����O      B  , ,  ����O  �����  ������  �����O  ����O      B  , ,  �Z���O  �Z����  �����  ����O  �Z���O      B  , ,  Ũ���O  Ũ����  �R����  �R���O  Ũ���O      B  , ,  �����O  ������  Ƞ����  Ƞ���O  �����O      B  , ,  �D���O  �D����  ������  �����O  �D���O      B  , ,  ̒���O  ̒����  �<����  �<���O  ̒���O      B  , ,  �����O  ������  ϊ����  ϊ���O  �����O      B  , ,  �.���O  �.����  ������  �����O  �.���O      B  , ,  �h����  �h���+  ����+  �����  �h����      B  , ,  �.���K  �.����  ������  �����K  �.���K      B  , ,  �h���}  �h���'  ����'  ����}  �h���}      B  , ,  �.����  �.����  ������  ������  �.����      B  , ,  �h���)  �h����  �����  ����)  �h���)      B  , ,  �.����  �.���M  �����M  ������  �.����      B  , ,  �h����  �h���  ����  �����  �h����      B  , ,  �.����  �.����  ������  ������  �.����      B  , ,  �h����  �h���s  ����s  �����  �h����      B  , ,  �.����  �.���Q  �����Q  ������  �.����      B  , ,  �h���u  �h���  ����  ����u  �h���u      B  , ,  �.���S  �.����  ������  �����S  �.���S      B  , ,  �h���!  �h����  �����  ����!  �h���!      B  , ,  �h����  �h���w  ����w  �����  �h����      B  , ,  �����  �����  б����  б����  �����      B  , ,  �h���y  �h���#  ����#  ����y  �h���y      B  , ,  �����  ����k  б���k  б����  �����      B  , ,  �h���%  �h����  �����  ����%  �h���%      B  , ,  �h����  �h���{  ����{  �����  �h����      B  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      B  , ,  ������  ������  Ƞ����  Ƞ����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �I����  �I����  ������  ������  �I����      B  , ,  ������  ������  �A����  �A����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �3����  �3����  ������  ������  �3����      B  , ,  ā����  ā����  �+����  �+����  ā����      B  , ,  ������  ������  �y����  �y����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �k����  �k����  �����  �����  �k����      B  , ,  ͹����  ͹����  �c����  �c����  ͹����      B  , ,  �"����  �"���Q  �����Q  ������  �"����      B  , ,  �p����  �p���Q  ����Q  �����  �p����      B  , ,  ������  �����k  �����k  ������  ������      B  , ,  �I����  �I���k  �����k  ������  �I����      B  , ,  ������  �����k  �A���k  �A����  ������      B  , ,  ������  �����k  �����k  ������  ������      B  , ,  �3����  �3���k  �����k  ������  �3����      B  , ,  ā����  ā���k  �+���k  �+����  ā����      B  , ,  ������  �����k  �y���k  �y����  ������      B  , ,  �����  ����k  �����k  ������  �����      B  , ,  �k����  �k���k  ����k  �����  �k����      B  , ,  ͹����  ͹���k  �c���k  �c����  ͹����      B  , ,  ������  �����Q  �h���Q  �h����  ������      B  , ,  �����  ����Q  �����Q  ������  �����      B  , ,  �Z����  �Z���Q  ����Q  �����  �Z����      B  , ,  �"���K  �"����  ������  �����K  �"���K      B  , ,  �p���K  �p����  �����  ����K  �p���K      B  , ,  �����K  ������  �h����  �h���K  �����K      B  , ,  ����K  �����  ������  �����K  ����K      B  , ,  �Z���K  �Z����  �����  ����K  �Z���K      B  , ,  Ũ���K  Ũ����  �R����  �R���K  Ũ���K      B  , ,  �����K  ������  Ƞ����  Ƞ���K  �����K      B  , ,  �D���K  �D����  ������  �����K  �D���K      B  , ,  ̒���K  ̒����  �<����  �<���K  ̒���K      B  , ,  �����K  ������  ϊ����  ϊ���K  �����K      B  , ,  Ũ����  Ũ���Q  �R���Q  �R����  Ũ����      B  , ,  ������  �����Q  Ƞ���Q  Ƞ����  ������      B  , ,  �"����  �"����  ������  ������  �"����      B  , ,  �p����  �p����  �����  �����  �p����      B  , ,  ������  ������  �h����  �h����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �Z����  �Z����  �����  �����  �Z����      B  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      B  , ,  ������  ������  Ƞ����  Ƞ����  ������      B  , ,  �D����  �D����  ������  ������  �D����      B  , ,  ̒����  ̒����  �<����  �<����  ̒����      B  , ,  ������  ������  ϊ����  ϊ����  ������      B  , ,  �D����  �D���Q  �����Q  ������  �D����      B  , ,  ̒����  ̒���Q  �<���Q  �<����  ̒����      B  , ,  �"����  �"���M  �����M  ������  �"����      B  , ,  �p����  �p���M  ����M  �����  �p����      B  , ,  ������  �����M  �h���M  �h����  ������      B  , ,  �����  ����M  �����M  ������  �����      B  , ,  �Z����  �Z���M  ����M  �����  �Z����      B  , ,  Ũ����  Ũ���M  �R���M  �R����  Ũ����      B  , ,  ������  �����M  Ƞ���M  Ƞ����  ������      B  , ,  �D����  �D���M  �����M  ������  �D����      B  , ,  ̒����  ̒���M  �<���M  �<����  ̒����      B  , ,  ������  �����M  ϊ���M  ϊ����  ������      B  , ,  ������  �����Q  ϊ���Q  ϊ����  ������      B  , ,  �D����  �D����  ������  ������  �D����      B  , ,  ̒����  ̒����  �<����  �<����  ̒����      B  , ,  �"���S  �"����  ������  �����S  �"���S      B  , ,  �p���S  �p����  �����  ����S  �p���S      B  , ,  �����S  ������  �h����  �h���S  �����S      B  , ,  ����S  �����  ������  �����S  ����S      B  , ,  �Z���S  �Z����  �����  ����S  �Z���S      B  , ,  Ũ���S  Ũ����  �R����  �R���S  Ũ���S      B  , ,  �����S  ������  Ƞ����  Ƞ���S  �����S      B  , ,  �D���S  �D����  ������  �����S  �D���S      B  , ,  ̒���S  ̒����  �<����  �<���S  ̒���S      B  , ,  �����S  ������  ϊ����  ϊ���S  �����S      B  , ,  ������  ������  ϊ����  ϊ����  ������      B  , ,  �"����  �"����  ������  ������  �"����      B  , ,  �p����  �p����  �����  �����  �p����      B  , ,  ������  ������  �h����  �h����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �Z����  �Z����  �����  �����  �Z����      B  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      B  , ,  ������  ������  Ƞ����  Ƞ����  ������      B  , ,  �D����  �D����  ������  ������  �D����      B  , ,  ̒����  ̒����  �<����  �<����  ̒����      B  , ,  ������  ������  ϊ����  ϊ����  ������      B  , ,  �"����  �"���Q  �����Q  ������  �"����      B  , ,  �p����  �p���Q  ����Q  �����  �p����      B  , ,  ������  �����Q  �h���Q  �h����  ������      B  , ,  �����  ����Q  �����Q  ������  �����      B  , ,  �Z����  �Z���Q  ����Q  �����  �Z����      B  , ,  Ũ����  Ũ���Q  �R���Q  �R����  Ũ����      B  , ,  ������  �����Q  Ƞ���Q  Ƞ����  ������      B  , ,  �D����  �D���Q  �����Q  ������  �D����      B  , ,  ̒����  ̒���Q  �<���Q  �<����  ̒����      B  , ,  ������  �����Q  ϊ���Q  ϊ����  ������      B  , ,  �"���S  �"����  ������  �����S  �"���S      B  , ,  �p���S  �p����  �����  ����S  �p���S      B  , ,  �����S  ������  �h����  �h���S  �����S      B  , ,  ����S  �����  ������  �����S  ����S      B  , ,  �Z���S  �Z����  �����  ����S  �Z���S      B  , ,  Ũ���S  Ũ����  �R����  �R���S  Ũ���S      B  , ,  �����S  ������  Ƞ����  Ƞ���S  �����S      B  , ,  �D���S  �D����  ������  �����S  �D���S      B  , ,  ̒���S  ̒����  �<����  �<���S  ̒���S      B  , ,  �����S  ������  ϊ����  ϊ���S  �����S      B  , ,  �"����  �"����  ������  ������  �"����      B  , ,  �p����  �p����  �����  �����  �p����      B  , ,  ������  ������  �h����  �h����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �Z����  �Z����  �����  �����  �Z����      B  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      B  , ,  ������  ������  Ƞ����  Ƞ����  ������      B  , ,  �D����  �D����  ������  ������  �D����      B  , ,  ̒����  ̒����  �<����  �<����  ̒����      B  , ,  ������  ������  ϊ����  ϊ����  ������      B  , ,  �"����  �"����  ������  ������  �"����      B  , ,  �n����  �n���5  ����5  �����  �n����      B  , ,  ������  �����5  �l���5  �l����  ������      B  , ,  �����  ����5  �����5  ������  �����      B  , ,  �j����  �j���5  ����5  �����  �j����      B  , ,  ������  �����5  �h���5  �h����  ������      B  , ,  �����  ����5  �����5  ������  �����      B  , ,  �f����  �f���5  ����5  �����  �f����      B  , ,  º����  º���5  �d���5  �d����  º����      B  , ,  �����  ����5  ĸ���5  ĸ����  �����      B  , ,  �b����  �b���5  ����5  �����  �b����      B  , ,  ƶ����  ƶ���5  �`���5  �`����  ƶ����      B  , ,  �
����  �
���5  ȴ���5  ȴ����  �
����      B  , ,  �^����  �^���5  ����5  �����  �^����      B  , ,  ʲ����  ʲ���5  �\���5  �\����  ʲ����      B  , ,  �����  ����5  ̰���5  ̰����  �����      B  , ,  �Z����  �Z���5  ����5  �����  �Z����      B  , ,  ή����  ή���5  �X���5  �X����  ή����      B  , ,  �p����  �p����  �����  �����  �p����      B  , ,  �n����  �n���}  ����}  �����  �n����      B  , ,  ������  �����}  �l���}  �l����  ������      B  , ,  �����  ����}  �����}  ������  �����      B  , ,  �j����  �j���}  ����}  �����  �j����      B  , ,  ������  �����}  �h���}  �h����  ������      B  , ,  �����  ����}  �����}  ������  �����      B  , ,  �f����  �f���}  ����}  �����  �f����      B  , ,  º����  º���}  �d���}  �d����  º����      B  , ,  �����  ����}  ĸ���}  ĸ����  �����      B  , ,  �b����  �b���}  ����}  �����  �b����      B  , ,  ƶ����  ƶ���}  �`���}  �`����  ƶ����      B  , ,  �
����  �
���}  ȴ���}  ȴ����  �
����      B  , ,  �^����  �^���}  ����}  �����  �^����      B  , ,  ʲ����  ʲ���}  �\���}  �\����  ʲ����      B  , ,  �����  ����}  ̰���}  ̰����  �����      B  , ,  �Z����  �Z���}  ����}  �����  �Z����      B  , ,  ή����  ή���}  �X���}  �X����  ή����      B  , ,  ������  ������  �h����  �h����  ������      B  , ,  �n���  �n����  �����  ����  �n���      B  , ,  �����  ������  �l����  �l���  �����      B  , ,  ����  �����  ������  �����  ����      B  , ,  �j���  �j����  �����  ����  �j���      B  , ,  �����  ������  �h����  �h���  �����      B  , ,  ����  �����  ������  �����  ����      B  , ,  �f���  �f����  �����  ����  �f���      B  , ,  º���  º����  �d����  �d���  º���      B  , ,  ����  �����  ĸ����  ĸ���  ����      B  , ,  �b���  �b����  �����  ����  �b���      B  , ,  ƶ���  ƶ����  �`����  �`���  ƶ���      B  , ,  �
���  �
����  ȴ����  ȴ���  �
���      B  , ,  �^���  �^����  �����  ����  �^���      B  , ,  ʲ���  ʲ����  �\����  �\���  ʲ���      B  , ,  ����  �����  ̰����  ̰���  ����      B  , ,  �Z���  �Z����  �����  ����  �Z���      B  , ,  ή���  ή����  �X����  �X���  ή���      B  , ,  �����  �����  ������  ������  �����      B  , ,  �Z����  �Z����  �����  �����  �Z����      B  , ,  �h����  �h����  �����  �����  �h����      B  , ,  �h����  �h���3  ����3  �����  �h����      B  , ,  �.���S  �.����  ������  �����S  �.���S      B  , ,  �h����  �h���/  ����/  �����  �h����      B  , ,  �.����  �.���Q  �����Q  ������  �.����      B  , ,  �h����  �h����  �����  �����  �h����      B  , ,  �����  ����}  Ь���}  Ь����  �����      B  , ,  �V����  �V���}  � ���}  � ����  �V����      B  , ,  �.����  �.����  ������  ������  �.����      B  , ,  �h���-  �h����  �����  ����-  �h���-      B  , ,  �.����  �.����  ������  ������  �.����      B  , ,  �h���1  �h����  �����  ����1  �h���1      B  , ,  ����  �����  Ь����  Ь���  ����      B  , ,  �V���  �V����  � ����  � ���  �V���      B  , ,  �����  ����5  Ь���5  Ь����  �����      B  , ,  �V����  �V���5  � ���5  � ����  �V����      B  , ,  �"���I  �"����  ������  �����I  �"���I      B  , ,  �p���I  �p����  �����  ����I  �p���I      B  , ,  �����I  ������  �h����  �h���I  �����I      B  , ,  ����I  �����  ������  �����I  ����I      B  , ,  �Z���I  �Z����  �����  ����I  �Z���I      B  , ,  Ũ���I  Ũ����  �R����  �R���I  Ũ���I      B  , ,  �����I  ������  Ƞ����  Ƞ���I  �����I      B  , ,  �D���I  �D����  ������  �����I  �D���I      B  , ,  �����A  ������  �h����  �h���A  �����A      B  , ,  ����A  �����  ������  �����A  ����A      B  , ,  �Z���A  �Z����  �����  ����A  �Z���A      B  , ,  Ũ���A  Ũ����  �R����  �R���A  Ũ���A      B  , ,  �����A  ������  Ƞ����  Ƞ���A  �����A      B  , ,  �D���A  �D����  ������  �����A  �D���A      B  , ,  �"����  �"����  ������  ������  �"����      B  , ,  �p����  �p����  �����  �����  �p����      B  , ,  ������  ������  �h����  �h����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �Z����  �Z����  �����  �����  �Z����      B  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      B  , ,  ������  ������  Ƞ����  Ƞ����  ������      B  , ,  �D����  �D����  ������  ������  �D����      B  , ,  �"����  �"���C  �����C  ������  �"����      B  , ,  �p����  �p���C  ����C  �����  �p����      B  , ,  ������  �����C  �h���C  �h����  ������      B  , ,  �����  ����C  �����C  ������  �����      B  , ,  �Z����  �Z���C  ����C  �����  �Z����      B  , ,  Ũ����  Ũ���C  �R���C  �R����  Ũ����      B  , ,  ������  �����C  Ƞ���C  Ƞ����  ������      B  , ,  �D����  �D���C  �����C  ������  �D����      B  , ,  �"���E  �"����  ������  �����E  �"���E      B  , ,  �p���E  �p����  �����  ����E  �p���E      B  , ,  �����E  ������  �h����  �h���E  �����E      B  , ,  ����E  �����  ������  �����E  ����E      B  , ,  �Z���E  �Z����  �����  ����E  �Z���E      B  , ,  Ũ���E  Ũ����  �R����  �R���E  Ũ���E      B  , ,  �����E  ������  Ƞ����  Ƞ���E  �����E      B  , ,  �D���E  �D����  ������  �����E  �D���E      B  , ,  �"����  �"����  ������  ������  �"����      B  , ,  �p����  �p����  �����  �����  �p����      B  , ,  ������  ������  �h����  �h����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �Z����  �Z����  �����  �����  �Z����      B  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      B  , ,  ������  ������  Ƞ����  Ƞ����  ������      B  , ,  �D����  �D����  ������  ������  �D����      B  , ,  �"����  �"���G  �����G  ������  �"����      B  , ,  �p����  �p���G  ����G  �����  �p����      B  , ,  ������  �����G  �h���G  �h����  ������      B  , ,  �����  ����G  �����G  ������  �����      B  , ,  �Z����  �Z���G  ����G  �����  �Z����      B  , ,  Ũ����  Ũ���G  �R���G  �R����  Ũ����      B  , ,  ������  �����G  Ƞ���G  Ƞ����  ������      B  , ,  �D����  �D���G  �����G  ������  �D����      B  , ,  ������  �����?  �h���?  �h����  ������      B  , ,  �����  ����?  �����?  ������  �����      B  , ,  �Z����  �Z���?  ����?  �����  �Z����      B  , ,  Ũ����  Ũ���?  �R���?  �R����  Ũ����      B  , ,  ������  �����?  Ƞ���?  Ƞ����  ������      B  , ,  �D����  �D���?  �����?  ������  �D����      B  , ,  �"���A  �"����  ������  �����A  �"���A      B  , ,  �p���A  �p����  �����  ����A  �p���A      B  , ,  �"����  �"���?  �����?  ������  �"����      B  , ,  �p����  �p���?  ����?  �����  �p����      B  , ,  ������  �����}  �A���}  �A����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �3����  �3���}  �����}  ������  �3����      B  , ,  ā����  ā���}  �+���}  �+����  ā����      B  , ,  ������  �����}  �y���}  �y����  ������      B  , ,  �����  ����}  �����}  ������  �����      B  , ,  �k����  �k���}  ����}  �����  �k����      B  , ,  ͹����  ͹���}  �c���}  �c����  ͹����      B  , ,  ������  �����a  �����a  ������  ������      B  , ,  �I����  �I���a  �����a  ������  �I����      B  , ,  ������  �����a  �A���a  �A����  ������      B  , ,  ������  �����a  �����a  ������  ������      B  , ,  �3����  �3���a  �����a  ������  �3����      B  , ,  ā����  ā���a  �+���a  �+����  ā����      B  , ,  ������  �����a  �y���a  �y����  ������      B  , ,  �����  ����a  �����a  ������  �����      B  , ,  �k����  �k���a  ����a  �����  �k����      B  , ,  ͹����  ͹���a  �c���a  �c����  ͹����      B  , ,  �"���A  �"����  ������  �����A  �"���A      B  , ,  �p���A  �p����  �����  ����A  �p���A      B  , ,  �����A  ������  �h����  �h���A  �����A      B  , ,  ����A  �����  ������  �����A  ����A      B  , ,  �Z���A  �Z����  �����  ����A  �Z���A      B  , ,  Ũ���A  Ũ����  �R����  �R���A  Ũ���A      B  , ,  �����A  ������  Ƞ����  Ƞ���A  �����A      B  , ,  �D���A  �D����  ������  �����A  �D���A      B  , ,  �"����  �"����  ������  ������  �"����      B  , ,  �p����  �p����  �����  �����  �p����      B  , ,  ������  ������  �h����  �h����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �Z����  �Z����  �����  �����  �Z����      B  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      B  , ,  ������  ������  Ƞ����  Ƞ����  ������      B  , ,  �D����  �D����  ������  ������  �D����      B  , ,  �"����  �"���C  �����C  ������  �"����      B  , ,  �p����  �p���C  ����C  �����  �p����      B  , ,  ������  �����C  �h���C  �h����  ������      B  , ,  �����  ����C  �����C  ������  �����      B  , ,  �Z����  �Z���C  ����C  �����  �Z����      B  , ,  Ũ����  Ũ���C  �R���C  �R����  Ũ����      B  , ,  ������  �����C  Ƞ���C  Ƞ����  ������      B  , ,  �D����  �D���C  �����C  ������  �D����      B  , ,  �"���E  �"����  ������  �����E  �"���E      B  , ,  �p���E  �p����  �����  ����E  �p���E      B  , ,  �����E  ������  �h����  �h���E  �����E      B  , ,  ����E  �����  ������  �����E  ����E      B  , ,  �Z���E  �Z����  �����  ����E  �Z���E      B  , ,  Ũ���E  Ũ����  �R����  �R���E  Ũ���E      B  , ,  �����E  ������  Ƞ����  Ƞ���E  �����E      B  , ,  �D���E  �D����  ������  �����E  �D���E      B  , ,  �"����  �"����  ������  ������  �"����      B  , ,  �p����  �p����  �����  �����  �p����      B  , ,  ������  ������  �h����  �h����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �Z����  �Z����  �����  �����  �Z����      B  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      B  , ,  ������  ������  Ƞ����  Ƞ����  ������      B  , ,  �D����  �D����  ������  ������  �D����      B  , ,  �"����  �"���G  �����G  ������  �"����      B  , ,  �p����  �p���G  ����G  �����  �p����      B  , ,  ������  �����G  �h���G  �h����  ������      B  , ,  �����  ����G  �����G  ������  �����      B  , ,  �Z����  �Z���G  ����G  �����  �Z����      B  , ,  Ũ����  Ũ���G  �R���G  �R����  Ũ����      B  , ,  ������  �����G  Ƞ���G  Ƞ����  ������      B  , ,  �D����  �D���G  �����G  ������  �D����      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �I����  �I���}  �����}  ������  �I����      B  , ,  �����  ����}  б���}  б����  �����      B  , ,  �����  ����a  б���a  б����  �����      B  , ,  ������  �����M  �f���M  �f����  ������      B  , ,  �����O  ������  �f����  �f���O  �����O      B  , ,  ������  ������  �f����  �f����  ������      B  , ,  ������  ������  �f����  �f����  ������      B  , ,  ������  �����Q  �f���Q  �f����  ������      B  , ,  �����S  ������  �f����  �f���S  �����S      B  , ,  �����S  ������  �f����  �f���S  �����S      B  , ,  ������  ������  �f����  �f����  ������      B  , ,  ������  �����5  �H���5  �H����  ������      B  , ,  ������  �����}  �H���}  �H����  ������      B  , ,  �����  ������  �H����  �H���  �����      B  , ,  �����K  ������  �f����  �f���K  �����K      B  , ,  ������  �����Q  �f���Q  �f����  ������      B  , ,  ������  ������  �f����  �f����  ������      B  , ,  ������  �����Q  �r���Q  �r����  ������      B  , ,  ������  �����M  �r���M  �r����  ������      B  , ,  �
���O  �
����  ������  �����O  �
���O      B  , ,  �X���O  �X����  �����  ����O  �X���O      B  , ,  �����O  ������  �P����  �P���O  �����O      B  , ,  �����O  ������  ������  �����O  �����O      B  , ,  �B���O  �B����  ������  �����O  �B���O      B  , ,  �����O  ������  �:����  �:���O  �����O      B  , ,  �����O  ������  ������  �����O  �����O      B  , ,  �,���O  �,����  ������  �����O  �,���O      B  , ,  �z���O  �z����  �$����  �$���O  �z���O      B  , ,  �����O  ������  �r����  �r���O  �����O      B  , ,  ����O  �����  ������  �����O  ����O      B  , ,  �d���O  �d����  �����  ����O  �d���O      B  , ,  �����O  ������  �\����  �\���O  �����O      B  , ,  � ���O  � ����  ������  �����O  � ���O      B  , ,  �N���O  �N����  ������  �����O  �N���O      B  , ,  �����O  ������  �F����  �F���O  �����O      B  , ,  �����O  ������  ������  �����O  �����O      B  , ,  �8���O  �8����  ������  �����O  �8���O      B  , ,  �����O  ������  �0����  �0���O  �����O      B  , ,  �����O  ������  �~����  �~���O  �����O      B  , ,  ������  ������  �r����  �r����  ������      B  , ,  ������  �����Q  �r���Q  �r����  ������      B  , ,  �����S  ������  �r����  �r���S  �����S      B  , ,  �����S  ������  �r����  �r���S  �����S      B  , ,  ������  ������  �r����  �r����  ������      B  , ,  ������  ������  �r����  �r����  ������      B  , ,  �����K  ������  �r����  �r���K  �����K      B  , ,  ������  ������  �r����  �r����  ������      B  , ,  � ����  � ���M  �����M  ������  � ����      B  , ,  �N����  �N���M  �����M  ������  �N����      B  , ,  ������  �����M  �F���M  �F����  ������      B  , ,  ������  �����M  �����M  ������  ������      B  , ,  �8����  �8���M  �����M  ������  �8����      B  , ,  ������  �����M  �0���M  �0����  ������      B  , ,  ������  �����M  �~���M  �~����  ������      B  , ,  ������  �����Q  �\���Q  �\����  ������      B  , ,  � ����  � ���Q  �����Q  ������  � ����      B  , ,  �N����  �N���Q  �����Q  ������  �N����      B  , ,  ������  �����Q  �F���Q  �F����  ������      B  , ,  ������  �����Q  �����Q  ������  ������      B  , ,  �8����  �8���Q  �����Q  ������  �8����      B  , ,  ������  �����Q  �0���Q  �0����  ������      B  , ,  �8����  �8����  ������  ������  �8����      B  , ,  ������  ������  �0����  �0����  ������      B  , ,  ������  �����Q  �~���Q  �~����  ������      B  , ,  ������  ������  �~����  �~����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �d����  �d���Q  ����Q  �����  �d����      B  , ,  ������  ������  �F����  �F����  ������      B  , ,  ����S  �����  ������  �����S  ����S      B  , ,  �d���S  �d����  �����  ����S  �d���S      B  , ,  �����S  ������  �\����  �\���S  �����S      B  , ,  � ���S  � ����  ������  �����S  � ���S      B  , ,  �N���S  �N����  ������  �����S  �N���S      B  , ,  �����S  ������  �F����  �F���S  �����S      B  , ,  �����S  ������  ������  �����S  �����S      B  , ,  �8���S  �8����  ������  �����S  �8���S      B  , ,  �����S  ������  �0����  �0���S  �����S      B  , ,  �����  ����Q  �����Q  ������  �����      B  , ,  �����S  ������  �~����  �~���S  �����S      B  , ,  �����  ����M  �����M  ������  �����      B  , ,  �����  �����  ������  ������  �����      B  , ,  �d����  �d����  �����  �����  �d����      B  , ,  ������  ������  �\����  �\����  ������      B  , ,  � ����  � ����  ������  ������  � ����      B  , ,  �N����  �N����  ������  ������  �N����      B  , ,  ������  ������  �F����  �F����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �=����  �=����  ������  ������  �=����      B  , ,  ������  ������  �5����  �5����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �'����  �'����  ������  ������  �'����      B  , ,  �u����  �u����  �����  �����  �u����      B  , ,  ������  ������  �m����  �m����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �_����  �_����  �	����  �	����  �_����      B  , ,  ������  ������  �W����  �W����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �8����  �8����  ������  ������  �8����      B  , ,  ������  ������  �0����  �0����  ������      B  , ,  ������  ������  �~����  �~����  ������      B  , ,  ������  �����k  �����k  ������  ������      B  , ,  �=����  �=���k  �����k  ������  �=����      B  , ,  ������  �����k  �5���k  �5����  ������      B  , ,  ������  �����k  �����k  ������  ������      B  , ,  �'����  �'���k  �����k  ������  �'����      B  , ,  �u����  �u���k  ����k  �����  �u����      B  , ,  ������  �����k  �m���k  �m����  ������      B  , ,  �����  ����k  �����k  ������  �����      B  , ,  �_����  �_���k  �	���k  �	����  �_����      B  , ,  ������  �����k  �W���k  �W����  ������      B  , ,  �d����  �d���M  ����M  �����  �d����      B  , ,  ����K  �����  ������  �����K  ����K      B  , ,  �d���K  �d����  �����  ����K  �d���K      B  , ,  �����K  ������  �\����  �\���K  �����K      B  , ,  � ���K  � ����  ������  �����K  � ���K      B  , ,  �N���K  �N����  ������  �����K  �N���K      B  , ,  �����K  ������  �F����  �F���K  �����K      B  , ,  �����K  ������  ������  �����K  �����K      B  , ,  �8���K  �8����  ������  �����K  �8���K      B  , ,  �����K  ������  �0����  �0���K  �����K      B  , ,  �����K  ������  �~����  �~���K  �����K      B  , ,  ������  �����M  �\���M  �\����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �d����  �d����  �����  �����  �d����      B  , ,  ������  ������  �\����  �\����  ������      B  , ,  � ����  � ����  ������  ������  � ����      B  , ,  �N����  �N����  ������  ������  �N����      B  , ,  ������  ������  �K����  �K����  ������      B  , ,  �X����  �X���Q  ����Q  �����  �X����      B  , ,  �
����  �
���M  �����M  ������  �
����      B  , ,  �,���S  �,����  ������  �����S  �,���S      B  , ,  �z���S  �z����  �$����  �$���S  �z���S      B  , ,  �X����  �X���M  ����M  �����  �X����      B  , ,  ������  �����M  �P���M  �P����  ������      B  , ,  ������  �����M  �����M  ������  ������      B  , ,  �B����  �B���M  �����M  ������  �B����      B  , ,  �
����  �
����  ������  ������  �
����      B  , ,  ������  �����Q  �:���Q  �:����  ������      B  , ,  �X����  �X����  �����  �����  �X����      B  , ,  ������  ������  �P����  �P����  ������      B  , ,  ������  �����M  �:���M  �:����  ������      B  , ,  ������  �����M  �����M  ������  ������      B  , ,  �,����  �,���M  �����M  ������  �,����      B  , ,  ������  �����k  �����k  ������  ������      B  , ,  �1����  �1���k  �����k  ������  �1����      B  , ,  �����  ����k  �)���k  �)����  �����      B  , ,  ������  �����k  �w���k  �w����  ������      B  , ,  �����  ����k  �����k  ������  �����      B  , ,  �i����  �i���k  ����k  �����  �i����      B  , ,  ������  �����k  �a���k  �a����  ������      B  , ,  �����  ����k  �����k  ������  �����      B  , ,  �S����  �S���k  �����k  ������  �S����      B  , ,  ������  �����k  �K���k  �K����  ������      B  , ,  ������  �����Q  �P���Q  �P����  ������      B  , ,  �z����  �z���M  �$���M  �$����  �z����      B  , ,  �
����  �
���Q  �����Q  ������  �
����      B  , ,  ������  ������  ������  ������  ������      B  , ,  �B����  �B����  ������  ������  �B����      B  , ,  ������  ������  �:����  �:����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �,����  �,����  ������  ������  �,����      B  , ,  �z����  �z����  �$����  �$����  �z����      B  , ,  �
���S  �
����  ������  �����S  �
���S      B  , ,  ������  �����Q  �����Q  ������  ������      B  , ,  �
���K  �
����  ������  �����K  �
���K      B  , ,  �X���K  �X����  �����  ����K  �X���K      B  , ,  �����K  ������  �P����  �P���K  �����K      B  , ,  �����K  ������  ������  �����K  �����K      B  , ,  �B���K  �B����  ������  �����K  �B���K      B  , ,  �����K  ������  �:����  �:���K  �����K      B  , ,  �����K  ������  ������  �����K  �����K      B  , ,  �,���K  �,����  ������  �����K  �,���K      B  , ,  �z���K  �z����  �$����  �$���K  �z���K      B  , ,  �X���S  �X����  �����  ����S  �X���S      B  , ,  �����S  ������  �P����  �P���S  �����S      B  , ,  �����S  ������  ������  �����S  �����S      B  , ,  �B���S  �B����  ������  �����S  �B���S      B  , ,  �����S  ������  �:����  �:���S  �����S      B  , ,  ������  �����Q  �����Q  ������  ������      B  , ,  �����S  ������  ������  �����S  �����S      B  , ,  �B����  �B���Q  �����Q  ������  �B����      B  , ,  ������  ������  ������  ������  ������      B  , ,  �1����  �1����  ������  ������  �1����      B  , ,  �����  �����  �)����  �)����  �����      B  , ,  �,����  �,���Q  �����Q  ������  �,����      B  , ,  �z����  �z���Q  �$���Q  �$����  �z����      B  , ,  �
����  �
����  ������  ������  �
����      B  , ,  �X����  �X����  �����  �����  �X����      B  , ,  ������  ������  �P����  �P����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �B����  �B����  ������  ������  �B����      B  , ,  ������  ������  �:����  �:����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �,����  �,����  ������  ������  �,����      B  , ,  �z����  �z����  �$����  �$����  �z����      B  , ,  ������  ������  �w����  �w����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �i����  �i����  �����  �����  �i����      B  , ,  ������  ������  �a����  �a����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �S����  �S����  ������  ������  �S����      B  , ,  ������  ������  ������  ������  ������      B  , ,  �B����  �B����  ������  ������  �B����      B  , ,  ������  ������  �:����  �:����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �,����  �,����  ������  ������  �,����      B  , ,  �z����  �z����  �$����  �$����  �z����      B  , ,  �z����  �z����  �$����  �$����  �z����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �F���  �F����  ������  �����  �F���      B  , ,  �����  ������  �D����  �D���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �B���  �B����  ������  �����  �B���      B  , ,  �����  ������  �@����  �@���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �>���  �>����  ������  �����  �>���      B  , ,  �����  ������  �<����  �<���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �:���  �:����  ������  �����  �:���      B  , ,  �����  ������  �8����  �8���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �6���  �6����  ������  �����  �6���      B  , ,  �����  ������  �4����  �4���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �2���  �2����  ������  �����  �2���      B  , ,  �
����  �
����  ������  ������  �
����      B  , ,  �X����  �X����  �����  �����  �X����      B  , ,  �
����  �
���Q  �����Q  ������  �
����      B  , ,  �
���S  �
����  ������  �����S  �
���S      B  , ,  �X���S  �X����  �����  ����S  �X���S      B  , ,  �����S  ������  �P����  �P���S  �����S      B  , ,  �����S  ������  ������  �����S  �����S      B  , ,  �B���S  �B����  ������  �����S  �B���S      B  , ,  �����S  ������  �:����  �:���S  �����S      B  , ,  �����S  ������  ������  �����S  �����S      B  , ,  �,���S  �,����  ������  �����S  �,���S      B  , ,  �z���S  �z����  �$����  �$���S  �z���S      B  , ,  �X����  �X���Q  ����Q  �����  �X����      B  , ,  ������  �����Q  �P���Q  �P����  ������      B  , ,  ������  �����5  �����5  ������  ������      B  , ,  �F����  �F���5  �����5  ������  �F����      B  , ,  ������  �����5  �D���5  �D����  ������      B  , ,  ������  �����5  �����5  ������  ������      B  , ,  �B����  �B���5  �����5  ������  �B����      B  , ,  ������  �����5  �@���5  �@����  ������      B  , ,  ������  �����5  �����5  ������  ������      B  , ,  �>����  �>���5  �����5  ������  �>����      B  , ,  ������  �����5  �<���5  �<����  ������      B  , ,  ������  �����5  �����5  ������  ������      B  , ,  �:����  �:���5  �����5  ������  �:����      B  , ,  ������  �����5  �8���5  �8����  ������      B  , ,  ������  �����5  �����5  ������  ������      B  , ,  �6����  �6���5  �����5  ������  �6����      B  , ,  ������  �����5  �4���5  �4����  ������      B  , ,  ������  �����5  �����5  ������  ������      B  , ,  �2����  �2���5  �����5  ������  �2����      B  , ,  ������  �����Q  �����Q  ������  ������      B  , ,  �B����  �B���Q  �����Q  ������  �B����      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �F����  �F���}  �����}  ������  �F����      B  , ,  ������  �����}  �D���}  �D����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �B����  �B���}  �����}  ������  �B����      B  , ,  ������  �����}  �@���}  �@����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �>����  �>���}  �����}  ������  �>����      B  , ,  ������  �����}  �<���}  �<����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �:����  �:���}  �����}  ������  �:����      B  , ,  ������  �����}  �8���}  �8����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �6����  �6���}  �����}  ������  �6����      B  , ,  ������  �����}  �4���}  �4����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �2����  �2���}  �����}  ������  �2����      B  , ,  ������  �����Q  �:���Q  �:����  ������      B  , ,  ������  �����Q  �����Q  ������  ������      B  , ,  �,����  �,���Q  �����Q  ������  �,����      B  , ,  �z����  �z���Q  �$���Q  �$����  �z����      B  , ,  ������  ������  �P����  �P����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �B����  �B����  ������  ������  �B����      B  , ,  ������  ������  �:����  �:����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �,����  �,����  ������  ������  �,����      B  , ,  �
����  �
����  ������  ������  �
����      B  , ,  �X����  �X����  �����  �����  �X����      B  , ,  ������  ������  �P����  �P����  ������      B  , ,  �*����  �*���5  �����5  ������  �*����      B  , ,  �~����  �~���5  �(���5  �(����  �~����      B  , ,  ������  �����5  �|���5  �|����  ������      B  , ,  �&����  �&���5  �����5  ������  �&����      B  , ,  �z����  �z���5  �$���5  �$����  �z����      B  , ,  ������  �����5  �x���5  �x����  ������      B  , ,  �"����  �"���5  �����5  ������  �"����      B  , ,  �v����  �v���5  � ���5  � ����  �v����      B  , ,  ������  �����5  �t���5  �t����  ������      B  , ,  �����  ����5  �����5  ������  �����      B  , ,  �r����  �r���5  ����5  �����  �r����      B  , ,  �����  ������  �0����  �0���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �.���  �.����  ������  �����  �.���      B  , ,  �����  ������  �,����  �,���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �*���  �*����  ������  �����  �*���      B  , ,  �~���  �~����  �(����  �(���  �~���      B  , ,  �����  ������  �|����  �|���  �����      B  , ,  �&���  �&����  ������  �����  �&���      B  , ,  �z���  �z����  �$����  �$���  �z���      B  , ,  �����  ������  �x����  �x���  �����      B  , ,  �"���  �"����  ������  �����  �"���      B  , ,  �v���  �v����  � ����  � ���  �v���      B  , ,  �����  ������  �t����  �t���  �����      B  , ,  ����  �����  ������  �����  ����      B  , ,  �r���  �r����  �����  ����  �r���      B  , ,  �����  ������  �p����  �p���  �����      B  , ,  ������  �����5  �p���5  �p����  ������      B  , ,  �d����  �d����  �����  �����  �d����      B  , ,  ������  ������  �\����  �\����  ������      B  , ,  � ����  � ����  ������  ������  � ����      B  , ,  �N����  �N����  ������  ������  �N����      B  , ,  ������  ������  �F����  �F����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �8����  �8����  ������  ������  �8����      B  , ,  ������  ������  �0����  �0����  ������      B  , ,  ������  ������  �~����  �~����  ������      B  , ,  � ���S  � ����  ������  �����S  � ���S      B  , ,  �N���S  �N����  ������  �����S  �N���S      B  , ,  �����S  ������  �F����  �F���S  �����S      B  , ,  �����S  ������  ������  �����S  �����S      B  , ,  �8���S  �8����  ������  �����S  �8���S      B  , ,  �����S  ������  �0����  �0���S  �����S      B  , ,  �����S  ������  �~����  �~���S  �����S      B  , ,  ������  �����Q  �~���Q  �~����  ������      B  , ,  �d����  �d����  �����  �����  �d����      B  , ,  ������  ������  �\����  �\����  ������      B  , ,  ������  �����}  �0���}  �0����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �.����  �.���}  �����}  ������  �.����      B  , ,  ������  �����}  �,���}  �,����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �*����  �*���}  �����}  ������  �*����      B  , ,  �~����  �~���}  �(���}  �(����  �~����      B  , ,  ������  �����}  �|���}  �|����  ������      B  , ,  �&����  �&���}  �����}  ������  �&����      B  , ,  �z����  �z���}  �$���}  �$����  �z����      B  , ,  ������  �����}  �x���}  �x����  ������      B  , ,  �"����  �"���}  �����}  ������  �"����      B  , ,  �v����  �v���}  � ���}  � ����  �v����      B  , ,  ������  �����}  �t���}  �t����  ������      B  , ,  �����  ����}  �����}  ������  �����      B  , ,  �r����  �r���}  ����}  �����  �r����      B  , ,  ������  �����}  �p���}  �p����  ������      B  , ,  � ����  � ����  ������  ������  � ����      B  , ,  �N����  �N����  ������  ������  �N����      B  , ,  ������  ������  �F����  �F����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �8����  �8����  ������  ������  �8����      B  , ,  ������  ������  �0����  �0����  ������      B  , ,  ������  ������  �~����  �~����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �����  ����Q  �����Q  ������  �����      B  , ,  �d����  �d���Q  ����Q  �����  �d����      B  , ,  ������  �����Q  �\���Q  �\����  ������      B  , ,  � ����  � ���Q  �����Q  ������  � ����      B  , ,  �N����  �N���Q  �����Q  ������  �N����      B  , ,  ������  �����Q  �F���Q  �F����  ������      B  , ,  ������  �����Q  �����Q  ������  ������      B  , ,  �8����  �8���Q  �����Q  ������  �8����      B  , ,  ������  �����Q  �0���Q  �0����  ������      B  , ,  ����S  �����  ������  �����S  ����S      B  , ,  �d���S  �d����  �����  ����S  �d���S      B  , ,  �����S  ������  �\����  �\���S  �����S      B  , ,  �����  �����  ������  ������  �����      B  , ,  ������  �����5  �0���5  �0����  ������      B  , ,  ������  �����5  �����5  ������  ������      B  , ,  �.����  �.���5  �����5  ������  �.����      B  , ,  ������  �����5  �,���5  �,����  ������      B  , ,  ������  �����5  �����5  ������  ������      B  , ,  [�����  [����+  \b���+  \b����  [�����      B  , ,  r����S  r�����  sZ����  sZ���S  r����S      B  , ,  r�����  r�����  sZ����  sZ����  r�����      B  , ,  ]����O  ]�����  ^�����  ^����O  ]����O      B  , ,  `@���O  `@����  `�����  `����O  `@���O      B  , ,  b����O  b�����  c8����  c8���O  b����O      B  , ,  d����O  d�����  e�����  e����O  d����O      B  , ,  g*���O  g*����  g�����  g����O  g*���O      B  , ,  ix���O  ix����  j"����  j"���O  ix���O      B  , ,  k����O  k�����  lp����  lp���O  k����O      B  , ,  n���O  n����  n�����  n����O  n���O      B  , ,  pb���O  pb����  q����  q���O  pb���O      B  , ,  r����O  r�����  sZ����  sZ���O  r����O      B  , ,  t����O  t�����  u�����  u����O  t����O      B  , ,  r�����  r�����  sZ����  sZ����  r�����      B  , ,  wL���O  wL����  w�����  w����O  wL���O      B  , ,  y����O  y�����  zD����  zD���O  y����O      B  , ,  {����O  {�����  |�����  |����O  {����O      B  , ,  ~6���O  ~6����  ~�����  ~����O  ~6���O      B  , ,  �����O  ������  �.����  �.���O  �����O      B  , ,  �����O  ������  �|����  �|���O  �����O      B  , ,  � ���O  � ����  ������  �����O  � ���O      B  , ,  �n���O  �n����  �����  ����O  �n���O      B  , ,  r�����  r����M  sZ���M  sZ����  r�����      B  , ,  r����S  r�����  sZ����  sZ���S  r����S      B  , ,  r�����  r����Q  sZ���Q  sZ����  r�����      B  , ,  r�����  r�����  sZ����  sZ����  r�����      B  , ,  r����K  r�����  sZ����  sZ���K  r����K      B  , ,  r�����  r����Q  sZ���Q  sZ����  r�����      B  , ,  r�����  r�����  sZ����  sZ����  r�����      B  , ,  t�����  t����M  u����M  u�����  t�����      B  , ,  wL����  wL���M  w����M  w�����  wL����      B  , ,  ������  ������  �?����  �?����  ������      B  , ,  y�����  y����M  zD���M  zD����  y�����      B  , ,  {�����  {����M  |����M  |�����  {�����      B  , ,  ~6����  ~6���M  ~����M  ~�����  ~6����      B  , ,  ������  �����M  �.���M  �.����  ������      B  , ,  ������  �����M  �|���M  �|����  ������      B  , ,  � ����  � ���M  �����M  ������  � ����      B  , ,  �n����  �n���M  ����M  �����  �n����      B  , ,  wL����  wL����  w�����  w�����  wL����      B  , ,  ������  ������  �.����  �.����  ������      B  , ,  ������  ������  �|����  �|����  ������      B  , ,  �����S  ������  �.����  �.���S  �����S      B  , ,  �����S  ������  �|����  �|���S  �����S      B  , ,  � ���S  � ����  ������  �����S  � ���S      B  , ,  �n���S  �n����  �����  ����S  �n���S      B  , ,  � ����  � ����  ������  ������  � ����      B  , ,  �n����  �n����  �����  �����  �n����      B  , ,  y�����  y�����  zD����  zD����  y�����      B  , ,  s�����  s�����  t�����  t�����  s�����      B  , ,  v%����  v%����  v�����  v�����  v%����      B  , ,  xs����  xs����  y����  y����  xs����      B  , ,  z�����  z�����  {k����  {k����  z�����      B  , ,  }����  }����  }�����  }�����  }����      B  , ,  s�����  s����k  t����k  t�����  s�����      B  , ,  v%����  v%���k  v����k  v�����  v%����      B  , ,  xs����  xs���k  y���k  y����  xs����      B  , ,  z�����  z����k  {k���k  {k����  z�����      B  , ,  }����  }���k  }����k  }�����  }����      B  , ,  ]����  ]���k  ����k  �����  ]����      B  , ,  ������  �����k  �U���k  �U����  ������      B  , ,  ������  �����k  �����k  ������  ������      B  , ,  �G����  �G���k  �����k  ������  �G����      B  , ,  ������  �����k  �?���k  �?����  ������      B  , ,  ]����  ]����  �����  �����  ]����      B  , ,  t����S  t�����  u�����  u����S  t����S      B  , ,  wL���S  wL����  w�����  w����S  wL���S      B  , ,  y����S  y�����  zD����  zD���S  y����S      B  , ,  {����S  {�����  |�����  |����S  {����S      B  , ,  ~6���S  ~6����  ~�����  ~����S  ~6���S      B  , ,  ������  ������  �U����  �U����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  t�����  t�����  u�����  u�����  t�����      B  , ,  �G����  �G����  ������  ������  �G����      B  , ,  t����K  t�����  u�����  u����K  t����K      B  , ,  wL���K  wL����  w�����  w����K  wL���K      B  , ,  y����K  y�����  zD����  zD���K  y����K      B  , ,  {����K  {�����  |�����  |����K  {����K      B  , ,  ~6���K  ~6����  ~�����  ~����K  ~6���K      B  , ,  �����K  ������  �.����  �.���K  �����K      B  , ,  �����K  ������  �|����  �|���K  �����K      B  , ,  � ���K  � ����  ������  �����K  � ���K      B  , ,  �n���K  �n����  �����  ����K  �n���K      B  , ,  {�����  {�����  |�����  |�����  {�����      B  , ,  t�����  t����Q  u����Q  u�����  t�����      B  , ,  wL����  wL���Q  w����Q  w�����  wL����      B  , ,  y�����  y����Q  zD���Q  zD����  y�����      B  , ,  {�����  {����Q  |����Q  |�����  {�����      B  , ,  ~6����  ~6���Q  ~����Q  ~�����  ~6����      B  , ,  ������  �����Q  �.���Q  �.����  ������      B  , ,  ������  �����Q  �|���Q  �|����  ������      B  , ,  � ����  � ���Q  �����Q  ������  � ����      B  , ,  �n����  �n���Q  ����Q  �����  �n����      B  , ,  ~6����  ~6����  ~�����  ~�����  ~6����      B  , ,  t�����  t�����  u�����  u�����  t�����      B  , ,  wL����  wL����  w�����  w�����  wL����      B  , ,  y�����  y�����  zD����  zD����  y�����      B  , ,  {�����  {�����  |�����  |�����  {�����      B  , ,  ~6����  ~6����  ~�����  ~�����  ~6����      B  , ,  ������  ������  �.����  �.����  ������      B  , ,  ������  ������  �|����  �|����  ������      B  , ,  � ����  � ����  ������  ������  � ����      B  , ,  �n����  �n����  �����  �����  �n����      B  , ,  hQ����  hQ����  h�����  h�����  hQ����      B  , ,  j�����  j�����  kI����  kI����  j�����      B  , ,  l�����  l�����  m�����  m�����  l�����      B  , ,  o;����  o;����  o�����  o�����  o;����      B  , ,  q�����  q�����  r3����  r3����  q�����      B  , ,  ]�����  ]����M  ^����M  ^�����  ]�����      B  , ,  `@����  `@���M  `����M  `�����  `@����      B  , ,  b�����  b����M  c8���M  c8����  b�����      B  , ,  d�����  d����M  e����M  e�����  d�����      B  , ,  g*����  g*���M  g����M  g�����  g*����      B  , ,  ix����  ix���M  j"���M  j"����  ix����      B  , ,  k�����  k����M  lp���M  lp����  k�����      B  , ,  n����  n���M  n����M  n�����  n����      B  , ,  [�����  [����  \b���  \b����  [�����      B  , ,  [����y  [����#  \b���#  \b���y  [����y      B  , ,  _����  _����  _�����  _�����  _����      B  , ,  n����  n����  n�����  n�����  n����      B  , ,  pb����  pb����  q����  q����  pb����      B  , ,  ag����  ag����  b����  b����  ag����      B  , ,  [����!  [�����  \b����  \b���!  [����!      B  , ,  [����u  [����  \b���  \b���u  [����u      B  , ,  ]�����  ]����Q  ^����Q  ^�����  ]�����      B  , ,  `@����  `@���Q  `����Q  `�����  `@����      B  , ,  b�����  b����Q  c8���Q  c8����  b�����      B  , ,  d�����  d����Q  e����Q  e�����  d�����      B  , ,  g*����  g*���Q  g����Q  g�����  g*����      B  , ,  ix����  ix���Q  j"���Q  j"����  ix����      B  , ,  k�����  k����Q  lp���Q  lp����  k�����      B  , ,  [�����  [����{  \b���{  \b����  [�����      B  , ,  n����  n���Q  n����Q  n�����  n����      B  , ,  [����}  [����'  \b���'  \b���}  [����}      B  , ,  ]����K  ]�����  ^�����  ^����K  ]����K      B  , ,  `@���K  `@����  `�����  `����K  `@���K      B  , ,  b����K  b�����  c8����  c8���K  b����K      B  , ,  d����K  d�����  e�����  e����K  d����K      B  , ,  g*���K  g*����  g�����  g����K  g*���K      B  , ,  ix���K  ix����  j"����  j"���K  ix���K      B  , ,  k����K  k�����  lp����  lp���K  k����K      B  , ,  n���K  n����  n�����  n����K  n���K      B  , ,  pb���K  pb����  q����  q���K  pb���K      B  , ,  ]����S  ]�����  ^�����  ^����S  ]����S      B  , ,  c�����  c�����  d_����  d_����  c�����      B  , ,  `@���S  `@����  `�����  `����S  `@���S      B  , ,  pb����  pb���M  q���M  q����  pb����      B  , ,  b����S  b�����  c8����  c8���S  b����S      B  , ,  d����S  d�����  e�����  e����S  d����S      B  , ,  g*���S  g*����  g�����  g����S  g*���S      B  , ,  ix���S  ix����  j"����  j"���S  ix���S      B  , ,  k����S  k�����  lp����  lp���S  k����S      B  , ,  n���S  n����  n�����  n����S  n���S      B  , ,  [�����  [����w  \b���w  \b����  [�����      B  , ,  pb����  pb���Q  q���Q  q����  pb����      B  , ,  pb���S  pb����  q����  q���S  pb���S      B  , ,  [�����  [����s  \b���s  \b����  [�����      B  , ,  ]�����  ]�����  ^�����  ^�����  ]�����      B  , ,  `@����  `@����  `�����  `�����  `@����      B  , ,  b�����  b�����  c8����  c8����  b�����      B  , ,  d�����  d�����  e�����  e�����  d�����      B  , ,  g*����  g*����  g�����  g�����  g*����      B  , ,  ix����  ix����  j"����  j"����  ix����      B  , ,  k�����  k�����  lp����  lp����  k�����      B  , ,  [����%  [�����  \b����  \b���%  [����%      B  , ,  [����)  [�����  \b����  \b���)  [����)      B  , ,  ]�����  ]�����  ^�����  ^�����  ]�����      B  , ,  `@����  `@����  `�����  `�����  `@����      B  , ,  b�����  b�����  c8����  c8����  b�����      B  , ,  d�����  d�����  e�����  e�����  d�����      B  , ,  g*����  g*����  g�����  g�����  g*����      B  , ,  ix����  ix����  j"����  j"����  ix����      B  , ,  k�����  k�����  lp����  lp����  k�����      B  , ,  n����  n����  n�����  n�����  n����      B  , ,  pb����  pb����  q����  q����  pb����      B  , ,  _����  _���k  _����k  _�����  _����      B  , ,  ag����  ag���k  b���k  b����  ag����      B  , ,  c�����  c����k  d_���k  d_����  c�����      B  , ,  f����  f���k  f����k  f�����  f����      B  , ,  hQ����  hQ���k  h����k  h�����  hQ����      B  , ,  j�����  j����k  kI���k  kI����  j�����      B  , ,  l�����  l����k  m����k  m�����  l�����      B  , ,  o;����  o;���k  o����k  o�����  o;����      B  , ,  q�����  q����k  r3���k  r3����  q�����      B  , ,  f����  f����  f�����  f�����  f����      B  , ,  g*����  g*���Q  g����Q  g�����  g*����      B  , ,  ix����  ix���Q  j"���Q  j"����  ix����      B  , ,  k�����  k����Q  lp���Q  lp����  k�����      B  , ,  n����  n���Q  n����Q  n�����  n����      B  , ,  pb����  pb���Q  q���Q  q����  pb����      B  , ,  c����  c���}  c����}  c�����  c����      B  , ,  [�����  [�����  \b����  \b����  [�����      B  , ,  [�����  [����3  \b���3  \b����  [�����      B  , ,  [����1  [�����  \b����  \b���1  [����1      B  , ,  ]�����  ]�����  ^�����  ^�����  ]�����      B  , ,  `@����  `@����  `�����  `�����  `@����      B  , ,  b�����  b�����  c8����  c8����  b�����      B  , ,  d�����  d�����  e�����  e�����  d�����      B  , ,  g*����  g*����  g�����  g�����  g*����      B  , ,  ix����  ix����  j"����  j"����  ix����      B  , ,  k�����  k�����  lp����  lp����  k�����      B  , ,  n����  n����  n�����  n�����  n����      B  , ,  pb����  pb����  q����  q����  pb����      B  , ,  [�����  [����/  \b���/  \b����  [�����      B  , ,  ]����S  ]�����  ^�����  ^����S  ]����S      B  , ,  `@���S  `@����  `�����  `����S  `@���S      B  , ,  b����S  b�����  c8����  c8���S  b����S      B  , ,  d����S  d�����  e�����  e����S  d����S      B  , ,  g*���S  g*����  g�����  g����S  g*���S      B  , ,  ix���S  ix����  j"����  j"���S  ix���S      B  , ,  k����S  k�����  lp����  lp���S  k����S      B  , ,  n���S  n����  n�����  n����S  n���S      B  , ,  pb���S  pb����  q����  q���S  pb���S      B  , ,  dn����  dn���}  e���}  e����  dn����      B  , ,  e�����  e����}  fl���}  fl����  e�����      B  , ,  g����  g���}  g����}  g�����  g����      B  , ,  [����-  [�����  \b����  \b���-  [����-      B  , ,  ]�����  ]�����  ^�����  ^�����  ]�����      B  , ,  `@����  `@����  `�����  `�����  `@����      B  , ,  b�����  b�����  c8����  c8����  b�����      B  , ,  d�����  d�����  e�����  e�����  d�����      B  , ,  g*����  g*����  g�����  g�����  g*����      B  , ,  ix����  ix����  j"����  j"����  ix����      B  , ,  k�����  k�����  lp����  lp����  k�����      B  , ,  hj����  hj���}  i���}  i����  hj����      B  , ,  n����  n����  n�����  n�����  n����      B  , ,  pb����  pb����  q����  q����  pb����      B  , ,  i�����  i����}  jh���}  jh����  i�����      B  , ,  ]�����  ]����5  ^t���5  ^t����  ]�����      B  , ,  _����  _���5  _����5  _�����  _����      B  , ,  `r����  `r���5  a���5  a����  `r����      B  , ,  a�����  a����5  bp���5  bp����  a�����      B  , ,  c����  c���5  c����5  c�����  c����      B  , ,  dn����  dn���5  e���5  e����  dn����      B  , ,  e�����  e����5  fl���5  fl����  e�����      B  , ,  g����  g���5  g����5  g�����  g����      B  , ,  hj����  hj���5  i���5  i����  hj����      B  , ,  i�����  i����5  jh���5  jh����  i�����      B  , ,  k����  k���5  k����5  k�����  k����      B  , ,  lf����  lf���5  m���5  m����  lf����      B  , ,  m�����  m����5  nd���5  nd����  m�����      B  , ,  o����  o���5  o����5  o�����  o����      B  , ,  pb����  pb���5  q���5  q����  pb����      B  , ,  q�����  q����5  r`���5  r`����  q�����      B  , ,  k����  k���}  k����}  k�����  k����      B  , ,  lf����  lf���}  m���}  m����  lf����      B  , ,  m�����  m����}  nd���}  nd����  m�����      B  , ,  o����  o���}  o����}  o�����  o����      B  , ,  pb����  pb���}  q���}  q����  pb����      B  , ,  q�����  q����}  r`���}  r`����  q�����      B  , ,  ]�����  ]����}  ^t���}  ^t����  ]�����      B  , ,  ]����  ]�����  ^t����  ^t���  ]����      B  , ,  _���  _����  _�����  _����  _���      B  , ,  `r���  `r����  a����  a���  `r���      B  , ,  a����  a�����  bp����  bp���  a����      B  , ,  c���  c����  c�����  c����  c���      B  , ,  dn���  dn����  e����  e���  dn���      B  , ,  e����  e�����  fl����  fl���  e����      B  , ,  g���  g����  g�����  g����  g���      B  , ,  hj���  hj����  i����  i���  hj���      B  , ,  i����  i�����  jh����  jh���  i����      B  , ,  k���  k����  k�����  k����  k���      B  , ,  lf���  lf����  m����  m���  lf���      B  , ,  m����  m�����  nd����  nd���  m����      B  , ,  o���  o����  o�����  o����  o���      B  , ,  pb���  pb����  q����  q���  pb���      B  , ,  q����  q�����  r`����  r`���  q����      B  , ,  _����  _���}  _����}  _�����  _����      B  , ,  `r����  `r���}  a���}  a����  `r����      B  , ,  a�����  a����}  bp���}  bp����  a�����      B  , ,  [�����  [�����  \b����  \b����  [�����      B  , ,  ]�����  ]����Q  ^����Q  ^�����  ]�����      B  , ,  `@����  `@���Q  `����Q  `�����  `@����      B  , ,  b�����  b����Q  c8���Q  c8����  b�����      B  , ,  d�����  d����Q  e����Q  e�����  d�����      B  , ,  �����S  ������  �|����  �|���S  �����S      B  , ,  � ���S  � ����  ������  �����S  � ���S      B  , ,  �n���S  �n����  �����  ����S  �n���S      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �N����  �N���}  �����}  ������  �N����      B  , ,  ������  �����}  �L���}  �L����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �J����  �J���}  �����}  ������  �J����      B  , ,  �n����  �n���Q  ����Q  �����  �n����      B  , ,  ������  �����Q  �.���Q  �.����  ������      B  , ,  s
���  s
����  s�����  s����  s
���      B  , ,  t^���  t^����  u����  u���  t^���      B  , ,  u����  u�����  v\����  v\���  u����      B  , ,  w���  w����  w�����  w����  w���      B  , ,  xZ���  xZ����  y����  y���  xZ���      B  , ,  y����  y�����  zX����  zX���  y����      B  , ,  {���  {����  {�����  {����  {���      B  , ,  |V���  |V����  } ����  } ���  |V���      B  , ,  }����  }�����  ~T����  ~T���  }����      B  , ,  ~����  ~�����  �����  ����  ~����      B  , ,  �R���  �R����  ������  �����  �R���      B  , ,  �����  ������  �P����  �P���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �N���  �N����  ������  �����  �N���      B  , ,  �����  ������  �L����  �L���  �����      B  , ,  �����  ������  ������  �����  �����      B  , ,  �J���  �J����  ������  �����  �J���      B  , ,  ������  �����Q  �|���Q  �|����  ������      B  , ,  � ����  � ���Q  �����Q  ������  � ����      B  , ,  s
����  s
���}  s����}  s�����  s
����      B  , ,  t^����  t^���}  u���}  u����  t^����      B  , ,  u�����  u����}  v\���}  v\����  u�����      B  , ,  w����  w���}  w����}  w�����  w����      B  , ,  xZ����  xZ���}  y���}  y����  xZ����      B  , ,  t�����  t�����  u�����  u�����  t�����      B  , ,  s
����  s
���5  s����5  s�����  s
����      B  , ,  t^����  t^���5  u���5  u����  t^����      B  , ,  u�����  u����5  v\���5  v\����  u�����      B  , ,  w����  w���5  w����5  w�����  w����      B  , ,  wL����  wL����  w�����  w�����  wL����      B  , ,  y�����  y�����  zD����  zD����  y�����      B  , ,  {�����  {�����  |�����  |�����  {�����      B  , ,  ~6����  ~6����  ~�����  ~�����  ~6����      B  , ,  ������  ������  �.����  �.����  ������      B  , ,  ������  ������  �|����  �|����  ������      B  , ,  � ����  � ����  ������  ������  � ����      B  , ,  t�����  t�����  u�����  u�����  t�����      B  , ,  wL����  wL����  w�����  w�����  wL����      B  , ,  y�����  y�����  zD����  zD����  y�����      B  , ,  {�����  {�����  |�����  |�����  {�����      B  , ,  xZ����  xZ���5  y���5  y����  xZ����      B  , ,  ~6����  ~6����  ~�����  ~�����  ~6����      B  , ,  ������  ������  �.����  �.����  ������      B  , ,  t�����  t����Q  u����Q  u�����  t�����      B  , ,  ������  ������  �|����  �|����  ������      B  , ,  � ����  � ����  ������  ������  � ����      B  , ,  �n����  �n����  �����  �����  �n����      B  , ,  �n����  �n����  �����  �����  �n����      B  , ,  y�����  y����}  zX���}  zX����  y�����      B  , ,  {����  {���}  {����}  {�����  {����      B  , ,  |V����  |V���}  } ���}  } ����  |V����      B  , ,  }�����  }����}  ~T���}  ~T����  }�����      B  , ,  ~�����  ~����}  ����}  �����  ~�����      B  , ,  �R����  �R���}  �����}  ������  �R����      B  , ,  ������  �����}  �P���}  �P����  ������      B  , ,  t����S  t�����  u�����  u����S  t����S      B  , ,  wL���S  wL����  w�����  w����S  wL���S      B  , ,  y����S  y�����  zD����  zD���S  y����S      B  , ,  {����S  {�����  |�����  |����S  {����S      B  , ,  ~6���S  ~6����  ~�����  ~����S  ~6���S      B  , ,  �����S  ������  �.����  �.���S  �����S      B  , ,  y�����  y����5  zX���5  zX����  y�����      B  , ,  {����  {���5  {����5  {�����  {����      B  , ,  |V����  |V���5  } ���5  } ����  |V����      B  , ,  }�����  }����5  ~T���5  ~T����  }�����      B  , ,  ~�����  ~����5  ����5  �����  ~�����      B  , ,  �R����  �R���5  �����5  ������  �R����      B  , ,  ������  �����5  �P���5  �P����  ������      B  , ,  ������  �����5  �����5  ������  ������      B  , ,  �N����  �N���5  �����5  ������  �N����      B  , ,  ������  �����5  �L���5  �L����  ������      B  , ,  ������  �����5  �����5  ������  ������      B  , ,  �J����  �J���5  �����5  ������  �J����      B  , ,  wL����  wL���Q  w����Q  w�����  wL����      B  , ,  y�����  y����Q  zD���Q  zD����  y�����      B  , ,  {�����  {����Q  |����Q  |�����  {�����      B  , ,  ~6����  ~6���Q  ~����Q  ~�����  ~6����      B  , ,  v%����  v%���a  v����a  v�����  v%����      B  , ,  xs����  xs���a  y���a  y����  xs����      B  , ,  z�����  z����a  {k���a  {k����  z�����      B  , ,  }����  }���a  }����a  }�����  }����      B  , ,  ]����  ]���a  ����a  �����  ]����      B  , ,  ������  �����a  �U���a  �U����  ������      B  , ,  ������  �����a  �����a  ������  ������      B  , ,  �G����  �G���a  �����a  ������  �G����      B  , ,  ������  �����a  �?���a  �?����  ������      B  , ,  wL����  wL���G  w����G  w�����  wL����      B  , ,  pb���E  pb����  q����  q���E  pb���E      B  , ,  r����E  r�����  sZ����  sZ���E  r����E      B  , ,  t����E  t�����  u�����  u����E  t����E      B  , ,  wL���E  wL����  w�����  w����E  wL���E      B  , ,  pb���A  pb����  q����  q���A  pb���A      B  , ,  r����A  r�����  sZ����  sZ���A  r����A      B  , ,  t����A  t�����  u�����  u����A  t����A      B  , ,  wL���A  wL����  w�����  w����A  wL���A      B  , ,  pb���I  pb����  q����  q���I  pb���I      B  , ,  r����I  r�����  sZ����  sZ���I  r����I      B  , ,  pb���A  pb����  q����  q���A  pb���A      B  , ,  r����A  r�����  sZ����  sZ���A  r����A      B  , ,  t����A  t�����  u�����  u����A  t����A      B  , ,  wL���A  wL����  w�����  w����A  wL���A      B  , ,  t����I  t�����  u�����  u����I  t����I      B  , ,  wL���I  wL����  w�����  w����I  wL���I      B  , ,  pb����  pb���C  q���C  q����  pb����      B  , ,  r�����  r����C  sZ���C  sZ����  r�����      B  , ,  t�����  t����C  u����C  u�����  t�����      B  , ,  wL����  wL���C  w����C  w�����  wL����      B  , ,  pb����  pb����  q����  q����  pb����      B  , ,  r�����  r�����  sZ����  sZ����  r�����      B  , ,  pb����  pb����  q����  q����  pb����      B  , ,  r�����  r�����  sZ����  sZ����  r�����      B  , ,  t�����  t�����  u�����  u�����  t�����      B  , ,  wL����  wL����  w�����  w�����  wL����      B  , ,  t�����  t�����  u�����  u�����  t�����      B  , ,  wL����  wL����  w�����  w�����  wL����      B  , ,  _����  _���}  _����}  _�����  _����      B  , ,  ag����  ag���}  b���}  b����  ag����      B  , ,  c�����  c����}  d_���}  d_����  c�����      B  , ,  f����  f���}  f����}  f�����  f����      B  , ,  hQ����  hQ���}  h����}  h�����  hQ����      B  , ,  j�����  j����}  kI���}  kI����  j�����      B  , ,  pb����  pb���C  q���C  q����  pb����      B  , ,  r�����  r����C  sZ���C  sZ����  r�����      B  , ,  t�����  t����C  u����C  u�����  t�����      B  , ,  wL����  wL���C  w����C  w�����  wL����      B  , ,  l�����  l����}  m����}  m�����  l�����      B  , ,  o;����  o;���}  o����}  o�����  o;����      B  , ,  q�����  q����}  r3���}  r3����  q�����      B  , ,  s�����  s����}  t����}  t�����  s�����      B  , ,  v%����  v%���}  v����}  v�����  v%����      B  , ,  xs����  xs���}  y���}  y����  xs����      B  , ,  z�����  z����}  {k���}  {k����  z�����      B  , ,  }����  }���}  }����}  }�����  }����      B  , ,  pb���E  pb����  q����  q���E  pb���E      B  , ,  r����E  r�����  sZ����  sZ���E  r����E      B  , ,  t����E  t�����  u�����  u����E  t����E      B  , ,  wL���E  wL����  w�����  w����E  wL���E      B  , ,  ]����  ]���}  ����}  �����  ]����      B  , ,  ������  �����}  �U���}  �U����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �G����  �G���}  �����}  ������  �G����      B  , ,  ������  �����}  �?���}  �?����  ������      B  , ,  pb����  pb����  q����  q����  pb����      B  , ,  r�����  r�����  sZ����  sZ����  r�����      B  , ,  t�����  t�����  u�����  u�����  t�����      B  , ,  pb����  pb����  q����  q����  pb����      B  , ,  r�����  r�����  sZ����  sZ����  r�����      B  , ,  t�����  t�����  u�����  u�����  t�����      B  , ,  wL����  wL����  w�����  w�����  wL����      B  , ,  wL����  wL����  w�����  w�����  wL����      B  , ,  pb����  pb���?  q���?  q����  pb����      B  , ,  r�����  r����?  sZ���?  sZ����  r�����      B  , ,  t�����  t����?  u����?  u�����  t�����      B  , ,  wL����  wL���?  w����?  w�����  wL����      B  , ,  pb����  pb���G  q���G  q����  pb����      B  , ,  r�����  r����G  sZ���G  sZ����  r�����      B  , ,  t�����  t����G  u����G  u�����  t�����      B  , ,  pb����  pb���G  q���G  q����  pb����      B  , ,  r�����  r����G  sZ���G  sZ����  r�����      B  , ,  t�����  t����G  u����G  u�����  t�����      B  , ,  wL����  wL���G  w����G  w�����  wL����      B  , ,  _����  _���a  _����a  _�����  _����      B  , ,  ag����  ag���a  b���a  b����  ag����      B  , ,  c�����  c����a  d_���a  d_����  c�����      B  , ,  f����  f���a  f����a  f�����  f����      B  , ,  hQ����  hQ���a  h����a  h�����  hQ����      B  , ,  j�����  j����a  kI���a  kI����  j�����      B  , ,  l�����  l����a  m����a  m�����  l�����      B  , ,  o;����  o;���a  o����a  o�����  o;����      B  , ,  q�����  q����a  r3���a  r3����  q�����      B  , ,  s�����  s����a  t����a  t�����  s�����      B  , ,  �=����  �=���}  �����}  ������  �=����      B  , ,  ������  �����}  �5���}  �5����  ������      B  , ,  �����A  ������  ������  �����A  �����A      B  , ,  �8���A  �8����  ������  �����A  �8���A      B  , ,  �����A  ������  �0����  �0���A  �����A      B  , ,  �����A  ������  �~����  �~���A  �����A      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  �'����  �'���}  �����}  ������  �'����      B  , ,  �u����  �u���}  ����}  �����  �u����      B  , ,  ������  �����}  �m���}  �m����  ������      B  , ,  �����  ����}  �����}  ������  �����      B  , ,  �_����  �_���}  �	���}  �	����  �_����      B  , ,  ������  �����}  �W���}  �W����  ������      B  , ,  ������  ������  �~����  �~����  ������      B  , ,  �����I  ������  ������  �����I  �����I      B  , ,  �8���I  �8����  ������  �����I  �8���I      B  , ,  �����I  ������  �0����  �0���I  �����I      B  , ,  �����I  ������  �~����  �~���I  �����I      B  , ,  ������  ������  ������  ������  ������      B  , ,  �8����  �8����  ������  ������  �8����      B  , ,  ������  ������  �0����  �0����  ������      B  , ,  ������  ������  �~����  �~����  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �8����  �8����  ������  ������  �8����      B  , ,  ������  ������  �0����  �0����  ������      B  , ,  ������  ������  �~����  �~����  ������      B  , ,  �����E  ������  ������  �����E  �����E      B  , ,  �8���E  �8����  ������  �����E  �8���E      B  , ,  �����E  ������  �0����  �0���E  �����E      B  , ,  �����E  ������  �~����  �~���E  �����E      B  , ,  ������  �����C  �����C  ������  ������      B  , ,  �8����  �8���C  �����C  ������  �8����      B  , ,  ������  �����C  �0���C  �0����  ������      B  , ,  ������  �����C  �~���C  �~����  ������      B  , ,  ������  �����C  �����C  ������  ������      B  , ,  �8����  �8���C  �����C  ������  �8����      B  , ,  ������  �����C  �0���C  �0����  ������      B  , ,  ������  �����C  �~���C  �~����  ������      B  , ,  ������  �����G  �����G  ������  ������      B  , ,  �8����  �8���G  �����G  ������  �8����      B  , ,  ������  �����G  �0���G  �0����  ������      B  , ,  ������  �����G  �~���G  �~����  ������      B  , ,  �����A  ������  ������  �����A  �����A      B  , ,  �8���A  �8����  ������  �����A  �8���A      B  , ,  �����A  ������  �0����  �0���A  �����A      B  , ,  �����A  ������  �~����  �~���A  �����A      B  , ,  ������  �����?  �����?  ������  ������      B  , ,  �8����  �8���?  �����?  ������  �8����      B  , ,  ������  �����?  �0���?  �0����  ������      B  , ,  ������  �����?  �~���?  �~����  ������      B  , ,  �����E  ������  ������  �����E  �����E      B  , ,  �8���E  �8����  ������  �����E  �8���E      B  , ,  �����E  ������  �0����  �0���E  �����E      B  , ,  �����E  ������  �~����  �~���E  �����E      B  , ,  ������  ������  ������  ������  ������      B  , ,  ������  �����a  �����a  ������  ������      B  , ,  �1����  �1���a  �����a  ������  �1����      B  , ,  �����  ����a  �)���a  �)����  �����      B  , ,  ������  �����a  �w���a  �w����  ������      B  , ,  �����  ����a  �����a  ������  �����      B  , ,  �i����  �i���a  ����a  �����  �i����      B  , ,  ������  �����a  �a���a  �a����  ������      B  , ,  �����  ����a  �����a  ������  �����      B  , ,  �S����  �S���a  �����a  ������  �S����      B  , ,  ������  �����a  �K���a  �K����  ������      B  , ,  ������  �����a  �����a  ������  ������      B  , ,  ������  ������  ������  ������  ������      B  , ,  �8����  �8����  ������  ������  �8����      B  , ,  ������  ������  �0����  �0����  ������      B  , ,  ������  ������  �~����  �~����  ������      B  , ,  �=����  �=���a  �����a  ������  �=����      B  , ,  ������  �����a  �5���a  �5����  ������      B  , ,  ������  �����a  �����a  ������  ������      B  , ,  �'����  �'���a  �����a  ������  �'����      B  , ,  �u����  �u���a  ����a  �����  �u����      B  , ,  ������  �����a  �m���a  �m����  ������      B  , ,  �����  ����a  �����a  ������  �����      B  , ,  �_����  �_���a  �	���a  �	����  �_����      B  , ,  ������  �����a  �W���a  �W����  ������      B  , ,  �8����  �8����  ������  ������  �8����      B  , ,  ������  ������  �0����  �0����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  ������  �����G  �����G  ������  ������      B  , ,  �8����  �8���G  �����G  ������  �8����      B  , ,  ������  �����G  �0���G  �0����  ������      B  , ,  ������  �����G  �~���G  �~����  ������      B  , ,  �1����  �1���}  �����}  ������  �1����      B  , ,  �����  ����}  �)���}  �)����  �����      B  , ,  ������  �����}  �w���}  �w����  ������      B  , ,  �����  ����}  �����}  ������  �����      B  , ,  �i����  �i���}  ����}  �����  �i����      B  , ,  ������  �����}  �a���}  �a����  ������      B  , ,  �����  ����}  �����}  ������  �����      B  , ,  �S����  �S���}  �����}  ������  �S����      B  , ,  ������  �����}  �K���}  �K����  ������      B  , ,  ������  �����}  �����}  ������  ������      B  , ,  ����}�  ����~s  �H��~s  �H��}�  ����}�      B  , ,  ����|  ����|�  �H��|�  �H��|  ����|      B  , ,  �����I  ������  �0����  �0���I  �����I      B  , ,  �����I  ������  �~����  �~���I  �����I      B  , ,  ������  ������  ������  ������  ������      B  , ,  �8����  �8����  ������  ������  �8����      B  , ,  ������  ������  �0����  �0����  ������      B  , ,  ������  ������  �~����  �~����  ������      B  , ,  �����I  ������  ������  �����I  �����I      B  , ,  ����}�  ����~s  �0��~s  �0��}�  ����}�      B  , ,  ����}�  ����~s  ����~s  ����}�  ����}�      B  , ,  �.��}�  �.��~s  ����~s  ����}�  �.��}�      B  , ,  ����}�  ����~s  �,��~s  �,��}�  ����}�      B  , ,  ����}�  ����~s  ����~s  ����}�  ����}�      B  , ,  �*��}�  �*��~s  ����~s  ����}�  �*��}�      B  , ,  �~��}�  �~��~s  �(��~s  �(��}�  �~��}�      B  , ,  ����}�  ����~s  �|��~s  �|��}�  ����}�      B  , ,  �&��}�  �&��~s  ����~s  ����}�  �&��}�      B  , ,  �z��}�  �z��~s  �$��~s  �$��}�  �z��}�      B  , ,  ����}�  ����~s  �x��~s  �x��}�  ����}�      B  , ,  �"��}�  �"��~s  ����~s  ����}�  �"��}�      B  , ,  �v��}�  �v��~s  � ��~s  � ��}�  �v��}�      B  , ,  ����}�  ����~s  �t��~s  �t��}�  ����}�      B  , ,  ���}�  ���~s  ����~s  ����}�  ���}�      B  , ,  �r��}�  �r��~s  ���~s  ���}�  �r��}�      B  , ,  ����}�  ����~s  �p��~s  �p��}�  ����}�      B  , ,  �8���I  �8����  ������  �����I  �8���I      B  , ,  ����|  ����|�  �0��|�  �0��|  ����|      B  , ,  ����|  ����|�  ����|�  ����|  ����|      B  , ,  �.��|  �.��|�  ����|�  ����|  �.��|      B  , ,  ����|  ����|�  �,��|�  �,��|  ����|      B  , ,  ����|  ����|�  ����|�  ����|  ����|      B  , ,  �*��|  �*��|�  ����|�  ����|  �*��|      B  , ,  �~��|  �~��|�  �(��|�  �(��|  �~��|      B  , ,  ����|  ����|�  �|��|�  �|��|  ����|      B  , ,  �&��|  �&��|�  ����|�  ����|  �&��|      B  , ,  �z��|  �z��|�  �$��|�  �$��|  �z��|      B  , ,  ����|  ����|�  �x��|�  �x��|  ����|      B  , ,  �"��|  �"��|�  ����|�  ����|  �"��|      B  , ,  �v��|  �v��|�  � ��|�  � ��|  �v��|      B  , ,  ����|  ����|�  �t��|�  �t��|  ����|      B  , ,  ���|  ���|�  ����|�  ����|  ���|      B  , ,  �r��|  �r��|�  ���|�  ���|  �r��|      B  , ,  ����|  ����|�  �p��|�  �p��|  ����|      B  , ,  ����|  ����|�  ����|�  ����|  ����|      B  , ,  �F��|  �F��|�  ����|�  ����|  �F��|      B  , ,  ����|  ����|�  �D��|�  �D��|  ����|      B  , ,  ����|  ����|�  ����|�  ����|  ����|      B  , ,  �B��|  �B��|�  ����|�  ����|  �B��|      B  , ,  ����|  ����|�  �@��|�  �@��|  ����|      B  , ,  ����|  ����|�  ����|�  ����|  ����|      B  , ,  �>��|  �>��|�  ����|�  ����|  �>��|      B  , ,  ����|  ����|�  �<��|�  �<��|  ����|      B  , ,  ����|  ����|�  ����|�  ����|  ����|      B  , ,  �:��|  �:��|�  ����|�  ����|  �:��|      B  , ,  ����|  ����|�  �8��|�  �8��|  ����|      B  , ,  ����|  ����|�  ����|�  ����|  ����|      B  , ,  �6��|  �6��|�  ����|�  ����|  �6��|      B  , ,  ����|  ����|�  �4��|�  �4��|  ����|      B  , ,  ����|  ����|�  ����|�  ����|  ����|      B  , ,  �2��|  �2��|�  ����|�  ����|  �2��|      B  , ,  �F��}�  �F��~s  ����~s  ����}�  �F��}�      B  , ,  ����}�  ����~s  �D��~s  �D��}�  ����}�      B  , ,  ����}�  ����~s  ����~s  ����}�  ����}�      B  , ,  �B��}�  �B��~s  ����~s  ����}�  �B��}�      B  , ,  ����}�  ����~s  �@��~s  �@��}�  ����}�      B  , ,  ����}�  ����~s  ����~s  ����}�  ����}�      B  , ,  �>��}�  �>��~s  ����~s  ����}�  �>��}�      B  , ,  ����}�  ����~s  �<��~s  �<��}�  ����}�      B  , ,  ����}�  ����~s  ����~s  ����}�  ����}�      B  , ,  �:��}�  �:��~s  ����~s  ����}�  �:��}�      B  , ,  ����}�  ����~s  �8��~s  �8��}�  ����}�      B  , ,  ����}�  ����~s  ����~s  ����}�  ����}�      B  , ,  �6��}�  �6��~s  ����~s  ����}�  �6��}�      B  , ,  ����}�  ����~s  �4��~s  �4��}�  ����}�      B  , ,  ����}�  ����~s  ����~s  ����}�  ����}�      B  , ,  �2��}�  �2��~s  ����~s  ����}�  �2��}�      B  , ,  ����}�  ����~s  ����~s  ����}�  ����}�      B  , ,  ����q�  ����rp  �t��rp  �t��q�  ����q�      B  , ,  ���q�  ���rp  ����rp  ����q�  ���q�      B  , ,  �f��q�  �f��rp  ���rp  ���q�  �f��q�      B  , ,  ����q�  ����rp  �^��rp  �^��q�  ����q�      B  , ,  ����pr  ����q  �t��q  �t��pr  ����pr      B  , ,  ���pr  ���q  ����q  ����pr  ���pr      B  , ,  �f��pr  �f��q  ���q  ���pr  �f��pr      B  , ,  ����pr  ����q  �^��q  �^��pr  ����pr      B  , ,  ����o  ����o�  �t��o�  �t��o  ����o      B  , ,  ���o  ���o�  ����o�  ����o  ���o      B  , ,  �f��o  �f��o�  ���o�  ���o  �f��o      B  , ,  ����o  ����o�  �^��o�  �^��o  ����o      B  , ,  ����m�  ����nt  �t��nt  �t��m�  ����m�      B  , ,  ���m�  ���nt  ����nt  ����m�  ���m�      B  , ,  �f��m�  �f��nt  ���nt  ���m�  �f��m�      B  , ,  ����m�  ����nt  �^��nt  �^��m�  ����m�      B  , ,  ����lv  ����m   �t��m   �t��lv  ����lv      B  , ,  ���lv  ���m   ����m   ����lv  ���lv      B  , ,  �f��lv  �f��m   ���m   ���lv  �f��lv      B  , ,  ����lv  ����m   �^��m   �^��lv  ����lv      B  , ,  ����k"  ����k�  �t��k�  �t��k"  ����k"      B  , ,  ���k"  ���k�  ����k�  ����k"  ���k"      B  , ,  �f��k"  �f��k�  ���k�  ���k"  �f��k"      B  , ,  ����k"  ����k�  �^��k�  �^��k"  ����k"      B  , ,  ����i�  ����jx  �t��jx  �t��i�  ����i�      B  , ,  ���i�  ���jx  ����jx  ����i�  ���i�      B  , ,  �f��i�  �f��jx  ���jx  ���i�  �f��i�      B  , ,  ����i�  ����jx  �^��jx  �^��i�  ����i�      B  , ,  �:��q�  �:��rp  ����rp  ����q�  �:��q�      B  , ,  ����q�  ����rp  �2��rp  �2��q�  ����q�      B  , ,  ����q�  ����rp  ����rp  ����q�  ����q�      B  , ,  �$��q�  �$��rp  ����rp  ����q�  �$��q�      B  , ,  ���o  ���o�  ����o�  ����o  ���o      B  , ,  �P��o  �P��o�  ����o�  ����o  �P��o      B  , ,  ����o  ����o�  �H��o�  �H��o  ����o      B  , ,  ����o  ����o�  ����o�  ����o  ����o      B  , ,  �:��o  �:��o�  ����o�  ����o  �:��o      B  , ,  ����o  ����o�  �2��o�  �2��o  ����o      B  , ,  ����o  ����o�  ����o�  ����o  ����o      B  , ,  �$��o  �$��o�  ����o�  ����o  �$��o      B  , ,  �r��o  �r��o�  ���o�  ���o  �r��o      B  , ,  ����o  ����o�  �j��o�  �j��o  ����o      B  , ,  �r��q�  �r��rp  ���rp  ���q�  �r��q�      B  , ,  ����q�  ����rp  �j��rp  �j��q�  ����q�      B  , ,  ���q�  ���rp  ����rp  ����q�  ���q�      B  , ,  �P��q�  �P��rp  ����rp  ����q�  �P��q�      B  , ,  ���m�  ���nt  ����nt  ����m�  ���m�      B  , ,  �P��m�  �P��nt  ����nt  ����m�  �P��m�      B  , ,  ����m�  ����nt  �H��nt  �H��m�  ����m�      B  , ,  ����m�  ����nt  ����nt  ����m�  ����m�      B  , ,  �:��m�  �:��nt  ����nt  ����m�  �:��m�      B  , ,  ����m�  ����nt  �2��nt  �2��m�  ����m�      B  , ,  ����m�  ����nt  ����nt  ����m�  ����m�      B  , ,  �$��m�  �$��nt  ����nt  ����m�  �$��m�      B  , ,  �r��m�  �r��nt  ���nt  ���m�  �r��m�      B  , ,  ����m�  ����nt  �j��nt  �j��m�  ����m�      B  , ,  ����q�  ����rp  �H��rp  �H��q�  ����q�      B  , ,  ����q�  ����rp  ����rp  ����q�  ����q�      B  , ,  ���pr  ���q  ����q  ����pr  ���pr      B  , ,  �P��pr  �P��q  ����q  ����pr  �P��pr      B  , ,  ���lv  ���m   ����m   ����lv  ���lv      B  , ,  �P��lv  �P��m   ����m   ����lv  �P��lv      B  , ,  ����lv  ����m   �H��m   �H��lv  ����lv      B  , ,  ����lv  ����m   ����m   ����lv  ����lv      B  , ,  �:��lv  �:��m   ����m   ����lv  �:��lv      B  , ,  ����lv  ����m   �2��m   �2��lv  ����lv      B  , ,  ����lv  ����m   ����m   ����lv  ����lv      B  , ,  �$��lv  �$��m   ����m   ����lv  �$��lv      B  , ,  �r��lv  �r��m   ���m   ���lv  �r��lv      B  , ,  ����lv  ����m   �j��m   �j��lv  ����lv      B  , ,  ����pr  ����q  �H��q  �H��pr  ����pr      B  , ,  ����pr  ����q  ����q  ����pr  ����pr      B  , ,  �:��pr  �:��q  ����q  ����pr  �:��pr      B  , ,  ����pr  ����q  �2��q  �2��pr  ����pr      B  , ,  ���k"  ���k�  ����k�  ����k"  ���k"      B  , ,  �P��k"  �P��k�  ����k�  ����k"  �P��k"      B  , ,  ����k"  ����k�  �H��k�  �H��k"  ����k"      B  , ,  ����k"  ����k�  ����k�  ����k"  ����k"      B  , ,  �:��k"  �:��k�  ����k�  ����k"  �:��k"      B  , ,  ����k"  ����k�  �2��k�  �2��k"  ����k"      B  , ,  ����k"  ����k�  ����k�  ����k"  ����k"      B  , ,  �$��k"  �$��k�  ����k�  ����k"  �$��k"      B  , ,  �r��k"  �r��k�  ���k�  ���k"  �r��k"      B  , ,  ����k"  ����k�  �j��k�  �j��k"  ����k"      B  , ,  ����pr  ����q  ����q  ����pr  ����pr      B  , ,  �$��pr  �$��q  ����q  ����pr  �$��pr      B  , ,  �r��pr  �r��q  ���q  ���pr  �r��pr      B  , ,  ����pr  ����q  �j��q  �j��pr  ����pr      B  , ,  ���i�  ���jx  ����jx  ����i�  ���i�      B  , ,  �P��i�  �P��jx  ����jx  ����i�  �P��i�      B  , ,  ����i�  ����jx  �H��jx  �H��i�  ����i�      B  , ,  ����i�  ����jx  ����jx  ����i�  ����i�      B  , ,  �:��i�  �:��jx  ����jx  ����i�  �:��i�      B  , ,  ����i�  ����jx  �2��jx  �2��i�  ����i�      B  , ,  ����i�  ����jx  ����jx  ����i�  ����i�      B  , ,  �$��i�  �$��jx  ����jx  ����i�  �$��i�      B  , ,  �r��i�  �r��jx  ���jx  ���i�  �r��i�      B  , ,  ����i�  ����jx  �j��jx  �j��i�  ����i�      B  , ,  r�����  r�����  sZ����  sZ����  r�����      B  , ,  r����I  r�����  sZ����  sZ���I  r����I      B  , ,  u���|  u���|�  v\��|�  v\��|  u���|      B  , ,  w��|  w��|�  w���|�  w���|  w��|      B  , ,  xZ��|  xZ��|�  y��|�  y��|  xZ��|      B  , ,  y���|  y���|�  zX��|�  zX��|  y���|      B  , ,  {��|  {��|�  {���|�  {���|  {��|      B  , ,  |V��|  |V��|�  } ��|�  } ��|  |V��|      B  , ,  }���|  }���|�  ~T��|�  ~T��|  }���|      B  , ,  ~���|  ~���|�  ���|�  ���|  ~���|      B  , ,  �R��|  �R��|�  ����|�  ����|  �R��|      B  , ,  ����|  ����|�  �P��|�  �P��|  ����|      B  , ,  ����|  ����|�  ����|�  ����|  ����|      B  , ,  �N��|  �N��|�  ����|�  ����|  �N��|      B  , ,  ����|  ����|�  �L��|�  �L��|  ����|      B  , ,  ����|  ����|�  ����|�  ����|  ����|      B  , ,  �J��|  �J��|�  ����|�  ����|  �J��|      B  , ,  �N��}�  �N��~s  ����~s  ����}�  �N��}�      B  , ,  ����}�  ����~s  �L��~s  �L��}�  ����}�      B  , ,  ����}�  ����~s  ����~s  ����}�  ����}�      B  , ,  �J��}�  �J��~s  ����~s  ����}�  �J��}�      B  , ,  t�����  t�����  u�����  u�����  t�����      B  , ,  wL����  wL����  w�����  w�����  wL����      B  , ,  t����I  t�����  u�����  u����I  t����I      B  , ,  wL���I  wL����  w�����  w����I  wL���I      B  , ,  s
��|  s
��|�  s���|�  s���|  s
��|      B  , ,  s
��}�  s
��~s  s���~s  s���}�  s
��}�      B  , ,  t^��}�  t^��~s  u��~s  u��}�  t^��}�      B  , ,  u���}�  u���~s  v\��~s  v\��}�  u���}�      B  , ,  w��}�  w��~s  w���~s  w���}�  w��}�      B  , ,  xZ��}�  xZ��~s  y��~s  y��}�  xZ��}�      B  , ,  y���}�  y���~s  zX��~s  zX��}�  y���}�      B  , ,  {��}�  {��~s  {���~s  {���}�  {��}�      B  , ,  |V��}�  |V��~s  } ��~s  } ��}�  |V��}�      B  , ,  }���}�  }���~s  ~T��~s  ~T��}�  }���}�      B  , ,  t^��|  t^��|�  u��|�  u��|  t^��|      B  , ,  ~���}�  ~���~s  ���~s  ���}�  ~���}�      B  , ,  �R��}�  �R��~s  ����~s  ����}�  �R��}�      B  , ,  ����}�  ����~s  �P��~s  �P��}�  ����}�      B  , ,  ����}�  ����~s  ����~s  ����}�  ����}�      B  , ,  hj��}�  hj��~s  i��~s  i��}�  hj��}�      B  , ,  i���}�  i���~s  jh��~s  jh��}�  i���}�      B  , ,  k��}�  k��~s  k���~s  k���}�  k��}�      B  , ,  lf��}�  lf��~s  m��~s  m��}�  lf��}�      B  , ,  m���}�  m���~s  nd��~s  nd��}�  m���}�      B  , ,  o��}�  o��~s  o���~s  o���}�  o��}�      B  , ,  pb��}�  pb��~s  q��~s  q��}�  pb��}�      B  , ,  q���}�  q���~s  r`��~s  r`��}�  q���}�      B  , ,  m���|  m���|�  nd��|�  nd��|  m���|      B  , ,  o��|  o��|�  o���|�  o���|  o��|      B  , ,  pb��|  pb��|�  q��|�  q��|  pb��|      B  , ,  q���|  q���|�  r`��|�  r`��|  q���|      B  , ,  pb����  pb����  q����  q����  pb����      B  , ,  lf��|  lf��|�  m��|�  m��|  lf��|      B  , ,  ]���}�  ]���~s  ^t��~s  ^t��}�  ]���}�      B  , ,  _��}�  _��~s  _���~s  _���}�  _��}�      B  , ,  `r��}�  `r��~s  a��~s  a��}�  `r��}�      B  , ,  a���}�  a���~s  bp��~s  bp��}�  a���}�      B  , ,  c��}�  c��~s  c���~s  c���}�  c��}�      B  , ,  dn��}�  dn��~s  e��~s  e��}�  dn��}�      B  , ,  e���}�  e���~s  fl��~s  fl��}�  e���}�      B  , ,  g��}�  g��~s  g���~s  g���}�  g��}�      B  , ,  pb���I  pb����  q����  q���I  pb���I      B  , ,  ]���|  ]���|�  ^t��|�  ^t��|  ]���|      B  , ,  _��|  _��|�  _���|�  _���|  _��|      B  , ,  `r��|  `r��|�  a��|�  a��|  `r��|      B  , ,  a���|  a���|�  bp��|�  bp��|  a���|      B  , ,  c��|  c��|�  c���|�  c���|  c��|      B  , ,  dn��|  dn��|�  e��|�  e��|  dn��|      B  , ,  e���|  e���|�  fl��|�  fl��|  e���|      B  , ,  g��|  g��|�  g���|�  g���|  g��|      B  , ,  hj��|  hj��|�  i��|�  i��|  hj��|      B  , ,  i���|  i���|�  jh��|�  jh��|  i���|      B  , ,  k��|  k��|�  k���|�  k���|  k��|      B  , ,  {���q�  {���rp  |���rp  |���q�  {���q�      B  , ,  ~J��q�  ~J��rp  ~���rp  ~���q�  ~J��q�      B  , ,  ����q�  ����rp  �B��rp  �B��q�  ����q�      B  , ,  ����q�  ����rp  ����rp  ����q�  ����q�      B  , ,  {���m�  {���nt  |���nt  |���m�  {���m�      B  , ,  ~J��m�  ~J��nt  ~���nt  ~���m�  ~J��m�      B  , ,  {���lv  {���m   |���m   |���lv  {���lv      B  , ,  ~J��lv  ~J��m   ~���m   ~���lv  ~J��lv      B  , ,  ����lv  ����m   �B��m   �B��lv  ����lv      B  , ,  ����lv  ����m   ����m   ����lv  ����lv      B  , ,  {���i�  {���jx  |���jx  |���i�  {���i�      B  , ,  ~J��i�  ~J��jx  ~���jx  ~���i�  ~J��i�      B  , ,  ����i�  ����jx  �B��jx  �B��i�  ����i�      B  , ,  ����i�  ����jx  ����jx  ����i�  ����i�      B  , ,  ����m�  ����nt  �B��nt  �B��m�  ����m�      B  , ,  ����m�  ����nt  ����nt  ����m�  ����m�      B  , ,  {���k"  {���k�  |���k�  |���k"  {���k"      B  , ,  ~J��k"  ~J��k�  ~���k�  ~���k"  ~J��k"      B  , ,  ����k"  ����k�  �B��k�  �B��k"  ����k"      B  , ,  ����k"  ����k�  ����k�  ����k"  ����k"      B  , ,  ����o  ����o�  �B��o�  �B��o  ����o      B  , ,  ����o  ����o�  ����o�  ����o  ����o      B  , ,  {���pr  {���q  |���q  |���pr  {���pr      B  , ,  ~J��pr  ~J��q  ~���q  ~���pr  ~J��pr      B  , ,  ����pr  ����q  �B��q  �B��pr  ����pr      B  , ,  ����pr  ����q  ����q  ����pr  ����pr      B  , ,  {���o  {���o�  |���o�  |���o  {���o      B  , ,  ~J��o  ~J��o�  ~���o�  ~���o  ~J��o      B  , ,  {���hz  {���i$  |���i$  |���hz  {���hz      B  , ,  ~J��hz  ~J��i$  ~���i$  ~���hz  ~J��hz      B  , ,  ����hz  ����i$  �B��i$  �B��hz  ����hz      B  , ,  ����hz  ����i$  ����i$  ����hz  ����hz      B  , ,  s���f1  s���f�  t���f�  t���f1  s���f1      B  , ,  v9��f1  v9��f�  v���f�  v���f1  v9��f1      B  , ,  x���f1  x���f�  y1��f�  y1��f1  x���f1      B  , ,  z���f1  z���f�  {��f�  {��f1  z���f1      B  , ,  }#��f1  }#��f�  }���f�  }���f1  }#��f1      B  , ,  q��f1  q��f�  ���f�  ���f1  q��f1      B  , ,  ����f1  ����f�  �i��f�  �i��f1  ����f1      B  , ,  ���f1  ���f�  ����f�  ����f1  ���f1      B  , ,  �[��f1  �[��f�  ���f�  ���f1  �[��f1      B  , ,  ����f1  ����f�  �S��f�  �S��f1  ����f1      B  , ,  s���d  s���d�  t���d�  t���d  s���d      B  , ,  v9��d  v9��d�  v���d�  v���d  v9��d      B  , ,  x���d  x���d�  y1��d�  y1��d  x���d      B  , ,  z���d  z���d�  {��d�  {��d  z���d      B  , ,  }#��d  }#��d�  }���d�  }���d  }#��d      B  , ,  q��d  q��d�  ���d�  ���d  q��d      B  , ,  ����d  ����d�  �i��d�  �i��d  ����d      B  , ,  ���d  ���d�  ����d�  ����d  ���d      B  , ,  �[��d  �[��d�  ���d�  ���d  �[��d      B  , ,  ����d  ����d�  �S��d�  �S��d  ����d      B  , ,  {���a�  {���bv  |���bv  |���a�  {���a�      B  , ,  ~J��a�  ~J��bv  ~���bv  ~���a�  ~J��a�      B  , ,  ����a�  ����bv  �B��bv  �B��a�  ����a�      B  , ,  ����a�  ����bv  ����bv  ����a�  ����a�      B  , ,  {���`x  {���a"  |���a"  |���`x  {���`x      B  , ,  ~J��`x  ~J��a"  ~���a"  ~���`x  ~J��`x      B  , ,  ����`x  ����a"  �B��a"  �B��`x  ����`x      B  , ,  ����`x  ����a"  ����a"  ����`x  ����`x      B  , ,  {���_$  {���_�  |���_�  |���_$  {���_$      B  , ,  ~J��_$  ~J��_�  ~���_�  ~���_$  ~J��_$      B  , ,  ����_$  ����_�  �B��_�  �B��_$  ����_$      B  , ,  ����_$  ����_�  ����_�  ����_$  ����_$      B  , ,  {���]�  {���^z  |���^z  |���]�  {���]�      B  , ,  ~J��]�  ~J��^z  ~���^z  ~���]�  ~J��]�      B  , ,  ����]�  ����^z  �B��^z  �B��]�  ����]�      B  , ,  ����]�  ����^z  ����^z  ����]�  ����]�      B  , ,  {���\|  {���]&  |���]&  |���\|  {���\|      B  , ,  ~J��\|  ~J��]&  ~���]&  ~���\|  ~J��\|      B  , ,  ����\|  ����]&  �B��]&  �B��\|  ����\|      B  , ,  ����\|  ����]&  ����]&  ����\|  ����\|      B  , ,  {���[(  {���[�  |���[�  |���[(  {���[(      B  , ,  ~J��[(  ~J��[�  ~���[�  ~���[(  ~J��[(      B  , ,  ����[(  ����[�  �B��[�  �B��[(  ����[(      B  , ,  ����[(  ����[�  ����[�  ����[(  ����[(      B  , ,  {���Y�  {���Z~  |���Z~  |���Y�  {���Y�      B  , ,  ~J��Y�  ~J��Z~  ~���Z~  ~���Y�  ~J��Y�      B  , ,  ����Y�  ����Z~  �B��Z~  �B��Y�  ����Y�      B  , ,  ����Y�  ����Z~  ����Z~  ����Y�  ����Y�      B  , ,  {���X�  {���Y*  |���Y*  |���X�  {���X�      B  , ,  ~J��X�  ~J��Y*  ~���Y*  ~���X�  ~J��X�      B  , ,  ����X�  ����Y*  �B��Y*  �B��X�  ����X�      B  , ,  ����X�  ����Y*  ����Y*  ����X�  ����X�      B  , ,  ���a�  ���bv  ����bv  ����a�  ���a�      B  , ,  �P��a�  �P��bv  ����bv  ����a�  �P��a�      B  , ,  ����a�  ����bv  �H��bv  �H��a�  ����a�      B  , ,  ����a�  ����bv  ����bv  ����a�  ����a�      B  , ,  �:��a�  �:��bv  ����bv  ����a�  �:��a�      B  , ,  ����a�  ����bv  �2��bv  �2��a�  ����a�      B  , ,  ����a�  ����bv  ����bv  ����a�  ����a�      B  , ,  �$��a�  �$��bv  ����bv  ����a�  �$��a�      B  , ,  �r��a�  �r��bv  ���bv  ���a�  �r��a�      B  , ,  ����a�  ����bv  �j��bv  �j��a�  ����a�      B  , ,  ���`x  ���a"  ����a"  ����`x  ���`x      B  , ,  �P��`x  �P��a"  ����a"  ����`x  �P��`x      B  , ,  ����`x  ����a"  �H��a"  �H��`x  ����`x      B  , ,  ����`x  ����a"  ����a"  ����`x  ����`x      B  , ,  �:��`x  �:��a"  ����a"  ����`x  �:��`x      B  , ,  ����`x  ����a"  �2��a"  �2��`x  ����`x      B  , ,  ����`x  ����a"  ����a"  ����`x  ����`x      B  , ,  �$��`x  �$��a"  ����a"  ����`x  �$��`x      B  , ,  �r��`x  �r��a"  ���a"  ���`x  �r��`x      B  , ,  ����`x  ����a"  �j��a"  �j��`x  ����`x      B  , ,  ����hz  ����i$  ����i$  ����hz  ����hz      B  , ,  �$��hz  �$��i$  ����i$  ����hz  �$��hz      B  , ,  �r��hz  �r��i$  ���i$  ���hz  �r��hz      B  , ,  ���_$  ���_�  ����_�  ����_$  ���_$      B  , ,  �P��_$  �P��_�  ����_�  ����_$  �P��_$      B  , ,  ����_$  ����_�  �H��_�  �H��_$  ����_$      B  , ,  ����_$  ����_�  ����_�  ����_$  ����_$      B  , ,  �:��_$  �:��_�  ����_�  ����_$  �:��_$      B  , ,  ����_$  ����_�  �2��_�  �2��_$  ����_$      B  , ,  ����_$  ����_�  ����_�  ����_$  ����_$      B  , ,  �$��_$  �$��_�  ����_�  ����_$  �$��_$      B  , ,  �r��_$  �r��_�  ���_�  ���_$  �r��_$      B  , ,  ����_$  ����_�  �j��_�  �j��_$  ����_$      B  , ,  ����hz  ����i$  �j��i$  �j��hz  ����hz      B  , ,  ���]�  ���^z  ����^z  ����]�  ���]�      B  , ,  �P��]�  �P��^z  ����^z  ����]�  �P��]�      B  , ,  ����]�  ����^z  �H��^z  �H��]�  ����]�      B  , ,  ����]�  ����^z  ����^z  ����]�  ����]�      B  , ,  �:��]�  �:��^z  ����^z  ����]�  �:��]�      B  , ,  ����]�  ����^z  �2��^z  �2��]�  ����]�      B  , ,  ����]�  ����^z  ����^z  ����]�  ����]�      B  , ,  �$��]�  �$��^z  ����^z  ����]�  �$��]�      B  , ,  �r��]�  �r��^z  ���^z  ���]�  �r��]�      B  , ,  ����]�  ����^z  �j��^z  �j��]�  ����]�      B  , ,  ���hz  ���i$  ����i$  ����hz  ���hz      B  , ,  �P��hz  �P��i$  ����i$  ����hz  �P��hz      B  , ,  ���\|  ���]&  ����]&  ����\|  ���\|      B  , ,  �P��\|  �P��]&  ����]&  ����\|  �P��\|      B  , ,  ����\|  ����]&  �H��]&  �H��\|  ����\|      B  , ,  ����\|  ����]&  ����]&  ����\|  ����\|      B  , ,  �:��\|  �:��]&  ����]&  ����\|  �:��\|      B  , ,  ����\|  ����]&  �2��]&  �2��\|  ����\|      B  , ,  ����\|  ����]&  ����]&  ����\|  ����\|      B  , ,  �$��\|  �$��]&  ����]&  ����\|  �$��\|      B  , ,  �r��\|  �r��]&  ���]&  ���\|  �r��\|      B  , ,  ����\|  ����]&  �j��]&  �j��\|  ����\|      B  , ,  ���[(  ���[�  ����[�  ����[(  ���[(      B  , ,  �P��[(  �P��[�  ����[�  ����[(  �P��[(      B  , ,  ����[(  ����[�  �H��[�  �H��[(  ����[(      B  , ,  ����[(  ����[�  ����[�  ����[(  ����[(      B  , ,  �:��[(  �:��[�  ����[�  ����[(  �:��[(      B  , ,  ����[(  ����[�  �2��[�  �2��[(  ����[(      B  , ,  ����[(  ����[�  ����[�  ����[(  ����[(      B  , ,  �$��[(  �$��[�  ����[�  ����[(  �$��[(      B  , ,  �r��[(  �r��[�  ���[�  ���[(  �r��[(      B  , ,  ����[(  ����[�  �j��[�  �j��[(  ����[(      B  , ,  ����hz  ����i$  �H��i$  �H��hz  ����hz      B  , ,  ����hz  ����i$  ����i$  ����hz  ����hz      B  , ,  �:��hz  �:��i$  ����i$  ����hz  �:��hz      B  , ,  ����hz  ����i$  �2��i$  �2��hz  ����hz      B  , ,  �f��\|  �f��]&  ���]&  ���\|  �f��\|      B  , ,  ����\|  ����]&  �^��]&  �^��\|  ����\|      B  , ,  ���_$  ���_�  ����_�  ����_$  ���_$      B  , ,  ����hz  ����i$  �t��i$  �t��hz  ����hz      B  , ,  ���hz  ���i$  ����i$  ����hz  ���hz      B  , ,  �f��hz  �f��i$  ���i$  ���hz  �f��hz      B  , ,  ����]�  ����^z  �t��^z  �t��]�  ����]�      B  , ,  ���]�  ���^z  ����^z  ����]�  ���]�      B  , ,  �f��]�  �f��^z  ���^z  ���]�  �f��]�      B  , ,  ����]�  ����^z  �^��^z  �^��]�  ����]�      B  , ,  �f��_$  �f��_�  ���_�  ���_$  �f��_$      B  , ,  ����_$  ����_�  �^��_�  �^��_$  ����_$      B  , ,  �E��d  �E��d�  ����d�  ����d  �E��d      B  , ,  ����d  ����d�  �=��d�  �=��d  ����d      B  , ,  ����d  ����d�  ����d�  ����d  ����d      B  , ,  �/��d  �/��d�  ����d�  ����d  �/��d      B  , ,  ����[(  ����[�  �t��[�  �t��[(  ����[(      B  , ,  ���[(  ���[�  ����[�  ����[(  ���[(      B  , ,  �f��[(  �f��[�  ���[�  ���[(  �f��[(      B  , ,  ����[(  ����[�  �^��[�  �^��[(  ����[(      B  , ,  ���`x  ���a"  ����a"  ����`x  ���`x      B  , ,  �f��`x  �f��a"  ���a"  ���`x  �f��`x      B  , ,  ����`x  ����a"  �^��a"  �^��`x  ����`x      B  , ,  ����f1  ����f�  ����f�  ����f1  ����f1      B  , ,  �E��f1  �E��f�  ����f�  ����f1  �E��f1      B  , ,  �/��f1  �/��f�  ����f�  ����f1  �/��f1      B  , ,  ����f1  ����f�  �=��f�  �=��f1  ����f1      B  , ,  ����f1  ����f�  ����f�  ����f1  ����f1      B  , ,  ����hz  ����i$  �^��i$  �^��hz  ����hz      B  , ,  ����`x  ����a"  �t��a"  �t��`x  ����`x      B  , ,  ����_$  ����_�  �t��_�  �t��_$  ����_$      B  , ,  ����d  ����d�  ����d�  ����d  ����d      B  , ,  ����\|  ����]&  �t��]&  �t��\|  ����\|      B  , ,  ���\|  ���]&  ����]&  ����\|  ���\|      B  , ,  ����a�  ����bv  �t��bv  �t��a�  ����a�      B  , ,  ���a�  ���bv  ����bv  ����a�  ���a�      B  , ,  �f��a�  �f��bv  ���bv  ���a�  �f��a�      B  , ,  ����a�  ����bv  �^��bv  �^��a�  ����a�      B  , ,  ����Y�  ����Z~  �t��Z~  �t��Y�  ����Y�      B  , ,  ���Y�  ���Z~  ����Z~  ����Y�  ���Y�      B  , ,  �f��Y�  �f��Z~  ���Z~  ���Y�  �f��Y�      B  , ,  ����Y�  ����Z~  �^��Z~  �^��Y�  ����Y�      B  , ,  ����X�  ����Y*  �t��Y*  �t��X�  ����X�      B  , ,  ���X�  ���Y*  ����Y*  ����X�  ���X�      B  , ,  �f��X�  �f��Y*  ���Y*  ���X�  �f��X�      B  , ,  ����X�  ����Y*  �^��Y*  �^��X�  ����X�      B  , ,  �r��Y�  �r��Z~  ���Z~  ���Y�  �r��Y�      B  , ,  ����Y�  ����Z~  �j��Z~  �j��Y�  ����Y�      B  , ,  ���Y�  ���Z~  ����Z~  ����Y�  ���Y�      B  , ,  �P��Y�  �P��Z~  ����Z~  ����Y�  �P��Y�      B  , ,  ����Y�  ����Z~  �H��Z~  �H��Y�  ����Y�      B  , ,  ����Y�  ����Z~  ����Z~  ����Y�  ����Y�      B  , ,  �:��Y�  �:��Z~  ����Z~  ����Y�  �:��Y�      B  , ,  ����Y�  ����Z~  �2��Z~  �2��Y�  ����Y�      B  , ,  ����Y�  ����Z~  ����Z~  ����Y�  ����Y�      B  , ,  �$��Y�  �$��Z~  ����Z~  ����Y�  �$��Y�      B  , ,  ���X�  ���Y*  ����Y*  ����X�  ���X�      B  , ,  �P��X�  �P��Y*  ����Y*  ����X�  �P��X�      B  , ,  ����X�  ����Y*  �H��Y*  �H��X�  ����X�      B  , ,  ����X�  ����Y*  ����Y*  ����X�  ����X�      B  , ,  �:��X�  �:��Y*  ����Y*  ����X�  �:��X�      B  , ,  ����X�  ����Y*  �2��Y*  �2��X�  ����X�      B  , ,  ����X�  ����Y*  ����Y*  ����X�  ����X�      B  , ,  �$��X�  �$��Y*  ����Y*  ����X�  �$��X�      B  , ,  �r��X�  �r��Y*  ���Y*  ���X�  �r��X�      B  , ,  ����X�  ����Y*  �j��Y*  �j��X�  ����X�      B  , , ���h� ���i� ���i� ���h� ���h�      B  , , ���h� ���i� |��i� |��h� ���h�      B  , , ���h� ���i� `��i� `��h� ���h�      B  , , ���h� ���i� D��i� D��h� ���h�      B  , , ���o� ���p, ���p, ���o� ���o�      B  , , ���o� ���p, |��p, |��o� ���o�      B  , , ���o� ���p, `��p, `��o� ���o�      B  , , ���o� ���p, D��p, D��o� ���o�      B  , , ���j2 ���j� ���j� ���j2 ���j2      B  , , ���j2 ���j� |��j� |��j2 ���j2      B  , , ���j2 ���j� `��j� `��j2 ���j2      B  , , ���j2 ���j� D��j� D��j2 ���j2      B  , , ���k� ���l0 ���l0 ���k� ���k�      B  , , ���k� ���l0 |��l0 |��k� ���k�      B  , , ���k� ���l0 `��l0 `��k� ���k�      B  , , ���k� ���l0 D��l0 D��k� ���k�      B  , , ���n. ���n� ���n� ���n. ���n.      B  , , ���n. ���n� |��n� |��n. ���n.      B  , , ���n. ���n� `��n� `��n. ���n.      B  , , ���n. ���n� D��n� D��n. ���n.      B  , , ���r* ���r� ���r� ���r* ���r*      B  , , ���r* ���r� |��r� |��r* ���r*      B  , , ���r* ���r� `��r� `��r* ���r*      B  , , ���r* ���r� D��r� D��r* ���r*      B  , , ���l� ���m� ���m� ���l� ���l�      B  , , ���l� ���m� |��m� |��l� ���l�      B  , , ���l� ���m� `��m� `��l� ���l�      B  , , ���l� ���m� D��m� D��l� ���l�      B  , , ���p� ���q� ���q� ���p� ���p�      B  , , ���p� ���q� |��q� |��p� ���p�      B  , , ���p� ���q� `��q� `��p� ���p�      B  , , ���p� ���q� D��q� D��p� ���p�      B  , ,  �"����  �"����  ������  ������  �"����      B  , ,  �p����  �p����  �����  �����  �p����      B  , ,  ������  ������  �h����  �h����  ������      B  , ,  �����  �����  ������  ������  �����      B  , ,  �Z����  �Z����  �����  �����  �Z����      B  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      B  , ,  ������  ������  Ƞ����  Ƞ����  ������      B  , ,  �D����  �D����  ������  ������  �D����      B  , ,  �"���I  �"����  ������  �����I  �"���I      B  , ,  �p���I  �p����  �����  ����I  �p���I      B  , ,  �����I  ������  �h����  �h���I  �����I      B  , ,  ����I  �����  ������  �����I  ����I      B  , ,  �Z���I  �Z����  �����  ����I  �Z���I      B  , ,  �n��}�  �n��~s  ���~s  ���}�  �n��}�      B  , ,  �Z��|  �Z��|�  ���|�  ���|  �Z��|      B  , ,  ή��|  ή��|�  �X��|�  �X��|  ή��|      B  , ,  ���|  ���|�  Ь��|�  Ь��|  ���|      B  , ,  �V��|  �V��|�  � ��|�  � ��|  �V��|      B  , ,  ���m�  ���nt  ����nt  ����m�  ���m�      B  , ,  �\��m�  �\��nt  ���nt  ���m�  �\��m�      B  , ,  ���o  ���o�  ����o�  ����o  ���o      B  , ,  �\��o  �\��o�  ���o�  ���o  �\��o      B  , ,  º��|  º��|�  �d��|�  �d��|  º��|      B  , ,  ���|  ���|�  ĸ��|�  ĸ��|  ���|      B  , ,  ���q�  ���rp  ����rp  ����q�  ���q�      B  , ,  �\��q�  �\��rp  ���rp  ���q�  �\��q�      B  , ,  �b��|  �b��|�  ���|�  ���|  �b��|      B  , ,  ƶ��|  ƶ��|�  �`��|�  �`��|  ƶ��|      B  , ,  ���i�  ���jx  ����jx  ����i�  ���i�      B  , ,  �\��i�  �\��jx  ���jx  ���i�  �\��i�      B  , ,  ����}�  ����~s  �l��~s  �l��}�  ����}�      B  , ,  ���}�  ���~s  ����~s  ����}�  ���}�      B  , ,  �j��}�  �j��~s  ���~s  ���}�  �j��}�      B  , ,  ����}�  ����~s  �h��~s  �h��}�  ����}�      B  , ,  ���}�  ���~s  ����~s  ����}�  ���}�      B  , ,  �f��}�  �f��~s  ���~s  ���}�  �f��}�      B  , ,  º��}�  º��~s  �d��~s  �d��}�  º��}�      B  , ,  ���}�  ���~s  ĸ��~s  ĸ��}�  ���}�      B  , ,  �b��}�  �b��~s  ���~s  ���}�  �b��}�      B  , ,  ƶ��}�  ƶ��~s  �`��~s  �`��}�  ƶ��}�      B  , ,  �
��}�  �
��~s  ȴ��~s  ȴ��}�  �
��}�      B  , ,  �^��}�  �^��~s  ���~s  ���}�  �^��}�      B  , ,  ���lv  ���m   ����m   ����lv  ���lv      B  , ,  �\��lv  �\��m   ���m   ���lv  �\��lv      B  , ,  �
��|  �
��|�  ȴ��|�  ȴ��|  �
��|      B  , ,  �^��|  �^��|�  ���|�  ���|  �^��|      B  , ,  ʲ��|  ʲ��|�  �\��|�  �\��|  ʲ��|      B  , ,  ���|  ���|�  ̰��|�  ̰��|  ���|      B  , ,  ʲ��}�  ʲ��~s  �\��~s  �\��}�  ʲ��}�      B  , ,  ���}�  ���~s  ̰��~s  ̰��}�  ���}�      B  , ,  �Z��}�  �Z��~s  ���~s  ���}�  �Z��}�      B  , ,  ή��}�  ή��~s  �X��~s  �X��}�  ή��}�      B  , ,  ���}�  ���~s  Ь��~s  Ь��}�  ���}�      B  , ,  �n��|  �n��|�  ���|�  ���|  �n��|      B  , ,  ���pr  ���q  ����q  ����pr  ���pr      B  , ,  �\��pr  �\��q  ���q  ���pr  �\��pr      B  , ,  �V��}�  �V��~s  � ��~s  � ��}�  �V��}�      B  , ,  Ũ���I  Ũ����  �R����  �R���I  Ũ���I      B  , ,  �����I  ������  Ƞ����  Ƞ���I  �����I      B  , ,  �D���I  �D����  ������  �����I  �D���I      B  , ,  ����|  ����|�  �l��|�  �l��|  ����|      B  , ,  ���|  ���|�  ����|�  ����|  ���|      B  , ,  �j��|  �j��|�  ���|�  ���|  �j��|      B  , ,  ����|  ����|�  �h��|�  �h��|  ����|      B  , ,  ���|  ���|�  ����|�  ����|  ���|      B  , ,  �f��|  �f��|�  ���|�  ���|  �f��|      B  , ,  ���k"  ���k�  ����k�  ����k"  ���k"      B  , ,  �\��k"  �\��k�  ���k�  ���k"  �\��k"      B  , ,  ���Y�  ���Z~  ����Z~  ����Y�  ���Y�      B  , ,  �\��Y�  �\��Z~  ���Z~  ���Y�  �\��Y�      B  , ,  ���hz  ���i$  ����i$  ����hz  ���hz      B  , ,  �\��hz  �\��i$  ���i$  ���hz  �\��hz      B  , ,  ���`x  ���a"  ����a"  ����`x  ���`x      B  , ,  �\��`x  �\��a"  ���a"  ���`x  �\��`x      B  , ,  ���_$  ���_�  ����_�  ����_$  ���_$      B  , ,  �\��_$  �\��_�  ���_�  ���_$  �\��_$      B  , ,  ���\|  ���]&  ����]&  ����\|  ���\|      B  , ,  �\��\|  �\��]&  ���]&  ���\|  �\��\|      B  , ,  ���[(  ���[�  ����[�  ����[(  ���[(      B  , ,  �\��[(  �\��[�  ���[�  ���[(  �\��[(      B  , ,  ���a�  ���bv  ����bv  ����a�  ���a�      B  , ,  �\��a�  �\��bv  ���bv  ���a�  �\��a�      B  , ,  ���]�  ���^z  ����^z  ����]�  ���]�      B  , ,  �\��]�  �\��^z  ���^z  ���]�  �\��]�      B  , ,  ���X�  ���Y*  ����Y*  ����X�  ���X�      B  , ,  �\��X�  �\��Y*  ���Y*  ���X�  �\��X�      B  , , ���c� ���d8 `��d8 `��c� ���c�      B  , , ���c� ���d8 D��d8 D��c� ���c�      B  , , ���f6 ���f� |��f� |��f6 ���f6      B  , , ���f6 ���f� `��f� `��f6 ���f6      B  , , ���f6 ���f� D��f� D��f6 ���f6      B  , , ���d� ���e� ���e� ���d� ���d�      B  , , ���d� ���e� |��e� |��d� ���d�      B  , , ���d� ���e� `��e� `��d� ���d�      B  , , ���d� ���e� D��e� D��d� ���d�      B  , , D��`U D��`� ���`� ���`U D��`U      B  , , ���`U ���`� z��`� z��`U ���`U      B  , , ���`U ���`� ^��`� ^��`U ���`U      B  , , ���`U ���`� B��`� B��`U ���`U      B  , , 
|��`U 
|��`� &��`� &��`U 
|��`U      B  , , ���^9 ���^� z��^� z��^9 ���^9      B  , , ���^9 ���^� ^��^� ^��^9 ���^9      B  , , ���^9 ���^� B��^� B��^9 ���^9      B  , , 
|��^9 
|��^� &��^� &��^9 
|��^9      B  , , `��^9 `��^� 
��^� 
��^9 `��^9      B  , , D��^9 D��^� ���^� ���^9 D��^9      B  , , ���g� ���h4 ���h4 ���g� ���g�      B  , , ���g� ���h4 |��h4 |��g� ���g�      B  , , ���g� ���h4 `��h4 `��g� ���g�      B  , , ���g� ���h4 D��h4 D��g� ���g�      B  , , ���b: ���b� ���b� ���b: ���b:      B  , , ���b: ���b� |��b� |��b: ���b:      B  , , ���b: ���b� `��b� `��b: ���b:      B  , , ���b: ���b� D��b� D��b: ���b:      B  , , `��`U `��`� 
��`� 
��`U `��`U      B  , , ���f6 ���f� ���f� ���f6 ���f6      B  , , ���c� ���d8 ���d8 ���c� ���c�      B  , , ���c� ���d8 |��d8 |��c� ���c�      B  , , ~��h� ~��i� (��i� (��h� ~��h�      B  , , b��h� b��i� ��i� ��h� b��h�      B  , , F��h� F��i� ���i� ���h� F��h�      B  , ,  *��h�  *��i�  ���i�  ���h�  *��h�      B  , , #��h� #��i� #���i� #���h� #��h�      B  , , %���h� %���i� &���i� &���h� %���h�      B  , , (���h� (���i� )���i� )���h� (���h�      B  , , +���h� +���i� ,d��i� ,d��h� +���h�      B  , , .���h� .���i� /H��i� /H��h� .���h�      B  , , 1���h� 1���i� 2,��i� 2,��h� 1���h�      B  , , 4f��h� 4f��i� 5��i� 5��h� 4f��h�      B  , , 7J��h� 7J��i� 7���i� 7���h� 7J��h�      B  , , :.��h� :.��i� :���i� :���h� :.��h�      B  , , =��h� =��i� =���i� =���h� =��h�      B  , , ?���h� ?���i� @���i� @���h� ?���h�      B  , , B���h� B���i� C���i� C���h� B���h�      B  , , E���h� E���i� Fh��i� Fh��h� E���h�      B  , , H���h� H���i� IL��i� IL��h� H���h�      B  , , K���h� K���i� L0��i� L0��h� K���h�      B  , , Nj��h� Nj��i� O��i� O��h� Nj��h�      B  , , QN��h� QN��i� Q���i� Q���h� QN��h�      B  , , T2��h� T2��i� T���i� T���h� T2��h�      B  , , W��h� W��i� W���i� W���h� W��h�      B  , , Y���h� Y���i� Z���i� Z���h� Y���h�      B  , , \���h� \���i� ]���i� ]���h� \���h�      B  , , _���h� _���i� `l��i� `l��h� _���h�      B  , , b���h� b���i� cP��i� cP��h� b���h�      B  , , e���h� e���i� f4��i� f4��h� e���h�      B  , , hn��h� hn��i� i��i� i��h� hn��h�      B  , , kR��h� kR��i� k���i� k���h� kR��h�      B  , , n6��h� n6��i� n���i� n���h� n6��h�      B  , , q��h� q��i� q���i� q���h� q��h�      B  , , E���j2 E���j� Fh��j� Fh��j2 E���j2      B  , , H���j2 H���j� IL��j� IL��j2 H���j2      B  , , K���j2 K���j� L0��j� L0��j2 K���j2      B  , , Nj��j2 Nj��j� O��j� O��j2 Nj��j2      B  , , QN��j2 QN��j� Q���j� Q���j2 QN��j2      B  , , T2��j2 T2��j� T���j� T���j2 T2��j2      B  , , W��j2 W��j� W���j� W���j2 W��j2      B  , , Y���j2 Y���j� Z���j� Z���j2 Y���j2      B  , , E���p� E���q� Fh��q� Fh��p� E���p�      B  , , H���p� H���q� IL��q� IL��p� H���p�      B  , , K���p� K���q� L0��q� L0��p� K���p�      B  , , Nj��p� Nj��q� O��q� O��p� Nj��p�      B  , , QN��p� QN��q� Q���q� Q���p� QN��p�      B  , , T2��p� T2��q� T���q� T���p� T2��p�      B  , , W��p� W��q� W���q� W���p� W��p�      B  , , Y���p� Y���q� Z���q� Z���p� Y���p�      B  , , E���k� E���l0 Fh��l0 Fh��k� E���k�      B  , , H���k� H���l0 IL��l0 IL��k� H���k�      B  , , K���k� K���l0 L0��l0 L0��k� K���k�      B  , , Nj��k� Nj��l0 O��l0 O��k� Nj��k�      B  , , QN��k� QN��l0 Q���l0 Q���k� QN��k�      B  , , T2��k� T2��l0 T���l0 T���k� T2��k�      B  , , W��k� W��l0 W���l0 W���k� W��k�      B  , , Y���k� Y���l0 Z���l0 Z���k� Y���k�      B  , , E���o� E���p, Fh��p, Fh��o� E���o�      B  , , H���o� H���p, IL��p, IL��o� H���o�      B  , , K���o� K���p, L0��p, L0��o� K���o�      B  , , Nj��o� Nj��p, O��p, O��o� Nj��o�      B  , , QN��o� QN��p, Q���p, Q���o� QN��o�      B  , , T2��o� T2��p, T���p, T���o� T2��o�      B  , , W��o� W��p, W���p, W���o� W��o�      B  , , Y���o� Y���p, Z���p, Z���o� Y���o�      B  , , E���n. E���n� Fh��n� Fh��n. E���n.      B  , , H���n. H���n� IL��n� IL��n. H���n.      B  , , K���n. K���n� L0��n� L0��n. K���n.      B  , , Nj��n. Nj��n� O��n� O��n. Nj��n.      B  , , QN��n. QN��n� Q���n� Q���n. QN��n.      B  , , T2��n. T2��n� T���n� T���n. T2��n.      B  , , W��n. W��n� W���n� W���n. W��n.      B  , , Y���n. Y���n� Z���n� Z���n. Y���n.      B  , , E���r* E���r� Fh��r� Fh��r* E���r*      B  , , H���r* H���r� IL��r� IL��r* H���r*      B  , , K���r* K���r� L0��r� L0��r* K���r*      B  , , Nj��r* Nj��r� O��r� O��r* Nj��r*      B  , , QN��r* QN��r� Q���r� Q���r* QN��r*      B  , , T2��r* T2��r� T���r� T���r* T2��r*      B  , , W��r* W��r� W���r� W���r* W��r*      B  , , Y���r* Y���r� Z���r� Z���r* Y���r*      B  , , E���l� E���m� Fh��m� Fh��l� E���l�      B  , , H���l� H���m� IL��m� IL��l� H���l�      B  , , K���l� K���m� L0��m� L0��l� K���l�      B  , , Nj��l� Nj��m� O��m� O��l� Nj��l�      B  , , QN��l� QN��m� Q���m� Q���l� QN��l�      B  , , T2��l� T2��m� T���m� T���l� T2��l�      B  , , W��l� W��m� W���m� W���l� W��l�      B  , , Y���l� Y���m� Z���m� Z���l� Y���l�      B  , , \���j2 \���j� ]���j� ]���j2 \���j2      B  , , _���j2 _���j� `l��j� `l��j2 _���j2      B  , , b���j2 b���j� cP��j� cP��j2 b���j2      B  , , e���j2 e���j� f4��j� f4��j2 e���j2      B  , , hn��j2 hn��j� i��j� i��j2 hn��j2      B  , , kR��j2 kR��j� k���j� k���j2 kR��j2      B  , , n6��j2 n6��j� n���j� n���j2 n6��j2      B  , , q��j2 q��j� q���j� q���j2 q��j2      B  , , \���o� \���p, ]���p, ]���o� \���o�      B  , , _���o� _���p, `l��p, `l��o� _���o�      B  , , b���o� b���p, cP��p, cP��o� b���o�      B  , , e���o� e���p, f4��p, f4��o� e���o�      B  , , hn��o� hn��p, i��p, i��o� hn��o�      B  , , kR��o� kR��p, k���p, k���o� kR��o�      B  , , n6��o� n6��p, n���p, n���o� n6��o�      B  , , q��o� q��p, q���p, q���o� q��o�      B  , , \���p� \���q� ]���q� ]���p� \���p�      B  , , _���p� _���q� `l��q� `l��p� _���p�      B  , , b���p� b���q� cP��q� cP��p� b���p�      B  , , e���p� e���q� f4��q� f4��p� e���p�      B  , , hn��p� hn��q� i��q� i��p� hn��p�      B  , , kR��p� kR��q� k���q� k���p� kR��p�      B  , , n6��p� n6��q� n���q� n���p� n6��p�      B  , , q��p� q��q� q���q� q���p� q��p�      B  , , \���n. \���n� ]���n� ]���n. \���n.      B  , , _���n. _���n� `l��n� `l��n. _���n.      B  , , b���n. b���n� cP��n� cP��n. b���n.      B  , , e���n. e���n� f4��n� f4��n. e���n.      B  , , hn��n. hn��n� i��n� i��n. hn��n.      B  , , kR��n. kR��n� k���n� k���n. kR��n.      B  , , n6��n. n6��n� n���n� n���n. n6��n.      B  , , q��n. q��n� q���n� q���n. q��n.      B  , , \���r* \���r� ]���r� ]���r* \���r*      B  , , _���r* _���r� `l��r� `l��r* _���r*      B  , , b���r* b���r� cP��r� cP��r* b���r*      B  , , e���r* e���r� f4��r� f4��r* e���r*      B  , , hn��r* hn��r� i��r� i��r* hn��r*      B  , , kR��r* kR��r� k���r� k���r* kR��r*      B  , , n6��r* n6��r� n���r� n���r* n6��r*      B  , , q��r* q��r� q���r� q���r* q��r*      B  , , \���k� \���l0 ]���l0 ]���k� \���k�      B  , , _���k� _���l0 `l��l0 `l��k� _���k�      B  , , b���k� b���l0 cP��l0 cP��k� b���k�      B  , , e���k� e���l0 f4��l0 f4��k� e���k�      B  , , hn��k� hn��l0 i��l0 i��k� hn��k�      B  , , kR��k� kR��l0 k���l0 k���k� kR��k�      B  , , n6��k� n6��l0 n���l0 n���k� n6��k�      B  , , q��k� q��l0 q���l0 q���k� q��k�      B  , , \���l� \���m� ]���m� ]���l� \���l�      B  , , _���l� _���m� `l��m� `l��l� _���l�      B  , , b���l� b���m� cP��m� cP��l� b���l�      B  , , e���l� e���m� f4��m� f4��l� e���l�      B  , , hn��l� hn��m� i��m� i��l� hn��l�      B  , , kR��l� kR��m� k���m� k���l� kR��l�      B  , , n6��l� n6��m� n���m� n���l� n6��l�      B  , , q��l� q��m� q���m� q���l� q��l�      B  , , #��j2 #��j� #���j� #���j2 #��j2      B  , , %���j2 %���j� &���j� &���j2 %���j2      B  , , (���j2 (���j� )���j� )���j2 (���j2      B  , , +���j2 +���j� ,d��j� ,d��j2 +���j2      B  , , ~��r* ~��r� (��r� (��r* ~��r*      B  , , b��r* b��r� ��r� ��r* b��r*      B  , , F��r* F��r� ���r� ���r* F��r*      B  , ,  *��r*  *��r�  ���r�  ���r*  *��r*      B  , , #��r* #��r� #���r� #���r* #��r*      B  , , %���r* %���r� &���r� &���r* %���r*      B  , , (���r* (���r� )���r� )���r* (���r*      B  , , +���r* +���r� ,d��r� ,d��r* +���r*      B  , , ~��n. ~��n� (��n� (��n. ~��n.      B  , , b��n. b��n� ��n� ��n. b��n.      B  , , F��n. F��n� ���n� ���n. F��n.      B  , ,  *��n.  *��n�  ���n�  ���n.  *��n.      B  , , #��n. #��n� #���n� #���n. #��n.      B  , , %���n. %���n� &���n� &���n. %���n.      B  , , (���n. (���n� )���n� )���n. (���n.      B  , , +���n. +���n� ,d��n� ,d��n. +���n.      B  , , ~��k� ~��l0 (��l0 (��k� ~��k�      B  , , b��k� b��l0 ��l0 ��k� b��k�      B  , , F��k� F��l0 ���l0 ���k� F��k�      B  , ,  *��k�  *��l0  ���l0  ���k�  *��k�      B  , , #��k� #��l0 #���l0 #���k� #��k�      B  , , %���k� %���l0 &���l0 &���k� %���k�      B  , , (���k� (���l0 )���l0 )���k� (���k�      B  , , +���k� +���l0 ,d��l0 ,d��k� +���k�      B  , , ~��o� ~��p, (��p, (��o� ~��o�      B  , , b��o� b��p, ��p, ��o� b��o�      B  , , F��o� F��p, ���p, ���o� F��o�      B  , ,  *��o�  *��p,  ���p,  ���o�  *��o�      B  , , ~��p� ~��q� (��q� (��p� ~��p�      B  , , b��p� b��q� ��q� ��p� b��p�      B  , , F��p� F��q� ���q� ���p� F��p�      B  , ,  *��p�  *��q�  ���q�  ���p�  *��p�      B  , , #��p� #��q� #���q� #���p� #��p�      B  , , %���p� %���q� &���q� &���p� %���p�      B  , , (���p� (���q� )���q� )���p� (���p�      B  , , +���p� +���q� ,d��q� ,d��p� +���p�      B  , , ~��l� ~��m� (��m� (��l� ~��l�      B  , , b��l� b��m� ��m� ��l� b��l�      B  , , F��l� F��m� ���m� ���l� F��l�      B  , ,  *��l�  *��m�  ���m�  ���l�  *��l�      B  , , #��l� #��m� #���m� #���l� #��l�      B  , , %���l� %���m� &���m� &���l� %���l�      B  , , (���l� (���m� )���m� )���l� (���l�      B  , , +���l� +���m� ,d��m� ,d��l� +���l�      B  , , #��o� #��p, #���p, #���o� #��o�      B  , , %���o� %���p, &���p, &���o� %���o�      B  , , (���o� (���p, )���p, )���o� (���o�      B  , , +���o� +���p, ,d��p, ,d��o� +���o�      B  , , ~��j2 ~��j� (��j� (��j2 ~��j2      B  , , b��j2 b��j� ��j� ��j2 b��j2      B  , , F��j2 F��j� ���j� ���j2 F��j2      B  , ,  *��j2  *��j�  ���j�  ���j2  *��j2      B  , , :.��r* :.��r� :���r� :���r* :.��r*      B  , , =��r* =��r� =���r� =���r* =��r*      B  , , ?���r* ?���r� @���r� @���r* ?���r*      B  , , B���r* B���r� C���r� C���r* B���r*      B  , , .���k� .���l0 /H��l0 /H��k� .���k�      B  , , 1���k� 1���l0 2,��l0 2,��k� 1���k�      B  , , 4f��k� 4f��l0 5��l0 5��k� 4f��k�      B  , , 7J��k� 7J��l0 7���l0 7���k� 7J��k�      B  , , :.��j2 :.��j� :���j� :���j2 :.��j2      B  , , =��j2 =��j� =���j� =���j2 =��j2      B  , , ?���j2 ?���j� @���j� @���j2 ?���j2      B  , , B���j2 B���j� C���j� C���j2 B���j2      B  , , .���n. .���n� /H��n� /H��n. .���n.      B  , , 1���n. 1���n� 2,��n� 2,��n. 1���n.      B  , , 4f��n. 4f��n� 5��n� 5��n. 4f��n.      B  , , 7J��n. 7J��n� 7���n� 7���n. 7J��n.      B  , , :.��n. :.��n� :���n� :���n. :.��n.      B  , , =��n. =��n� =���n� =���n. =��n.      B  , , ?���n. ?���n� @���n� @���n. ?���n.      B  , , B���n. B���n� C���n� C���n. B���n.      B  , , .���p� .���q� /H��q� /H��p� .���p�      B  , , 1���p� 1���q� 2,��q� 2,��p� 1���p�      B  , , 4f��p� 4f��q� 5��q� 5��p� 4f��p�      B  , , 7J��p� 7J��q� 7���q� 7���p� 7J��p�      B  , , :.��k� :.��l0 :���l0 :���k� :.��k�      B  , , =��k� =��l0 =���l0 =���k� =��k�      B  , , ?���k� ?���l0 @���l0 @���k� ?���k�      B  , , B���k� B���l0 C���l0 C���k� B���k�      B  , , :.��p� :.��q� :���q� :���p� :.��p�      B  , , =��p� =��q� =���q� =���p� =��p�      B  , , ?���p� ?���q� @���q� @���p� ?���p�      B  , , B���p� B���q� C���q� C���p� B���p�      B  , , .���l� .���m� /H��m� /H��l� .���l�      B  , , 1���l� 1���m� 2,��m� 2,��l� 1���l�      B  , , 4f��l� 4f��m� 5��m� 5��l� 4f��l�      B  , , 7J��l� 7J��m� 7���m� 7���l� 7J��l�      B  , , :.��l� :.��m� :���m� :���l� :.��l�      B  , , =��l� =��m� =���m� =���l� =��l�      B  , , ?���l� ?���m� @���m� @���l� ?���l�      B  , , B���l� B���m� C���m� C���l� B���l�      B  , , .���r* .���r� /H��r� /H��r* .���r*      B  , , 1���r* 1���r� 2,��r� 2,��r* 1���r*      B  , , 4f��r* 4f��r� 5��r� 5��r* 4f��r*      B  , , 7J��r* 7J��r� 7���r� 7���r* 7J��r*      B  , , .���o� .���p, /H��p, /H��o� .���o�      B  , , 1���o� 1���p, 2,��p, 2,��o� 1���o�      B  , , 4f��o� 4f��p, 5��p, 5��o� 4f��o�      B  , , 7J��o� 7J��p, 7���p, 7���o� 7J��o�      B  , , :.��o� :.��p, :���p, :���o� :.��o�      B  , , =��o� =��p, =���p, =���o� =��o�      B  , , ?���o� ?���p, @���p, @���o� ?���o�      B  , , B���o� B���p, C���p, C���o� B���o�      B  , , .���j2 .���j� /H��j� /H��j2 .���j2      B  , , 1���j2 1���j� 2,��j� 2,��j2 1���j2      B  , , 4f��j2 4f��j� 5��j� 5��j2 4f��j2      B  , , 7J��j2 7J��j� 7���j� 7���j2 7J��j2      B  , , =��f6 =��f� =���f� =���f6 =��f6      B  , , ?���f6 ?���f� @���f� @���f6 ?���f6      B  , , B���f6 B���f� C���f� C���f6 B���f6      B  , ,  *��g�  *��h4  ���h4  ���g�  *��g�      B  , , 0��`U 0��`� 0���`� 0���`U 0��`U      B  , , 2���`U 2���`� 3���`� 3���`U 2���`U      B  , , 5���`U 5���`� 6���`� 6���`U 5���`U      B  , , 8���`U 8���`� 9f��`� 9f��`U 8���`U      B  , , ;���`U ;���`� <J��`� <J��`U ;���`U      B  , , >���`U >���`� ?.��`� ?.��`U >���`U      B  , , Ah��`U Ah��`� B��`� B��`U Ah��`U      B  , , #��g� #��h4 #���h4 #���g� #��g�      B  , , %���g� %���h4 &���h4 &���g� %���g�      B  , , (���g� (���h4 )���h4 )���g� (���g�      B  , , ~��d� ~��e� (��e� (��d� ~��d�      B  , , b��d� b��e� ��e� ��d� b��d�      B  , , F��d� F��e� ���e� ���d� F��d�      B  , ,  *��d�  *��e�  ���e�  ���d�  *��d�      B  , , #��d� #��e� #���e� #���d� #��d�      B  , , %���d� %���e� &���e� &���d� %���d�      B  , , (���d� (���e� )���e� )���d� (���d�      B  , , +���d� +���e� ,d��e� ,d��d� +���d�      B  , , .���d� .���e� /H��e� /H��d� .���d�      B  , , 1���d� 1���e� 2,��e� 2,��d� 1���d�      B  , , 4f��d� 4f��e� 5��e� 5��d� 4f��d�      B  , , 7J��d� 7J��e� 7���e� 7���d� 7J��d�      B  , , :.��d� :.��e� :���e� :���d� :.��d�      B  , , =��d� =��e� =���e� =���d� =��d�      B  , , ?���d� ?���e� @���e� @���d� ?���d�      B  , , B���d� B���e� C���e� C���d� B���d�      B  , , +���g� +���h4 ,d��h4 ,d��g� +���g�      B  , , 0��^9 0��^� 0���^� 0���^9 0��^9      B  , , 2���^9 2���^� 3���^� 3���^9 2���^9      B  , , 5���^9 5���^� 6���^� 6���^9 5���^9      B  , , 8���^9 8���^� 9f��^� 9f��^9 8���^9      B  , , ;���^9 ;���^� <J��^� <J��^9 ;���^9      B  , , >���^9 >���^� ?.��^� ?.��^9 >���^9      B  , , Ah��^9 Ah��^� B��^� B��^9 Ah��^9      B  , , .���g� .���h4 /H��h4 /H��g� .���g�      B  , , 1���g� 1���h4 2,��h4 2,��g� 1���g�      B  , , 4f��g� 4f��h4 5��h4 5��g� 4f��g�      B  , , 7J��g� 7J��h4 7���h4 7���g� 7J��g�      B  , , ~��c� ~��d8 (��d8 (��c� ~��c�      B  , , b��c� b��d8 ��d8 ��c� b��c�      B  , , F��c� F��d8 ���d8 ���c� F��c�      B  , ,  *��c�  *��d8  ���d8  ���c�  *��c�      B  , , #��c� #��d8 #���d8 #���c� #��c�      B  , , %���c� %���d8 &���d8 &���c� %���c�      B  , , (���c� (���d8 )���d8 )���c� (���c�      B  , , +���c� +���d8 ,d��d8 ,d��c� +���c�      B  , , .���c� .���d8 /H��d8 /H��c� .���c�      B  , , 1���c� 1���d8 2,��d8 2,��c� 1���c�      B  , , 4f��c� 4f��d8 5��d8 5��c� 4f��c�      B  , , 7J��c� 7J��d8 7���d8 7���c� 7J��c�      B  , , :.��c� :.��d8 :���d8 :���c� :.��c�      B  , , =��c� =��d8 =���d8 =���c� =��c�      B  , , ?���c� ?���d8 @���d8 @���c� ?���c�      B  , , B���c� B���d8 C���d8 C���c� B���c�      B  , , ~��b: ~��b� (��b� (��b: ~��b:      B  , , b��b: b��b� ��b� ��b: b��b:      B  , , F��b: F��b� ���b� ���b: F��b:      B  , ,  *��b:  *��b�  ���b�  ���b:  *��b:      B  , , #��b: #��b� #���b� #���b: #��b:      B  , , %���b: %���b� &���b� &���b: %���b:      B  , , (���b: (���b� )���b� )���b: (���b:      B  , , +���b: +���b� ,d��b� ,d��b: +���b:      B  , , .���b: .���b� /H��b� /H��b: .���b:      B  , , 1���b: 1���b� 2,��b� 2,��b: 1���b:      B  , , 4f��b: 4f��b� 5��b� 5��b: 4f��b:      B  , , 7J��b: 7J��b� 7���b� 7���b: 7J��b:      B  , , :.��b: :.��b� :���b� :���b: :.��b:      B  , , =��b: =��b� =���b� =���b: =��b:      B  , , ?���b: ?���b� @���b� @���b: ?���b:      B  , , B���b: B���b� C���b� C���b: B���b:      B  , , :.��g� :.��h4 :���h4 :���g� :.��g�      B  , , =��g� =��h4 =���h4 =���g� =��g�      B  , , ?���g� ?���h4 @���h4 @���g� ?���g�      B  , , B���g� B���h4 C���h4 C���g� B���g�      B  , , ~��g� ~��h4 (��h4 (��g� ~��g�      B  , , b��g� b��h4 ��h4 ��g� b��g�      B  , , F��g� F��h4 ���h4 ���g� F��g�      B  , , ~��f6 ~��f� (��f� (��f6 ~��f6      B  , , b��f6 b��f� ��f� ��f6 b��f6      B  , , F��f6 F��f� ���f� ���f6 F��f6      B  , ,  *��f6  *��f�  ���f�  ���f6  *��f6      B  , , #��f6 #��f� #���f� #���f6 #��f6      B  , , %���f6 %���f� &���f� &���f6 %���f6      B  , , (���f6 (���f� )���f� )���f6 (���f6      B  , , +���f6 +���f� ,d��f� ,d��f6 +���f6      B  , , .���f6 .���f� /H��f� /H��f6 .���f6      B  , , 1���f6 1���f� 2,��f� 2,��f6 1���f6      B  , , 4f��f6 4f��f� 5��f� 5��f6 4f��f6      B  , , 7J��f6 7J��f� 7���f� 7���f6 7J��f6      B  , , :.��f6 :.��f� :���f� :���f6 :.��f6      B  , , [l��`U [l��`� \��`� \��`U [l��`U      B  , , ^P��`U ^P��`� ^���`� ^���`U ^P��`U      B  , , a4��`U a4��`� a���`� a���`U a4��`U      B  , , d��`U d��`� d���`� d���`U d��`U      B  , , f���`U f���`� g���`� g���`U f���`U      B  , , e���g� e���h4 f4��h4 f4��g� e���g�      B  , , \���c� \���d8 ]���d8 ]���c� \���c�      B  , , _���c� _���d8 `l��d8 `l��c� _���c�      B  , , b���c� b���d8 cP��d8 cP��c� b���c�      B  , , e���c� e���d8 f4��d8 f4��c� e���c�      B  , , hn��c� hn��d8 i��d8 i��c� hn��c�      B  , , kR��c� kR��d8 k���d8 k���c� kR��c�      B  , , n6��c� n6��d8 n���d8 n���c� n6��c�      B  , , q��c� q��d8 q���d8 q���c� q��c�      B  , , hn��g� hn��h4 i��h4 i��g� hn��g�      B  , , kR��g� kR��h4 k���h4 k���g� kR��g�      B  , , n6��g� n6��h4 n���h4 n���g� n6��g�      B  , , q��g� q��h4 q���h4 q���g� q��g�      B  , , [l��^9 [l��^� \��^� \��^9 [l��^9      B  , , ^P��^9 ^P��^� ^���^� ^���^9 ^P��^9      B  , , a4��^9 a4��^� a���^� a���^9 a4��^9      B  , , d��^9 d��^� d���^� d���^9 d��^9      B  , , f���^9 f���^� g���^� g���^9 f���^9      B  , , \���b: \���b� ]���b� ]���b: \���b:      B  , , _���b: _���b� `l��b� `l��b: _���b:      B  , , b���b: b���b� cP��b� cP��b: b���b:      B  , , e���b: e���b� f4��b� f4��b: e���b:      B  , , hn��b: hn��b� i��b� i��b: hn��b:      B  , , kR��b: kR��b� k���b� k���b: kR��b:      B  , , n6��b: n6��b� n���b� n���b: n6��b:      B  , , q��b: q��b� q���b� q���b: q��b:      B  , , \���d� \���e� ]���e� ]���d� \���d�      B  , , _���d� _���e� `l��e� `l��d� _���d�      B  , , b���d� b���e� cP��e� cP��d� b���d�      B  , , e���d� e���e� f4��e� f4��d� e���d�      B  , , hn��d� hn��e� i��e� i��d� hn��d�      B  , , kR��d� kR��e� k���e� k���d� kR��d�      B  , , n6��d� n6��e� n���e� n���d� n6��d�      B  , , q��d� q��e� q���e� q���d� q��d�      B  , , \���f6 \���f� ]���f� ]���f6 \���f6      B  , , _���f6 _���f� `l��f� `l��f6 _���f6      B  , , b���f6 b���f� cP��f� cP��f6 b���f6      B  , , e���f6 e���f� f4��f� f4��f6 e���f6      B  , , hn��f6 hn��f� i��f� i��f6 hn��f6      B  , , kR��f6 kR��f� k���f� k���f6 kR��f6      B  , , n6��f6 n6��f� n���f� n���f6 n6��f6      B  , , q��f6 q��f� q���f� q���f6 q��f6      B  , , \���g� \���h4 ]���h4 ]���g� \���g�      B  , , _���g� _���h4 `l��h4 `l��g� _���g�      B  , , b���g� b���h4 cP��h4 cP��g� b���g�      B  , , Nj��f6 Nj��f� O��f� O��f6 Nj��f6      B  , , E���d� E���e� Fh��e� Fh��d� E���d�      B  , , H���d� H���e� IL��e� IL��d� H���d�      B  , , K���d� K���e� L0��e� L0��d� K���d�      B  , , Nj��d� Nj��e� O��e� O��d� Nj��d�      B  , , QN��d� QN��e� Q���e� Q���d� QN��d�      B  , , E���b: E���b� Fh��b� Fh��b: E���b:      B  , , H���b: H���b� IL��b� IL��b: H���b:      B  , , K���b: K���b� L0��b� L0��b: K���b:      B  , , Nj��b: Nj��b� O��b� O��b: Nj��b:      B  , , QN��b: QN��b� Q���b� Q���b: QN��b:      B  , , T2��b: T2��b� T���b� T���b: T2��b:      B  , , W��b: W��b� W���b� W���b: W��b:      B  , , Y���b: Y���b� Z���b� Z���b: Y���b:      B  , , L���`U L���`� M���`� M���`U L���`U      B  , , E���c� E���d8 Fh��d8 Fh��c� E���c�      B  , , H���c� H���d8 IL��d8 IL��c� H���c�      B  , , K���c� K���d8 L0��d8 L0��c� K���c�      B  , , Nj��c� Nj��d8 O��d8 O��c� Nj��c�      B  , , QN��c� QN��d8 Q���d8 Q���c� QN��c�      B  , , T2��c� T2��d8 T���d8 T���c� T2��c�      B  , , W��c� W��d8 W���d8 W���c� W��c�      B  , , T2��d� T2��e� T���e� T���d� T2��d�      B  , , W��d� W��e� W���e� W���d� W��d�      B  , , Y���d� Y���e� Z���e� Z���d� Y���d�      B  , , E���g� E���h4 Fh��h4 Fh��g� E���g�      B  , , H���g� H���h4 IL��h4 IL��g� H���g�      B  , , K���g� K���h4 L0��h4 L0��g� K���g�      B  , , E���f6 E���f� Fh��f� Fh��f6 E���f6      B  , , H���f6 H���f� IL��f� IL��f6 H���f6      B  , , K���f6 K���f� L0��f� L0��f6 K���f6      B  , , DL��^9 DL��^� D���^� D���^9 DL��^9      B  , , G0��^9 G0��^� G���^� G���^9 G0��^9      B  , , QN��f6 QN��f� Q���f� Q���f6 QN��f6      B  , , T2��f6 T2��f� T���f� T���f6 T2��f6      B  , , W��f6 W��f� W���f� W���f6 W��f6      B  , , Y���f6 Y���f� Z���f� Z���f6 Y���f6      B  , , J��^9 J��^� J���^� J���^9 J��^9      B  , , L���^9 L���^� M���^� M���^9 L���^9      B  , , O���^9 O���^� P���^� P���^9 O���^9      B  , , R���^9 R���^� Sj��^� Sj��^9 R���^9      B  , , U���^9 U���^� VN��^� VN��^9 U���^9      B  , , X���^9 X���^� Y2��^� Y2��^9 X���^9      B  , , Y���c� Y���d8 Z���d8 Z���c� Y���c�      B  , , O���`U O���`� P���`� P���`U O���`U      B  , , Nj��g� Nj��h4 O��h4 O��g� Nj��g�      B  , , QN��g� QN��h4 Q���h4 Q���g� QN��g�      B  , , T2��g� T2��h4 T���h4 T���g� T2��g�      B  , , W��g� W��h4 W���h4 W���g� W��g�      B  , , Y���g� Y���h4 Z���h4 Z���g� Y���g�      B  , , R���`U R���`� Sj��`� Sj��`U R���`U      B  , , U���`U U���`� VN��`� VN��`U U���`U      B  , , X���`U X���`� Y2��`� Y2��`U X���`U      B  , , DL��`U DL��`� D���`� D���`U DL��`U      B  , , G0��`U G0��`� G���`� G���`U G0��`U      B  , , J��`U J��`� J���`� J���`U J��`U      B  , , �"��h� �"��i� ����i� ����h� �"��h�      B  , , ���h� ���i� ����i� ����h� ���h�      B  , , ����h� ����i� ����i� ����h� ����h�      B  , , ����h� ����i� �x��i� �x��h� ����h�      B  , , ����h� ����i� �\��i� �\��h� ����h�      B  , , ����h� ����i� �@��i� �@��h� ����h�      B  , , �z��h� �z��i� �$��i� �$��h� �z��h�      B  , , �^��h� �^��i� ���i� ���h� �^��h�      B  , , �B��h� �B��i� ����i� ����h� �B��h�      B  , , �&��h� �&��i� ����i� ����h� �&��h�      B  , , �
��h� �
��i� ´��i� ´��h� �
��h�      B  , , s���h� s���i� t���i� t���h� s���h�      B  , , v���h� v���i� w���i� w���h� v���h�      B  , , y���h� y���i� zp��i� zp��h� y���h�      B  , , |���h� |���i� }T��i� }T��h� |���h�      B  , , ���h� ���i� �8��i� �8��h� ���h�      B  , , �r��h� �r��i� ���i� ���h� �r��h�      B  , , �V��h� �V��i� � ��i� � ��h� �V��h�      B  , , �:��h� �:��i� ����i� ����h� �:��h�      B  , , ���h� ���i� ����i� ����h� ���h�      B  , , ���h� ���i� ����i� ����h� ���h�      B  , , ����h� ����i� ����i� ����h� ����h�      B  , , ����h� ����i� �t��i� �t��h� ����h�      B  , , ����h� ����i� �X��i� �X��h� ����h�      B  , , ����h� ����i� �<��i� �<��h� ����h�      B  , , �v��h� �v��i� � ��i� � ��h� �v��h�      B  , , �Z��h� �Z��i� ���i� ���h� �Z��h�      B  , , �>��h� �>��i� ����i� ����h� �>��h�      B  , , �
��o� �
��p, ´��p, ´��o� �
��o�      B  , , �>��r* �>��r� ����r� ����r* �>��r*      B  , , �"��r* �"��r� ����r� ����r* �"��r*      B  , , ���r* ���r� ����r� ����r* ���r*      B  , , ����r* ����r� ����r� ����r* ����r*      B  , , ����r* ����r� �x��r� �x��r* ����r*      B  , , ����r* ����r� �\��r� �\��r* ����r*      B  , , ����r* ����r� �@��r� �@��r* ����r*      B  , , �z��r* �z��r� �$��r� �$��r* �z��r*      B  , , �^��r* �^��r� ���r� ���r* �^��r*      B  , , �B��r* �B��r� ����r� ����r* �B��r*      B  , , �&��r* �&��r� ����r� ����r* �&��r*      B  , , �
��r* �
��r� ´��r� ´��r* �
��r*      B  , , �>��j2 �>��j� ����j� ����j2 �>��j2      B  , , �"��j2 �"��j� ����j� ����j2 �"��j2      B  , , ���j2 ���j� ����j� ����j2 ���j2      B  , , ����j2 ����j� ����j� ����j2 ����j2      B  , , ����j2 ����j� �x��j� �x��j2 ����j2      B  , , ����j2 ����j� �\��j� �\��j2 ����j2      B  , , ����j2 ����j� �@��j� �@��j2 ����j2      B  , , �z��j2 �z��j� �$��j� �$��j2 �z��j2      B  , , �^��j2 �^��j� ���j� ���j2 �^��j2      B  , , �B��j2 �B��j� ����j� ����j2 �B��j2      B  , , �&��j2 �&��j� ����j� ����j2 �&��j2      B  , , �
��j2 �
��j� ´��j� ´��j2 �
��j2      B  , , ����k� ����l0 �@��l0 �@��k� ����k�      B  , , �z��k� �z��l0 �$��l0 �$��k� �z��k�      B  , , �^��k� �^��l0 ���l0 ���k� �^��k�      B  , , �B��k� �B��l0 ����l0 ����k� �B��k�      B  , , �&��k� �&��l0 ����l0 ����k� �&��k�      B  , , �
��k� �
��l0 ´��l0 ´��k� �
��k�      B  , , �>��p� �>��q� ����q� ����p� �>��p�      B  , , �"��p� �"��q� ����q� ����p� �"��p�      B  , , ���p� ���q� ����q� ����p� ���p�      B  , , �>��n. �>��n� ����n� ����n. �>��n.      B  , , �"��n. �"��n� ����n� ����n. �"��n.      B  , , ���n. ���n� ����n� ����n. ���n.      B  , , ����n. ����n� ����n� ����n. ����n.      B  , , ����n. ����n� �x��n� �x��n. ����n.      B  , , ����n. ����n� �\��n� �\��n. ����n.      B  , , ����n. ����n� �@��n� �@��n. ����n.      B  , , �z��n. �z��n� �$��n� �$��n. �z��n.      B  , , �^��n. �^��n� ���n� ���n. �^��n.      B  , , �B��n. �B��n� ����n� ����n. �B��n.      B  , , �&��n. �&��n� ����n� ����n. �&��n.      B  , , �
��n. �
��n� ´��n� ´��n. �
��n.      B  , , ����p� ����q� ����q� ����p� ����p�      B  , , ����p� ����q� �x��q� �x��p� ����p�      B  , , ����p� ����q� �\��q� �\��p� ����p�      B  , , ����p� ����q� �@��q� �@��p� ����p�      B  , , �z��p� �z��q� �$��q� �$��p� �z��p�      B  , , �^��p� �^��q� ���q� ���p� �^��p�      B  , , �B��p� �B��q� ����q� ����p� �B��p�      B  , , �&��p� �&��q� ����q� ����p� �&��p�      B  , , �
��p� �
��q� ´��q� ´��p� �
��p�      B  , , �&��l� �&��m� ����m� ����l� �&��l�      B  , , �
��l� �
��m� ´��m� ´��l� �
��l�      B  , , ����l� ����m� �@��m� �@��l� ����l�      B  , , �z��l� �z��m� �$��m� �$��l� �z��l�      B  , , �^��l� �^��m� ���m� ���l� �^��l�      B  , , �B��l� �B��m� ����m� ����l� �B��l�      B  , , �>��k� �>��l0 ����l0 ����k� �>��k�      B  , , �"��k� �"��l0 ����l0 ����k� �"��k�      B  , , ���k� ���l0 ����l0 ����k� ���k�      B  , , ����k� ����l0 ����l0 ����k� ����k�      B  , , ����k� ����l0 �x��l0 �x��k� ����k�      B  , , ����k� ����l0 �\��l0 �\��k� ����k�      B  , , �>��o� �>��p, ����p, ����o� �>��o�      B  , , �"��o� �"��p, ����p, ����o� �"��o�      B  , , ���o� ���p, ����p, ����o� ���o�      B  , , ����o� ����p, ����p, ����o� ����o�      B  , , ����o� ����p, �x��p, �x��o� ����o�      B  , , ����o� ����p, �\��p, �\��o� ����o�      B  , , ����o� ����p, �@��p, �@��o� ����o�      B  , , �z��o� �z��p, �$��p, �$��o� �z��o�      B  , , �^��o� �^��p, ���p, ���o� �^��o�      B  , , �B��o� �B��p, ����p, ����o� �B��o�      B  , , �&��o� �&��p, ����p, ����o� �&��o�      B  , , �>��l� �>��m� ����m� ����l� �>��l�      B  , , �"��l� �"��m� ����m� ����l� �"��l�      B  , , ���l� ���m� ����m� ����l� ���l�      B  , , ����l� ����m� ����m� ����l� ����l�      B  , , ����l� ����m� �x��m� �x��l� ����l�      B  , , ����l� ����m� �\��m� �\��l� ����l�      B  , , |���r* |���r� }T��r� }T��r* |���r*      B  , , ���r* ���r� �8��r� �8��r* ���r*      B  , , �r��r* �r��r� ���r� ���r* �r��r*      B  , , �V��r* �V��r� � ��r� � ��r* �V��r*      B  , , �:��r* �:��r� ����r� ����r* �:��r*      B  , , �V��p� �V��q� � ��q� � ��p� �V��p�      B  , , �:��p� �:��q� ����q� ����p� �:��p�      B  , , ���o� ���p, �8��p, �8��o� ���o�      B  , , �r��o� �r��p, ���p, ���o� �r��o�      B  , , s���k� s���l0 t���l0 t���k� s���k�      B  , , s���n. s���n� t���n� t���n. s���n.      B  , , v���n. v���n� w���n� w���n. v���n.      B  , , y���n. y���n� zp��n� zp��n. y���n.      B  , , |���n. |���n� }T��n� }T��n. |���n.      B  , , ���n. ���n� �8��n� �8��n. ���n.      B  , , �r��n. �r��n� ���n� ���n. �r��n.      B  , , �V��n. �V��n� � ��n� � ��n. �V��n.      B  , , �:��n. �:��n� ����n� ����n. �:��n.      B  , , v���k� v���l0 w���l0 w���k� v���k�      B  , , y���k� y���l0 zp��l0 zp��k� y���k�      B  , , |���k� |���l0 }T��l0 }T��k� |���k�      B  , , ���k� ���l0 �8��l0 �8��k� ���k�      B  , , �r��k� �r��l0 ���l0 ���k� �r��k�      B  , , �V��k� �V��l0 � ��l0 � ��k� �V��k�      B  , , �:��k� �:��l0 ����l0 ����k� �:��k�      B  , , ���j2 ���j� �8��j� �8��j2 ���j2      B  , , �r��j2 �r��j� ���j� ���j2 �r��j2      B  , , �V��j2 �V��j� � ��j� � ��j2 �V��j2      B  , , �:��j2 �:��j� ����j� ����j2 �:��j2      B  , , s���p� s���q� t���q� t���p� s���p�      B  , , v���p� v���q� w���q� w���p� v���p�      B  , , y���p� y���q� zp��q� zp��p� y���p�      B  , , |���p� |���q� }T��q� }T��p� |���p�      B  , , �V��o� �V��p, � ��p, � ��o� �V��o�      B  , , �:��o� �:��p, ����p, ����o� �:��o�      B  , , s���j2 s���j� t���j� t���j2 s���j2      B  , , v���j2 v���j� w���j� w���j2 v���j2      B  , , y���j2 y���j� zp��j� zp��j2 y���j2      B  , , |���j2 |���j� }T��j� }T��j2 |���j2      B  , , s���o� s���p, t���p, t���o� s���o�      B  , , v���o� v���p, w���p, w���o� v���o�      B  , , y���o� y���p, zp��p, zp��o� y���o�      B  , , s���l� s���m� t���m� t���l� s���l�      B  , , v���l� v���m� w���m� w���l� v���l�      B  , , y���l� y���m� zp��m� zp��l� y���l�      B  , , |���l� |���m� }T��m� }T��l� |���l�      B  , , ���l� ���m� �8��m� �8��l� ���l�      B  , , �r��l� �r��m� ���m� ���l� �r��l�      B  , , �V��l� �V��m� � ��m� � ��l� �V��l�      B  , , �:��l� �:��m� ����m� ����l� �:��l�      B  , , |���o� |���p, }T��p, }T��o� |���o�      B  , , ���p� ���q� �8��q� �8��p� ���p�      B  , , �r��p� �r��q� ���q� ���p� �r��p�      B  , , s���r* s���r� t���r� t���r* s���r*      B  , , v���r* v���r� w���r� w���r* v���r*      B  , , y���r* y���r� zp��r� zp��r* y���r*      B  , , ����r* ����r� �<��r� �<��r* ����r*      B  , , �v��r* �v��r� � ��r� � ��r* �v��r*      B  , , �Z��r* �Z��r� ���r� ���r* �Z��r*      B  , , ���j2 ���j� ����j� ����j2 ���j2      B  , , ���j2 ���j� ����j� ����j2 ���j2      B  , , ����j2 ����j� ����j� ����j2 ����j2      B  , , ����j2 ����j� �t��j� �t��j2 ����j2      B  , , ����j2 ����j� �X��j� �X��j2 ����j2      B  , , ����j2 ����j� �<��j� �<��j2 ����j2      B  , , �v��k� �v��l0 � ��l0 � ��k� �v��k�      B  , , �Z��k� �Z��l0 ���l0 ���k� �Z��k�      B  , , ���r* ���r� ����r� ����r* ���r*      B  , , ���r* ���r� ����r� ����r* ���r*      B  , , ���p� ���q� ����q� ����p� ���p�      B  , , ���p� ���q� ����q� ����p� ���p�      B  , , �v��j2 �v��j� � ��j� � ��j2 �v��j2      B  , , �Z��j2 �Z��j� ���j� ���j2 �Z��j2      B  , , ����p� ����q� ����q� ����p� ����p�      B  , , ���n. ���n� ����n� ����n. ���n.      B  , , ���o� ���p, ����p, ����o� ���o�      B  , , ���o� ���p, ����p, ����o� ���o�      B  , , ����o� ����p, ����p, ����o� ����o�      B  , , ����o� ����p, �t��p, �t��o� ����o�      B  , , ���n. ���n� ����n� ����n. ���n.      B  , , ����n. ����n� ����n� ����n. ����n.      B  , , ����n. ����n� �t��n� �t��n. ����n.      B  , , ����n. ����n� �X��n� �X��n. ����n.      B  , , �v��o� �v��p, � ��p, � ��o� �v��o�      B  , , �Z��o� �Z��p, ���p, ���o� �Z��o�      B  , , ����o� ����p, �X��p, �X��o� ����o�      B  , , ����o� ����p, �<��p, �<��o� ����o�      B  , , ����n. ����n� �<��n� �<��n. ����n.      B  , , �v��n. �v��n� � ��n� � ��n. �v��n.      B  , , �Z��n. �Z��n� ���n� ���n. �Z��n.      B  , , ����p� ����q� �t��q� �t��p� ����p�      B  , , ����p� ����q� �X��q� �X��p� ����p�      B  , , ����p� ����q� �<��q� �<��p� ����p�      B  , , �v��p� �v��q� � ��q� � ��p� �v��p�      B  , , �Z��p� �Z��q� ���q� ���p� �Z��p�      B  , , ����r* ����r� ����r� ����r* ����r*      B  , , ����r* ����r� �t��r� �t��r* ����r*      B  , , ���k� ���l0 ����l0 ����k� ���k�      B  , , ���l� ���m� ����m� ����l� ���l�      B  , , ���l� ���m� ����m� ����l� ���l�      B  , , ����l� ����m� ����m� ����l� ����l�      B  , , ����l� ����m� �t��m� �t��l� ����l�      B  , , ����l� ����m� �X��m� �X��l� ����l�      B  , , ����l� ����m� �<��m� �<��l� ����l�      B  , , �v��l� �v��m� � ��m� � ��l� �v��l�      B  , , �Z��l� �Z��m� ���m� ���l� �Z��l�      B  , , ���k� ���l0 ����l0 ����k� ���k�      B  , , ����k� ����l0 ����l0 ����k� ����k�      B  , , ����k� ����l0 �t��l0 �t��k� ����k�      B  , , ����k� ����l0 �X��l0 �X��k� ����k�      B  , , ����k� ����l0 �<��l0 �<��k� ����k�      B  , , ����r* ����r� �X��r� �X��r* ����r*      B  , , ����f6 ����f� �X��f� �X��f6 ����f6      B  , , ����f6 ����f� �<��f� �<��f6 ����f6      B  , , �v��f6 �v��f� � ��f� � ��f6 �v��f6      B  , , �Z��f6 �Z��f� ���f� ���f6 �Z��f6      B  , , �Z��g� �Z��h4 ���h4 ���g� �Z��g�      B  , , s���b: s���b� t���b� t���b: s���b:      B  , , v���b: v���b� w���b� w���b: v���b:      B  , , y���b: y���b� zp��b� zp��b: y���b:      B  , , |���b: |���b� }T��b� }T��b: |���b:      B  , , ���b: ���b� �8��b� �8��b: ���b:      B  , , �r��b: �r��b� ���b� ���b: �r��b:      B  , , �V��b: �V��b� � ��b� � ��b: �V��b:      B  , , �:��b: �:��b� ����b� ����b: �:��b:      B  , , ���b: ���b� ����b� ����b: ���b:      B  , , ���b: ���b� ����b� ����b: ���b:      B  , , ����b: ����b� ����b� ����b: ����b:      B  , , ����b: ����b� �t��b� �t��b: ����b:      B  , , ����b: ����b� �X��b� �X��b: ����b:      B  , , ����b: ����b� �<��b� �<��b: ����b:      B  , , �v��b: �v��b� � ��b� � ��b: �v��b:      B  , , �Z��b: �Z��b� ���b� ���b: �Z��b:      B  , , y���c� y���d8 zp��d8 zp��c� y���c�      B  , , |���c� |���d8 }T��d8 }T��c� |���c�      B  , , ���c� ���d8 �8��d8 �8��c� ���c�      B  , , �r��c� �r��d8 ���d8 ���c� �r��c�      B  , , �V��c� �V��d8 � ��d8 � ��c� �V��c�      B  , , s���f6 s���f� t���f� t���f6 s���f6      B  , , v���f6 v���f� w���f� w���f6 v���f6      B  , , y���f6 y���f� zp��f� zp��f6 y���f6      B  , , |���f6 |���f� }T��f� }T��f6 |���f6      B  , , ���f6 ���f� �8��f� �8��f6 ���f6      B  , , �r��f6 �r��f� ���f� ���f6 �r��f6      B  , , �V��f6 �V��f� � ��f� � ��f6 �V��f6      B  , , �:��c� �:��d8 ����d8 ����c� �:��c�      B  , , ���c� ���d8 ����d8 ����c� ���c�      B  , , ���c� ���d8 ����d8 ����c� ���c�      B  , , ����c� ����d8 ����d8 ����c� ����c�      B  , , ����c� ����d8 �t��d8 �t��c� ����c�      B  , , ����c� ����d8 �X��d8 �X��c� ����c�      B  , , ����c� ����d8 �<��d8 �<��c� ����c�      B  , , �v��c� �v��d8 � ��d8 � ��c� �v��c�      B  , , �Z��c� �Z��d8 ���d8 ���c� �Z��c�      B  , , s���d� s���e� t���e� t���d� s���d�      B  , , v���d� v���e� w���e� w���d� v���d�      B  , , y���d� y���e� zp��e� zp��d� y���d�      B  , , |���d� |���e� }T��e� }T��d� |���d�      B  , , ���d� ���e� �8��e� �8��d� ���d�      B  , , �r��d� �r��e� ���e� ���d� �r��d�      B  , , �V��d� �V��e� � ��e� � ��d� �V��d�      B  , , �:��d� �:��e� ����e� ����d� �:��d�      B  , , ���d� ���e� ����e� ����d� ���d�      B  , , ���d� ���e� ����e� ����d� ���d�      B  , , ����d� ����e� ����e� ����d� ����d�      B  , , ����d� ����e� �t��e� �t��d� ����d�      B  , , ����d� ����e� �X��e� �X��d� ����d�      B  , , ����d� ����e� �<��e� �<��d� ����d�      B  , , �v��d� �v��e� � ��e� � ��d� �v��d�      B  , , �Z��d� �Z��e� ���e� ���d� �Z��d�      B  , , s���c� s���d8 t���d8 t���c� s���c�      B  , , v���c� v���d8 w���d8 w���c� v���c�      B  , , s���g� s���h4 t���h4 t���g� s���g�      B  , , v���g� v���h4 w���h4 w���g� v���g�      B  , , y���g� y���h4 zp��h4 zp��g� y���g�      B  , , |���g� |���h4 }T��h4 }T��g� |���g�      B  , , ���g� ���h4 �8��h4 �8��g� ���g�      B  , , �r��g� �r��h4 ���h4 ���g� �r��g�      B  , , �V��g� �V��h4 � ��h4 � ��g� �V��g�      B  , , �:��g� �:��h4 ����h4 ����g� �:��g�      B  , , ���g� ���h4 ����h4 ����g� ���g�      B  , , ���g� ���h4 ����h4 ����g� ���g�      B  , , ����g� ����h4 ����h4 ����g� ����g�      B  , , ����g� ����h4 �t��h4 �t��g� ����g�      B  , , ����g� ����h4 �X��h4 �X��g� ����g�      B  , , ����g� ����h4 �<��h4 �<��g� ����g�      B  , , �v��g� �v��h4 � ��h4 � ��g� �v��g�      B  , , �:��f6 �:��f� ����f� ����f6 �:��f6      B  , , ���f6 ���f� ����f� ����f6 ���f6      B  , , ���f6 ���f� ����f� ����f6 ���f6      B  , , ����f6 ����f� ����f� ����f6 ����f6      B  , , ����f6 ����f� �t��f� �t��f6 ����f6      B  , , �^��d� �^��e� ���e� ���d� �^��d�      B  , , �B��d� �B��e� ����e� ����d� �B��d�      B  , , �^��b: �^��b� ���b� ���b: �^��b:      B  , , �B��b: �B��b� ����b� ����b: �B��b:      B  , , �&��b: �&��b� ����b� ����b: �&��b:      B  , , �
��b: �
��b� ´��b� ´��b: �
��b:      B  , , �&��d� �&��e� ����e� ����d� �&��d�      B  , , �
��d� �
��e� ´��e� ´��d� �
��d�      B  , , �^��g� �^��h4 ���h4 ���g� �^��g�      B  , , �B��g� �B��h4 ����h4 ����g� �B��g�      B  , , �&��g� �&��h4 ����h4 ����g� �&��g�      B  , , �
��g� �
��h4 ´��h4 ´��g� �
��g�      B  , , �^��f6 �^��f� ���f� ���f6 �^��f6      B  , , �B��f6 �B��f� ����f� ����f6 �B��f6      B  , , �&��f6 �&��f� ����f� ����f6 �&��f6      B  , , �
��f6 �
��f� ´��f� ´��f6 �
��f6      B  , , �^��c� �^��d8 ���d8 ���c� �^��c�      B  , , �B��c� �B��d8 ����d8 ����c� �B��c�      B  , , �&��c� �&��d8 ����d8 ����c� �&��c�      B  , , �
��c� �
��d8 ´��d8 ´��c� �
��c�      B  , , ����\T ����\� ����\� ����\T ����\T      B  , , ����\T ����\� �x��\� �x��\T ����\T      B  , , ����\T ����\� �\��\� �\��\T ����\T      B  , , ����\T ����\� �@��\� �@��\T ����\T      B  , , �z��\T �z��\� �$��\� �$��\T �z��\T      B  , , ����g� ����h4 �@��h4 �@��g� ����g�      B  , , �z��g� �z��h4 �$��h4 �$��g� �z��g�      B  , , �z��d� �z��e� �$��e� �$��d� �z��d�      B  , , �>��[  �>��[� ����[� ����[  �>��[       B  , , �"��[  �"��[� ����[� ����[  �"��[       B  , , ���[  ���[� ����[� ����[  ���[       B  , , ����[  ����[� ����[� ����[  ����[       B  , , ����[  ����[� �x��[� �x��[  ����[       B  , , ����[  ����[� �\��[� �\��[  ����[       B  , , ����[  ����[� �@��[� �@��[  ����[       B  , , �z��[  �z��[� �$��[� �$��[  �z��[       B  , , �>��\T �>��\� ����\� ����\T �>��\T      B  , , �"��\T �"��\� ����\� ����\T �"��\T      B  , , �>��b: �>��b� ����b� ����b: �>��b:      B  , , ����d� ����e� ����e� ����d� ����d�      B  , , ����d� ����e� �x��e� �x��d� ����d�      B  , , ����d� ����e� �\��e� �\��d� ����d�      B  , , �>��f6 �>��f� ����f� ����f6 �>��f6      B  , , �"��f6 �"��f� ����f� ����f6 �"��f6      B  , , ���f6 ���f� ����f� ����f6 ���f6      B  , , ����f6 ����f� ����f� ����f6 ����f6      B  , , ����f6 ����f� �x��f� �x��f6 ����f6      B  , , ����f6 ����f� �\��f� �\��f6 ����f6      B  , , ����f6 ����f� �@��f� �@��f6 ����f6      B  , , �z��f6 �z��f� �$��f� �$��f6 �z��f6      B  , , �"��b: �"��b� ����b� ����b: �"��b:      B  , , �>��d� �>��e� ����e� ����d� �>��d�      B  , , �"��d� �"��e� ����e� ����d� �"��d�      B  , , ���d� ���e� ����e� ����d� ���d�      B  , , ���b: ���b� ����b� ����b: ���b:      B  , , ����b: ����b� ����b� ����b: ����b:      B  , , �>��g� �>��h4 ����h4 ����g� �>��g�      B  , , �"��g� �"��h4 ����h4 ����g� �"��g�      B  , , ����b: ����b� �x��b� �x��b: ����b:      B  , , ���g� ���h4 ����h4 ����g� ���g�      B  , , ����g� ����h4 ����h4 ����g� ����g�      B  , , ����g� ����h4 �x��h4 �x��g� ����g�      B  , , ����g� ����h4 �\��h4 �\��g� ����g�      B  , , ����d� ����e� �@��e� �@��d� ����d�      B  , , �>��c� �>��d8 ����d8 ����c� �>��c�      B  , , �"��c� �"��d8 ����d8 ����c� �"��c�      B  , , ���c� ���d8 ����d8 ����c� ���c�      B  , , ����c� ����d8 ����d8 ����c� ����c�      B  , , ����c� ����d8 �x��d8 �x��c� ����c�      B  , , ����c� ����d8 �\��d8 �\��c� ����c�      B  , , ����c� ����d8 �@��d8 �@��c� ����c�      B  , , �z��c� �z��d8 �$��d8 �$��c� �z��c�      B  , , ����b: ����b� �\��b� �\��b: ����b:      B  , , ����b: ����b� �@��b� �@��b: ����b:      B  , , �z��b: �z��b� �$��b� �$��b: �z��b:      B  , , ���\T ���\� ����\� ����\T ���\T      B  , , ����Y� ����ZV �x��ZV �x��Y� ����Y�      B  , , ����Y� ����ZV �\��ZV �\��Y� ����Y�      B  , , ����Y� ����ZV �@��ZV �@��Y� ����Y�      B  , , �z��Y� �z��ZV �$��ZV �$��Y� �z��Y�      B  , , �>��Y� �>��ZV ����ZV ����Y� �>��Y�      B  , , �"��Y� �"��ZV ����ZV ����Y� �"��Y�      B  , , ���Y� ���ZV ����ZV ����Y� ���Y�      B  , , ����Y� ����ZV ����ZV ����Y� ����Y�      B  , , �>��XX �>��Y ����Y ����XX �>��XX      B  , , �"��XX �"��Y ����Y ����XX �"��XX      B  , , ���XX ���Y ����Y ����XX ���XX      B  , , ����XX ����Y ����Y ����XX ����XX      B  , , ����XX ����Y �x��Y �x��XX ����XX      B  , , ����XX ����Y �\��Y �\��XX ����XX      B  , , ����XX ����Y �@��Y �@��XX ����XX      B  , , �z��XX �z��Y �$��Y �$��XX �z��XX      B  , , �>��W �>��W� ����W� ����W �>��W      B  , , �"��W �"��W� ����W� ����W �"��W      B  , , ���W ���W� ����W� ����W ���W      B  , , ����W ����W� ����W� ����W ����W      B  , , ����W ����W� �x��W� �x��W ����W      B  , , ����W ����W� �\��W� �\��W ����W      B  , , ����W ����W� �@��W� �@��W ����W      B  , , �z��W �z��W� �$��W� �$��W �z��W      B  , , �>��U� �>��VZ ����VZ ����U� �>��U�      B  , , �"��U� �"��VZ ����VZ ����U� �"��U�      B  , , ���U� ���VZ ����VZ ����U� ���U�      B  , , ����U� ����VZ ����VZ ����U� ����U�      B  , , ����U� ����VZ �x��VZ �x��U� ����U�      B  , , ����U� ����VZ �\��VZ �\��U� ����U�      B  , , ����U� ����VZ �@��VZ �@��U� ����U�      B  , , �z��U� �z��VZ �$��VZ �$��U� �z��U�      B  , , �>��T\ �>��U ����U ����T\ �>��T\      B  , , �"��T\ �"��U ����U ����T\ �"��T\      B  , , ���T\ ���U ����U ����T\ ���T\      B  , , ����T\ ����U ����U ����T\ ����T\      B  , , ����T\ ����U �x��U �x��T\ ����T\      B  , , ����T\ ����U �\��U �\��T\ ����T\      B  , , ����T\ ����U �@��U �@��T\ ����T\      B  , , �z��T\ �z��U �$��U �$��T\ �z��T\      B  , , �>��S �>��S� ����S� ����S �>��S      B  , , �"��S �"��S� ����S� ����S �"��S      B  , , ���S ���S� ����S� ����S ���S      B  , , ����S ����S� ����S� ����S ����S      B  , , ����S ����S� �x��S� �x��S ����S      B  , , ����S ����S� �\��S� �\��S ����S      B  , , ����S ����S� �@��S� �@��S ����S      B  , , �z��S �z��S� �$��S� �$��S �z��S      B  , , �>��Q� �>��R^ ����R^ ����Q� �>��Q�      B  , , �"��Q� �"��R^ ����R^ ����Q� �"��Q�      B  , , ���Q� ���R^ ����R^ ����Q� ���Q�      B  , , ����Q� ����R^ ����R^ ����Q� ����Q�      B  , , ����Q� ����R^ �x��R^ �x��Q� ����Q�      B  , , ����Q� ����R^ �\��R^ �\��Q� ����Q�      B  , , ����Q� ����R^ �@��R^ �@��Q� ����Q�      B  , , �z��Q� �z��R^ �$��R^ �$��Q� �z��Q�      B  , , �>��P` �>��Q
 ����Q
 ����P` �>��P`      B  , , �"��P` �"��Q
 ����Q
 ����P` �"��P`      B  , , ���P` ���Q
 ����Q
 ����P` ���P`      B  , , ����P` ����Q
 ����Q
 ����P` ����P`      B  , , ����P` ����Q
 �x��Q
 �x��P` ����P`      B  , , ����P` ����Q
 �\��Q
 �\��P` ����P`      B  , , ����P` ����Q
 �@��Q
 �@��P` ����P`      B  , , �z��P` �z��Q
 �$��Q
 �$��P` �z��P`      B  , , �>��O �>��O� ����O� ����O �>��O      B  , , �"��O �"��O� ����O� ����O �"��O      B  , , ���O ���O� ����O� ����O ���O      B  , , ����O ����O� ����O� ����O ����O      B  , , ����O ����O� �x��O� �x��O ����O      B  , , ����O ����O� �\��O� �\��O ����O      B  , , ����O ����O� �@��O� �@��O ����O      B  , , �z��O �z��O� �$��O� �$��O �z��O      B  , , �>��M� �>��Nb ����Nb ����M� �>��M�      B  , , �"��M� �"��Nb ����Nb ����M� �"��M�      B  , , ���M� ���Nb ����Nb ����M� ���M�      B  , , ����M� ����Nb ����Nb ����M� ����M�      B  , , ����M� ����Nb �x��Nb �x��M� ����M�      B  , , ����M� ����Nb �\��Nb �\��M� ����M�      B  , , ����M� ����Nb �@��Nb �@��M� ����M�      B  , , �z��M� �z��Nb �$��Nb �$��M� �z��M�      B  , , �>��Ld �>��M ����M ����Ld �>��Ld      B  , , �"��Ld �"��M ����M ����Ld �"��Ld      B  , , ���Ld ���M ����M ����Ld ���Ld      B  , , ����Ld ����M ����M ����Ld ����Ld      B  , , ����Ld ����M �x��M �x��Ld ����Ld      B  , , ����Ld ����M �\��M �\��Ld ����Ld      B  , , ����Ld ����M �@��M �@��Ld ����Ld      B  , , �z��Ld �z��M �$��M �$��Ld �z��Ld      _   ,  �+  &�  �+  (<  �q  (<  �q  &�  �+  &�      _   ,  ��  &�  ��  (<  �w  (<  �w  &�  ��  &�      _   ,  �5  $�  �5  (7 -�  (7 -�  $�  �5  $�      _   , G�  $� G�  (7 ~0  (7 ~0  $� G�  $�      _   , �C  $� �C  (7 η  (7 η  $� �C  $�      _   ,  ^�  q  ^�  
�  �  
�  �  q  ^�  q      _   ,  ^����g  ^�����  �����  ����g  ^����g      _   ,  ^����]  ^�����  �����  ����]  ^����]      _   ,  ^����S  ^�����  �����  ����S  ^����S      _   ,  s���c�  s���g?  �=��g?  �=��c�  s���c�      _   , l��]� l��ac ���ac ���]� l��]�      _   , P��]� P��ac ���ac ���]� P��]�      _   , 4��]� 4��ac ���ac ���]� 4��]�      _   , 
��]� 
��ac ���ac ���]� 
��]�      _   , ���]� ���ac n��ac n��]� ���]�      _   , ���]� ���ac R��ac R��]� ���]�      _   , /���]� /���ac 1��ac 1��]� /���]�      _   , 2���]� 2���ac 4��ac 4��]� 2���]�      _   , 5t��]� 5t��ac 6���ac 6���]� 5t��]�      _   , 8X��]� 8X��ac 9���ac 9���]� 8X��]�      _   , ;<��]� ;<��ac <���ac <���]� ;<��]�      _   , > ��]� > ��ac ?���ac ?���]� > ��]�      _   , A��]� A��ac Bv��ac Bv��]� A��]�      _   , C���]� C���ac EZ��ac EZ��]� C���]�      _   , F���]� F���ac H>��ac H>��]� F���]�      _   , I���]� I���ac K"��ac K"��]� I���]�      _   , L���]� L���ac N��ac N��]� L���]�      _   , Ox��]� Ox��ac P���ac P���]� Ox��]�      _   , R\��]� R\��ac S���ac S���]� R\��]�      _   , U@��]� U@��ac V���ac V���]� U@��]�      _   , X$��]� X$��ac Y���ac Y���]� X$��]�      _   , [��]� [��ac \z��ac \z��]� [��]�      _   , ]���]� ]���ac _^��ac _^��]� ]���]�      _   , `���]� `���ac bB��ac bB��]� `���]�      _   , c���]� c���ac e&��ac e&��]� c���]�      _   , f���]� f���ac h
��ac h
��]� f���]�      C   , �  (� �  4: J  4: J  (� �  (�      C   , �  � �  #� J  #� J  � �  �      C   ,  [����5  [����  \b���  \b���5  [����5      C   ,  ]����^  ]����>  ^����>  ^����^  ]����^      C   ,  `@���^  `@���>  `����>  `����^  `@���^      C   ,  b����^  b����>  c8���>  c8���^  b����^      C   ,  d����^  d����>  e����>  e����^  d����^      C   ,  g*���^  g*���>  g����>  g����^  g*���^      C   ,  ix���^  ix���>  j"���>  j"���^  ix���^      C   ,  k����^  k����>  lp���>  lp���^  k����^      C   ,  n���^  n���>  n����>  n����^  n���^      C   ,  pb���^  pb���>  q���>  q���^  pb���^      C   ,  r����^  r����>  sZ���>  sZ���^  r����^      C   ,  t����^  t����>  u����>  u����^  t����^      C   ,  wL���^  wL���>  w����>  w����^  wL���^      C   ,  y����^  y����>  zD���>  zD���^  y����^      C   ,  {����^  {����>  |����>  |����^  {����^      C   ,  ~6���^  ~6���>  ~����>  ~����^  ~6���^      C   ,  �����^  �����>  �.���>  �.���^  �����^      C   ,  �����^  �����>  �|���>  �|���^  �����^      C   ,  � ���^  � ���>  �����>  �����^  � ���^      C   ,  �n���^  �n���>  ����>  ����^  �n���^      C   ,  �����^  �����>  �f���>  �f���^  �����^      C   ,  �
���^  �
���>  �����>  �����^  �
���^      C   ,  �X���^  �X���>  ����>  ����^  �X���^      C   ,  �����^  �����>  �P���>  �P���^  �����^      C   ,  �����^  �����>  �����>  �����^  �����^      C   ,  �B���^  �B���>  �����>  �����^  �B���^      C   ,  �����^  �����>  �:���>  �:���^  �����^      C   ,  �����^  �����>  �����>  �����^  �����^      C   ,  �,���^  �,���>  �����>  �����^  �,���^      C   ,  �z���^  �z���>  �$���>  �$���^  �z���^      C   ,  �����^  �����>  �r���>  �r���^  �����^      C   ,  ����^  ����>  �����>  �����^  ����^      C   ,  �d���^  �d���>  ����>  ����^  �d���^      C   ,  �����^  �����>  �\���>  �\���^  �����^      C   ,  � ���^  � ���>  �����>  �����^  � ���^      C   ,  �N���^  �N���>  �����>  �����^  �N���^      C   ,  �����^  �����>  �F���>  �F���^  �����^      C   ,  �����^  �����>  �����>  �����^  �����^      C   ,  �8���^  �8���>  �����>  �����^  �8���^      C   ,  �����^  �����>  �0���>  �0���^  �����^      C   ,  �����^  �����>  �~���>  �~���^  �����^      C   ,  �"���^  �"���>  �����>  �����^  �"���^      C   ,  �p���^  �p���>  ����>  ����^  �p���^      C   ,  �����^  �����>  �h���>  �h���^  �����^      C   ,  ����^  ����>  �����>  �����^  ����^      C   ,  �Z���^  �Z���>  ����>  ����^  �Z���^      C   ,  Ũ���^  Ũ���>  �R���>  �R���^  Ũ���^      C   ,  �����^  �����>  Ƞ���>  Ƞ���^  �����^      C   ,  �D���^  �D���>  �����>  �����^  �D���^      C   ,  ̒���^  ̒���>  �<���>  �<���^  ̒���^      C   ,  �����^  �����>  ϊ���>  ϊ���^  �����^      C   ,  �.���^  �.���>  �����>  �����^  �.���^      C   ,  �h���5  �h���  ����  ����5  �h���5      C   , F��a� F��s ���s ���a� F��a�      C   , F��L# F��]? ���]? ���L# F��L#      C   , ��  (� ��  4: ��  4: ��  (� ��  (�      C   , �(  (� �(  4: ��  4: ��  (� �(  (�      C   , �v  (� �v  4: �   4: �   (� �v  (�      C   , ��  (� ��  4: �n  4: �n  (� ��  (�      C   , �  (� �  4: ��  4: ��  (� �  (�      C   , �`  (� �`  4: �
  4: �
  (� �`  (�      C   , ��  (� ��  4: �X  4: �X  (� ��  (�      C   , ��  (� ��  4: ��  4: ��  (� ��  (�      C   , �J  (� �J  4: ��  4: ��  (� �J  (�      C   , Ř  (� Ř  4: �B  4: �B  (� Ř  (�      C   , ��  (� ��  4: Ȑ  4: Ȑ  (� ��  (�      C   , �4  (� �4  4: ��  4: ��  (� �4  (�      C   , ̂  (� ̂  4: �,  4: �,  (� ̂  (�      C   , ��  (� ��  4: �z  4: �z  (� ��  (�      C   , ��  3� ��  4{ �  4{ �  3� ��  3�      C   , ��  2_ ��  3	 �  3	 �  2_ ��  2_      C   , ��  0� ��  1� �  1� �  0� ��  0�      C   , ��  /{ ��  0% �  0% �  /{ ��  /{      C   , ��  .	 ��  .� �  .� �  .	 ��  .	      C   , ��  ,� ��  -A �  -A �  ,� ��  ,�      C   , ��  +% ��  +� �  +� �  +% ��  +%      C   , ��  )� ��  *] �  *] �  )� ��  )�      C   , ��  (A ��  (� �  (� �  (A ��  (A      C   , ��  ') ��  '� ��  '� ��  ') ��  ')      C   , ��  ') ��  '� �I  '� �I  ') ��  ')      C   , �M  ') �M  '� ��  '� ��  ') �M  ')      C   , ��  ') ��  '� ��  '� ��  ') ��  ')      C   , ��  ') ��  '� �3  '� �3  ') ��  ')      C   , �7  ') �7  '� ��  '� ��  ') �7  ')      C   , ��  ') ��  '� ��  '� ��  ') ��  ')      C   , ��  ') ��  '� �  '� �  ') ��  ')      C   , �!  ') �!  '� �k  '� �k  ') �!  ')      C   , �o  ') �o  '� ǹ  '� ǹ  ') �o  ')      C   , Ƚ  ') Ƚ  '� �  '� �  ') Ƚ  ')      C   , �  ') �  '� �U  '� �U  ') �  ')      C   , �Y  ') �Y  '� Σ  '� Σ  ') �Y  ')      C   , ��  &� ��  'y �  'y �  &� ��  &�      C   , ��  % ��  %� ��  %� ��  % ��  %      C   , ��  % ��  %� �I  %� �I  % ��  %      C   , �M  % �M  %� ��  %� ��  % �M  %      C   , ��  % ��  %� ��  %� ��  % ��  %      C   , ��  % ��  %� �3  %� �3  % ��  %      C   , �7  % �7  %� ��  %� ��  % �7  %      C   , ��  % ��  %� ��  %� ��  % ��  %      C   , ��  % ��  %� �  %� �  % ��  %      C   , �!  % �!  %� �k  %� �k  % �!  %      C   , �o  % �o  %� ǹ  %� ǹ  % �o  %      C   , Ƚ  % Ƚ  %� �  %� �  % Ƚ  %      C   , �  % �  %� �U  %� �U  % �  %      C   , �Y  % �Y  %� Σ  %� Σ  % �Y  %      C   , ��  %] ��  & �  & �  %] ��  %]      C   , ��  #� ��  $� �  $� �  #� ��  #�      C   , ��  � ��  #� ��  #� ��  � ��  �      C   , �(  � �(  #� ��  #� ��  � �(  �      C   , �v  � �v  #� �   #� �   � �v  �      C   , ��  � ��  #� �n  #� �n  � ��  �      C   , �  � �  #� ��  #� ��  � �  �      C   , �`  � �`  #� �
  #� �
  � �`  �      C   , ��  � ��  #� �X  #� �X  � ��  �      C   , ��  � ��  #� ��  #� ��  � ��  �      C   , �J  � �J  #� ��  #� ��  � �J  �      C   , Ř  � Ř  #� �B  #� �B  � Ř  �      C   , ��  � ��  #� Ȑ  #� Ȑ  � ��  �      C   , �4  � �4  #� ��  #� ��  � �4  �      C   , ̂  � ̂  #� �,  #� �,  � ̂  �      C   , ��  � ��  #� �z  #� �z  � ��  �      C   , ��  "y ��  ## �  ## �  "y ��  "y      C   , ��  ! ��  !� �  !� �  ! ��  !      C   , ��  � ��   ? �   ? �  � ��  �      C   , ��  # ��  � �  � �  # ��  #      C   , ��  � ��  [ �  [ �  � ��  �      C   , ��  ? ��  � �  � �  ? ��  ?      C   , ��  � ��  w �  w �  � ��  �      C   , ��  [ ��   �   �  [ ��  [      C   , ��  ') ��  '� �  '� �  ') ��  ')      C   , �  ') �  '� �_  '� �_  ') �  ')      C   , �c  ') �c  '� ��  '� ��  ') �c  ')      C   , �^  #� �^  $� �  $� �  #� �^  #�      C   , �^  %] �^  & �  & �  %] �^  %]      C   , �^  "y �^  ## �  ## �  "y �^  "y      C   , �^  ! �^  !� �  !� �  ! �^  !      C   , �^  � �^   ? �   ? �  � �^  �      C   , �^  # �^  � �  � �  # �^  #      C   , �^  � �^  [ �  [ �  � �^  �      C   , �^  ? �^  � �  � �  ? �^  ?      C   , �^  � �^  w �  w �  � �^  �      C   , �^  [ �^   �   �  [ �^  [      C   , �2  � �2  #� ��  #� ��  � �2  �      C   , ��  � ��  #� �*  #� �*  � ��  �      C   , ��  � ��  #� �x  #� �x  � ��  �      C   , �  � �  #� ��  #� ��  � �  �      C   , �j  � �j  #� �  #� �  � �j  �      C   , ��  � ��  #� �b  #� �b  � ��  �      C   , �  � �  #� ��  #� ��  � �  �      C   , �T  � �T  #� ��  #� ��  � �T  �      C   , ��  � ��  #� �L  #� �L  � ��  �      C   , ��  � ��  #� ��  #� ��  � ��  �      C   , �>  � �>  #� ��  #� ��  � �>  �      C   , ��  � ��  #� �6  #� �6  � ��  �      C   , �k  % �k  %� ��  %� ��  % �k  %      C   , ��  % ��  %� ��  %� ��  % ��  %      C   , ��  % ��  %� �=  %� �=  % ��  %      C   , �A  % �A  %� ��  %� ��  % �A  %      C   , ��  % ��  %� ��  %� ��  % ��  %      C   , ��  % ��  %� �'  %� �'  % ��  %      C   , �+  % �+  %� �u  %� �u  % �+  %      C   , �y  % �y  %� ��  %� ��  % �y  %      C   , ��  % ��  %� �  %� �  % ��  %      C   , �  % �  %� �_  %� �_  % �  %      C   , �c  % �c  %� ��  %� ��  % �c  %      C   , �^  (A �^  (� �  (� �  (A �^  (A      C   , ��  (� ��  4: �6  4: �6  (� ��  (�      C   , �^  &� �^  'y �  'y �  &� �^  &�      C   , �k  ') �k  '� ��  '� ��  ') �k  ')      C   , ��  ') ��  '� ��  '� ��  ') ��  ')      C   , ��  ') ��  '� �=  '� �=  ') ��  ')      C   , �A  ') �A  '� ��  '� ��  ') �A  ')      C   , ��  ') ��  '� ��  '� ��  ') ��  ')      C   , ��  ') ��  '� �'  '� �'  ') ��  ')      C   , �+  ') �+  '� �u  '� �u  ') �+  ')      C   , �y  ') �y  '� ��  '� ��  ') �y  ')      C   , �^  3� �^  4{ �  4{ �  3� �^  3�      C   , �^  2_ �^  3	 �  3	 �  2_ �^  2_      C   , �^  0� �^  1� �  1� �  0� �^  0�      C   , �^  /{ �^  0% �  0% �  /{ �^  /{      C   , �^  .	 �^  .� �  .� �  .	 �^  .	      C   , �^  ,� �^  -A �  -A �  ,� �^  ,�      C   , �^  +% �^  +� �  +� �  +% �^  +%      C   , �^  )� �^  *] �  *] �  )� �^  )�      C   , ��  (� ��  4: �x  4: �x  (� ��  (�      C   , �  (� �  4: ��  4: ��  (� �  (�      C   , �j  (� �j  4: �  4: �  (� �j  (�      C   , ��  (� ��  4: �b  4: �b  (� ��  (�      C   , �  (� �  4: ��  4: ��  (� �  (�      C   , �T  (� �T  4: ��  4: ��  (� �T  (�      C   , ��  (� ��  4: �L  4: �L  (� ��  (�      C   , ��  (� ��  4: ��  4: ��  (� ��  (�      C   , �>  (� �>  4: ��  4: ��  (� �>  (�      C   , N�  % N�  %� P  %� P  % N�  %      C   , N�  ') N�  '� P  '� P  ') N�  ')      C   , Z@  ') Z@  '� [�  '� [�  ') Z@  ')      C   , \�  ') \�  '� ]�  '� ]�  ') \�  ')      C   , ^�  ') ^�  '� `&  '� `&  ') ^�  ')      C   , a*  ') a*  '� bt  '� bt  ') a*  ')      C   , P1  � P1  #� P�  #� P�  � P1  �      C   , R  � R  #� S)  #� S)  � R  �      C   , T�  � T�  #� Uw  #� Uw  � T�  �      C   , W  � W  #� W�  #� W�  � W  �      C   , Yi  � Yi  #� Z  #� Z  � Yi  �      C   , [�  � [�  #� \a  #� \a  � [�  �      C   , ^  � ^  #� ^�  #� ^�  � ^  �      C   , `S  � `S  #� `�  #� `�  � `S  �      C   , b�  � b�  #� cK  #� cK  � b�  �      C   , d�  � d�  #� e�  #� e�  � d�  �      C   , g=  � g=  #� g�  #� g�  � g=  �      C   , i�  � i�  #� j5  #� j5  � i�  �      C   , k�  � k�  #� l�  #� l�  � k�  �      C   , n'  � n'  #� n�  #� n�  � n'  �      C   , pu  � pu  #� q  #� q  � pu  �      C   , r�  � r�  #� sm  #� sm  � r�  �      C   , u  � u  #� u�  #� u�  � u  �      C   , w_  � w_  #� x	  #� x	  � w_  �      C   , y�  � y�  #� zW  #� zW  � y�  �      C   , {�  � {�  #� |�  #� |�  � {�  �      C   , ~I  � ~I  #� ~�  #� ~�  � ~I  �      C   , cx  ') cx  '� d�  '� d�  ') cx  ')      C   , e�  ') e�  '� g  '� g  ') e�  ')      C   , h  ') h  '� i^  '� i^  ') h  ')      C   , jb  ') jb  '� k�  '� k�  ') jb  ')      C   , l�  ') l�  '� m�  '� m�  ') l�  ')      C   , U�  ') U�  '� V�  '� V�  ') U�  ')      C   , Q  % Q  %� RR  %� RR  % Q  %      C   , SV  % SV  %� T�  %� T�  % SV  %      C   , U�  % U�  %� V�  %� V�  % U�  %      C   , W�  % W�  %� Y<  %� Y<  % W�  %      C   , Z@  % Z@  %� [�  %� [�  % Z@  %      C   , \�  % \�  %� ]�  %� ]�  % \�  %      C   , ^�  % ^�  %� `&  %� `&  % ^�  %      C   , a*  % a*  %� bt  %� bt  % a*  %      C   , cx  % cx  %� d�  %� d�  % cx  %      C   , e�  % e�  %� g  %� g  % e�  %      C   , h  % h  %� i^  %� i^  % h  %      C   , jb  % jb  %� k�  %� k�  % jb  %      C   , l�  % l�  %� m�  %� m�  % l�  %      C   , n�  % n�  %� pH  %� pH  % n�  %      C   , qL  % qL  %� r�  %� r�  % qL  %      C   , s�  % s�  %� t�  %� t�  % s�  %      C   , u�  % u�  %� w2  %� w2  % u�  %      C   , x6  % x6  %� y�  %� y�  % x6  %      C   , z�  % z�  %� {�  %� {�  % z�  %      C   , |�  % |�  %� ~  %� ~  % |�  %      C   , n�  ') n�  '� pH  '� pH  ') n�  ')      C   , qL  ') qL  '� r�  '� r�  ') qL  ')      C   , s�  ') s�  '� t�  '� t�  ') s�  ')      C   , u�  ') u�  '� w2  '� w2  ') u�  ')      C   , x6  ') x6  '� y�  '� y�  ') x6  ')      C   , P1  (� P1  4: P�  4: P�  (� P1  (�      C   , R  (� R  4: S)  4: S)  (� R  (�      C   , T�  (� T�  4: Uw  4: Uw  (� T�  (�      C   , W  (� W  4: W�  4: W�  (� W  (�      C   , Yi  (� Yi  4: Z  4: Z  (� Yi  (�      C   , [�  (� [�  4: \a  4: \a  (� [�  (�      C   , ^  (� ^  4: ^�  4: ^�  (� ^  (�      C   , `S  (� `S  4: `�  4: `�  (� `S  (�      C   , b�  (� b�  4: cK  4: cK  (� b�  (�      C   , d�  (� d�  4: e�  4: e�  (� d�  (�      C   , g=  (� g=  4: g�  4: g�  (� g=  (�      C   , i�  (� i�  4: j5  4: j5  (� i�  (�      C   , k�  (� k�  4: l�  4: l�  (� k�  (�      C   , n'  (� n'  4: n�  4: n�  (� n'  (�      C   , pu  (� pu  4: q  4: q  (� pu  (�      C   , r�  (� r�  4: sm  4: sm  (� r�  (�      C   , u  (� u  4: u�  4: u�  (� u  (�      C   , w_  (� w_  4: x	  4: x	  (� w_  (�      C   , y�  (� y�  4: zW  4: zW  (� y�  (�      C   , {�  (� {�  4: |�  4: |�  (� {�  (�      C   , ~I  (� ~I  4: ~�  4: ~�  (� ~I  (�      C   , z�  ') z�  '� {�  '� {�  ') z�  ')      C   , |�  ') |�  '� ~  '� ~  ') |�  ')      C   , W�  ') W�  '� Y<  '� Y<  ') W�  ')      C   , Q  ') Q  '� RR  '� RR  ') Q  ')      C   , SV  ') SV  '� T�  '� T�  ') SV  ')      C   , �  (� �  4:  �  4:  �  (� �  (�      C   , �  � �  #�  �  #�  �  � �  �      C   , "<  � "<  #� "�  #� "�  � "<  �      C   , w  % w  %� �  %� �  % w  %      C   ,  �  %  �  %� "  %� "  %  �  %      C   , #  % #  %� $]  %� $]  % #  %      C   , %a  % %a  %� &�  %� &�  % %a  %      C   , "<  (� "<  4: "�  4: "�  (� "<  (�      C   , $�  (� $�  4: %4  4: %4  (� $�  (�      C   , &�  (� &�  4: '�  4: '�  (� &�  (�      C   , )&  (� )&  4: )�  4: )�  (� )&  (�      C   , +t  (� +t  4: ,  4: ,  (� +t  (�      C   , -�  (� -�  4: .l  4: .l  (� -�  (�      C   , 1�  3� 1�  4{ @�  4{ @�  3� 1�  3�      C   , 1�  2_ 1�  3	 @�  3	 @�  2_ 1�  2_      C   , 1�  0� 1�  1� @�  1� @�  0� 1�  0�      C   , 1�  /{ 1�  0% @�  0% @�  /{ 1�  /{      C   , 1�  .	 1�  .� @�  .� @�  .	 1�  .	      C   , 1�  ,� 1�  -A @�  -A @�  ,� 1�  ,�      C   , 1�  +% 1�  +� @�  +� @�  +% 1�  +%      C   , 1�  )� 1�  *] @�  *] @�  )� 1�  )�      C   , IG  (� IG  4: I�  4: I�  (� IG  (�      C   , K�  (� K�  4: L?  4: L?  (� K�  (�      C   , M�  (� M�  4: N�  4: N�  (� M�  (�      C   , '�  % '�  %� (�  %� (�  % '�  %      C   , )�  % )�  %� +G  %� +G  % )�  %      C   , ,K  % ,K  %� -�  %� -�  % ,K  %      C   , 1�  %] 1�  & @�  & @�  %] 1�  %]      C   , G�  % G�  %� I  %� I  % G�  %      C   , J  % J  %� Kh  %� Kh  % J  %      C   , Ll  % Ll  %� M�  %� M�  % Ll  %      C   , $�  � $�  #� %4  #� %4  � $�  �      C   , &�  � &�  #� '�  #� '�  � &�  �      C   , )&  � )&  #� )�  #� )�  � )&  �      C   , +t  � +t  #� ,  #� ,  � +t  �      C   , -�  � -�  #� .l  #� .l  � -�  �      C   , 1�  "y 1�  ## @�  ## @�  "y 1�  "y      C   , 1�  ! 1�  !� @�  !� @�  ! 1�  !      C   , 1�  � 1�   ? @�   ? @�  � 1�  �      C   , 1�  # 1�  � @�  � @�  # 1�  #      C   , 1�  � 1�  [ @�  [ @�  � 1�  �      C   , 1�  ? 1�  � @�  � @�  ? 1�  ?      C   , 1�  � 1�  w @�  w @�  � 1�  �      C   , 1�  [ 1�   @�   @�  [ 1�  [      C   , D�  � D�  #� EU  #� EU  � D�  �      C   , F�  � F�  #� G�  #� G�  � F�  �      C   , IG  � IG  #� I�  #� I�  � IG  �      C   , 1�  (A 1�  (� @�  (� @�  (A 1�  (A      C   , w  ') w  '� �  '� �  ') w  ')      C   ,  �  ')  �  '� "  '� "  ')  �  ')      C   , #  ') #  '� $]  '� $]  ') #  ')      C   , %a  ') %a  '� &�  '� &�  ') %a  ')      C   , '�  ') '�  '� (�  '� (�  ') '�  ')      C   , )�  ') )�  '� +G  '� +G  ') )�  ')      C   , ,K  ') ,K  '� -�  '� -�  ') ,K  ')      C   , 1�  &� 1�  'y @�  'y @�  &� 1�  &�      C   , G�  ') G�  '� I  '� I  ') G�  ')      C   , J  ') J  '� Kh  '� Kh  ') J  ')      C   , Ll  ') Ll  '� M�  '� M�  ') Ll  ')      C   , K�  � K�  #� L?  #� L?  � K�  �      C   , M�  � M�  #� N�  #� N�  � M�  �      C   , 1�  #� 1�  $� @�  $� @�  #� 1�  #�      C   ,  ��  	�  ��  
�  �C  
�  �C  	�  ��  	�      C   ,  ��  �  ��    �C    �C  �  ��  �      C   ,  �h���I  �h  '  �  '  ����I  �h���I      C   ,  [�����  [����I  ����I  �����  [�����      C   ,  \�����  \�����  ������  ������  \�����      C   ,  \����/  \�����  ������  �����/  \����/      C   ,  [����  [�����  �����  ����  [����      C   ,  ������  �����  �C���  �C����  ������      C   ,  ������  �����u  �C���u  �C����  ������      C   ,  [���ϕ  [����?  ����?  ���ϕ  [���ϕ      C   ,  \�����  \���·  ����·  ������  \�����      C   ,  \����%  \�����  ������  �����%  \����%      C   ,  [����  [���ʽ  ���ʽ  ����  [����      C   ,  ]H  �  ]H  �  ҂  �  ҂  �  ]H  �      C   ,  [�  '  [�  �  �  �  �  '  [�  '      C   ,  [����I  [�  '  \b  '  \b���I  [����I      C   ,  �$  �  �$  #�  ��  #�  ��  �  �$  �      C   ,  �r  �  �r  #�  �  #�  �  �  �r  �      C   ,  ��  �  ��  #�  �j  #�  �j  �  ��  �      C   ,  �  �  �  #�  ��  #�  ��  �  �  �      C   ,  �\  �  �\  #�  �  #�  �  �  �\  �      C   ,  ��  �  ��  #�  T  #�  T  �  ��  �      C   , �  � �  #� �  #� �  � �  �      C   , F  � F  #� �  #� �  � F  �      C   , �  � �  #� >  #� >  � �  �      C   , �  � �  #� 	�  #� 	�  � �  �      C   , 0  � 0  #� �  #� �  � 0  �      C   , ~  � ~  #� (  #� (  � ~  �      C   , �  � �  #� v  #� v  � �  �      C   ,   �   #� �  #� �  �   �      C   , h  � h  #�   #�   � h  �      C   , �  � �  #� `  #� `  � �  �      C   ,   �   #� �  #� �  �   �      C   , R  � R  #� �  #� �  � R  �      C   ,  �]  %  �]  %�  �  %�  �  %  �]  %      C   ,  ��  %  ��  %�  ��  %�  ��  %  ��  %      C   ,  ��  %  ��  %�  �/  %�  �/  %  ��  %      C   ,  �3  %  �3  %�  �}  %�  �}  %  �3  %      C   ,  �  %  �  %� �  %� �  %  �  %      C   , �  % �  %�   %�   % �  %      C   ,   %   %� g  %� g  %   %      C   , k  % k  %� �  %� �  % k  %      C   , 	�  % 	�  %�   %�   % 	�  %      C   ,   %   %� Q  %� Q  %   %      C   , U  % U  %� �  %� �  % U  %      C   , �  % �  %� �  %� �  % �  %      C   , �  % �  %� ;  %� ;  % �  %      C   , ?  % ?  %� �  %� �  % ?  %      C   , �  % �  %� �  %� �  % �  %      C   , �  % �  %� %  %� %  % �  %      C   , )  % )  %� s  %� s  % )  %      C   ,  �]  ')  �]  '�  �  '�  �  ')  �]  ')      C   ,  ��  ')  ��  '�  ��  '�  ��  ')  ��  ')      C   ,  ��  ')  ��  '�  �/  '�  �/  ')  ��  ')      C   ,  �3  ')  �3  '�  �}  '�  �}  ')  �3  ')      C   ,  �  ')  �  '� �  '� �  ')  �  ')      C   , �  ') �  '�   '�   ') �  ')      C   ,   ')   '� g  '� g  ')   ')      C   , k  ') k  '� �  '� �  ') k  ')      C   , 	�  ') 	�  '�   '�   ') 	�  ')      C   ,   ')   '� Q  '� Q  ')   ')      C   , U  ') U  '� �  '� �  ') U  ')      C   , �  ') �  '� �  '� �  ') �  ')      C   , �  ') �  '� ;  '� ;  ') �  ')      C   , ?  ') ?  '� �  '� �  ') ?  ')      C   , �  ') �  '� �  '� �  ') �  ')      C   , �  ') �  '� %  '� %  ') �  ')      C   , )  ') )  '� s  '� s  ') )  ')      C   ,   (�   4: �  4: �  (�   (�      C   , R  (� R  4: �  4: �  (� R  (�      C   ,  ��  (�  ��  4:  �j  4:  �j  (�  ��  (�      C   ,  �  (�  �  4:  ��  4:  ��  (�  �  (�      C   ,  �\  (�  �\  4:  �  4:  �  (�  �\  (�      C   ,  ��  (�  ��  4:  T  4:  T  (�  ��  (�      C   , �  (� �  4: �  4: �  (� �  (�      C   , F  (� F  4: �  4: �  (� F  (�      C   , �  (� �  4: >  4: >  (� �  (�      C   , �  (� �  4: 	�  4: 	�  (� �  (�      C   , 0  (� 0  4: �  4: �  (� 0  (�      C   , ~  (� ~  4: (  4: (  (� ~  (�      C   , �  (� �  4: v  4: v  (� �  (�      C   ,   (�   4: �  4: �  (�   (�      C   , h  (� h  4:   4:   (� h  (�      C   , �  (� �  4: `  4: `  (� �  (�      C   ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      C   ,  ��  '.  ��  '�  �  '�  �  '.  ��  '.      C   ,  �  '.  �  '�  �c  '�  �c  '.  �  '.      C   ,  ��  '.  ��  '�  �+  '�  �+  '.  ��  '.      C   ,  �/  '.  �/  '�  �y  '�  �y  '.  �/  '.      C   ,  �}  '.  �}  '�  ��  '�  ��  '.  �}  '.      C   ,  Ϸ  	�  Ϸ  
�  �  
�  �  	�  Ϸ  	�      C   ,  �  r  �  R  ��  R  ��  r  �  r      C   ,  �G  �  �G    ��    ��  �  �G  �      C   ,  ��  �  ��    ��    ��  �  ��  �      C   ,  ��  �  ��    �-    �-  �  ��  �      C   ,  �1  �  �1    �{    �{  �  �1  �      C   ,  �  �  �    ��    ��  �  �  �      C   ,  ��  �  ��    �    �  �  ��  �      C   ,  �  �  �    �e    �e  �  �  �      C   ,  �i  �  �i    γ    γ  �  �i  �      C   ,  Ϸ  �  Ϸ    �    �  �  Ϸ  �      C   ,  �p���  �p  �  �  �  ����  �p���      C   ,  �����  ��  �  �h  �  �h���  �����      C   ,  ����  �  �  ��  �  �����  ����      C   ,  �Z���  �Z  �  �  �  ����  �Z���      C   ,  Ũ���  Ũ  �  �R  �  �R���  Ũ���      C   ,  �����  ��  �  Ƞ  �  Ƞ���  �����      C   ,  �D���  �D  �  ��  �  �����  �D���      C   ,  ̒���  ̒  �  �<  �  �<���  ̒���      C   ,  �����  ��  �  ϊ  �  ϊ���  �����      C   ,  �.���  �.  �  ��  �  �����  �.���      C   ,  �Z  r  �Z  R  �  R  �  r  �Z  r      C   ,  �  	�  �  
�  �e  
�  �e  	�  �  	�      C   ,  �i  	�  �i  
�  γ  
�  γ  	�  �i  	�      C   ,  Ũ  r  Ũ  R  �R  R  �R  r  Ũ  r      C   ,  ��  r  ��  R  Ƞ  R  Ƞ  r  ��  r      C   ,  �D  r  �D  R  ��  R  ��  r  �D  r      C   ,  ̒  r  ̒  R  �<  R  �<  r  ̒  r      C   ,  ��  r  ��  R  ϊ  R  ϊ  r  ��  r      C   ,  �.  r  �.  R  ��  R  ��  r  �.  r      C   ,  ��  r  ��  R  �h  R  �h  r  ��  r      C   ,  �G  	�  �G  
�  ��  
�  ��  	�  �G  	�      C   ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C   ,  ��  	�  ��  
�  �-  
�  �-  	�  ��  	�      C   ,  �1  	�  �1  
�  �{  
�  �{  	�  �1  	�      C   ,  �  	�  �  
�  ��  
�  ��  	�  �  	�      C   ,  ��  	�  ��  
�  �  
�  �  	�  ��  	�      C   ,  �p  r  �p  R  �  R  �  r  �p  r      C   ,  ��  �  ��    ��    ��  �  ��  �      C   ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C   ,  �  '.  �  '�  �]  '�  �]  '.  �  '.      C   ,  ��  '.  ��  '�  �  '�  �  '.  ��  '.      C   ,  �#  '.  �#  '�  �m  '�  �m  '.  �#  '.      C   ,  �q  '.  �q  '�  ��  '�  ��  '.  �q  '.      C   ,  ��  '.  ��  '�  �	  '�  �	  '.  ��  '.      C   ,  �  '.  �  '�  �W  '�  �W  '.  �  '.      C   ,  �[  '.  �[  '�  ��  '�  ��  '.  �[  '.      C   ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      C   ,  ��  '.  ��  '�  �A  '�  �A  '.  ��  '.      C   ,  �E  '.  �E  '�  ��  '�  ��  '.  �E  '.      C   ,  �w  '.  �w  '�  ��  '�  ��  '.  �w  '.      C   ,  ��  '.  ��  '�  �  '�  �  '.  ��  '.      C   ,  ��  '.  ��  '�  �O  '�  �O  '.  ��  '.      C   ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      C   ,  �A  '.  �A  '�  ��  '�  ��  '.  �A  '.      C   ,  �?  '.  �?  '�  ��  '�  ��  '.  �?  '.      C   ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      C   ,  ��  '.  ��  '�  �%  '�  �%  '.  ��  '.      C   ,  �)  '.  �)  '�  �s  '�  �s  '.  �)  '.      C   ,  g�  '.  g�  '�  h�  '�  h�  '.  g�  '.      C   ,  j;  '.  j;  '�  j�  '�  j�  '.  j;  '.      C   ,  l�  '.  l�  '�  m3  '�  m3  '.  l�  '.      C   ,  n�  '.  n�  '�  o�  '�  o�  '.  n�  '.      C   ,  q%  '.  q%  '�  q�  '�  q�  '.  q%  '.      C   ,  ss  '.  ss  '�  t  '�  t  '.  ss  '.      C   ,  u�  '.  u�  '�  vk  '�  vk  '.  u�  '.      C   ,  x  '.  x  '�  x�  '�  x�  '.  x  '.      C   ,  z]  '.  z]  '�  {  '�  {  '.  z]  '.      C   ,  ��  '.  ��  '�  �e  '�  �e  '.  ��  '.      C   ,  �	  '.  �	  '�  ��  '�  ��  '.  �	  '.      C   ,  �W  '.  �W  '�  �  '�  �  '.  �W  '.      C   ,  ��  (�  ��  4?  �>  4?  �>  (�  ��  (�      C   ,  Z  '.  Z  '�  Z�  '�  Z�  '.  Z  '.      C   ,  \g  '.  \g  '�  ]  '�  ]  '.  \g  '.      C   ,  ^�  '.  ^�  '�  __  '�  __  '.  ^�  '.      C   ,  a  '.  a  '�  a�  '�  a�  '.  a  '.      C   ,  cQ  '.  cQ  '�  c�  '�  c�  '.  cQ  '.      C   ,  e�  '.  e�  '�  fI  '�  fI  '.  e�  '.      C   ,  ��  �  ��    �A    �A  �  ��  �      C   ,  �E  �  �E    ��    ��  �  �E  �      C   ,  a  	�  a  
�  ba  
�  ba  	�  a  	�      C   ,  u�  	�  u�  
�  w  
�  w  	�  u�  	�      C   ,  ce  	�  ce  
�  d�  
�  d�  	�  ce  	�      C   ,  x#  	�  x#  
�  ym  
�  ym  	�  x#  	�      C   ,  zq  	�  zq  
�  {�  
�  {�  	�  zq  	�      C   ,  |�  	�  |�  
�  ~	  
�  ~	  	�  |�  	�      C   ,    	�    
�  �W  
�  �W  	�    	�      C   ,  �[  	�  �[  
�  ��  
�  ��  	�  �[  	�      C   ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C   ,  ��  	�  ��  
�  �A  
�  �A  	�  ��  	�      C   ,  �E  	�  �E  
�  ��  
�  ��  	�  �E  	�      C   ,  e�  	�  e�  
�  f�  
�  f�  	�  e�  	�      C   ,  ]����  ]�  �  ^�  �  ^����  ]����      C   ,  `@���  `@  �  `�  �  `����  `@���      C   ,  b����  b�  �  c8  �  c8���  b����      C   ,  d����  d�  �  e�  �  e����  d����      C   ,  g*���  g*  �  g�  �  g����  g*���      C   ,  h  	�  h  
�  iK  
�  iK  	�  h  	�      C   ,  jO  	�  jO  
�  k�  
�  k�  	�  jO  	�      C   ,  l�  	�  l�  
�  m�  
�  m�  	�  l�  	�      C   ,  n�  	�  n�  
�  p5  
�  p5  	�  n�  	�      C   ,  q9  	�  q9  
�  r�  
�  r�  	�  q9  	�      C   ,  �����  ��  �  �f  �  �f���  �����      C   ,  ^�  	�  ^�  
�  `  
�  `  	�  ^�  	�      C   ,  s�  	�  s�  
�  t�  
�  t�  	�  s�  	�      C   ,  ^�  �  ^�    `    `  �  ^�  �      C   ,  a  �  a    ba    ba  �  a  �      C   ,  ce  �  ce    d�    d�  �  ce  �      C   ,  e�  �  e�    f�    f�  �  e�  �      C   ,  h  �  h    iK    iK  �  h  �      C   ,  jO  �  jO    k�    k�  �  jO  �      C   ,  l�  �  l�    m�    m�  �  l�  �      C   ,  ix���  ix  �  j"  �  j"���  ix���      C   ,  k����  k�  �  lp  �  lp���  k����      C   ,  n���  n  �  n�  �  n����  n���      C   ,  pb���  pb  �  q  �  q���  pb���      C   ,  r����  r�  �  sZ  �  sZ���  r����      C   ,  t����  t�  �  u�  �  u����  t����      C   ,  wL���  wL  �  w�  �  w����  wL���      C   ,  y����  y�  �  zD  �  zD���  y����      C   ,  {����  {�  �  |�  �  |����  {����      C   ,  ~6���  ~6  �  ~�  �  ~����  ~6���      C   ,  n�  �  n�    p5    p5  �  n�  �      C   ,  q9  �  q9    r�    r�  �  q9  �      C   ,  s�  �  s�    t�    t�  �  s�  �      C   ,  u�  �  u�    w    w  �  u�  �      C   ,  x#  �  x#    ym    ym  �  x#  �      C   ,  zq  �  zq    {�    {�  �  zq  �      C   ,  |�  �  |�    ~	    ~	  �  |�  �      C   ,    �      �W    �W  �    �      C   ,  �[  �  �[    ��    ��  �  �[  �      C   ,  ��  �  ��    ��    ��  �  ��  �      C   ,  �����  ��  �  �.  �  �.���  �����      C   ,  �����  ��  �  �|  �  �|���  �����      C   ,  � ���  �   �  ��  �  �����  � ���      C   ,  ]�  r  ]�  R  ^�  R  ^�  r  ]�  r      C   ,  `@  r  `@  R  `�  R  `�  r  `@  r      C   ,  b�  r  b�  R  c8  R  c8  r  b�  r      C   ,  d�  r  d�  R  e�  R  e�  r  d�  r      C   ,  g*  r  g*  R  g�  R  g�  r  g*  r      C   ,  ix  r  ix  R  j"  R  j"  r  ix  r      C   ,  k�  r  k�  R  lp  R  lp  r  k�  r      C   ,  n  r  n  R  n�  R  n�  r  n  r      C   ,  pb  r  pb  R  q  R  q  r  pb  r      C   ,  r�  r  r�  R  sZ  R  sZ  r  r�  r      C   ,  t�  r  t�  R  u�  R  u�  r  t�  r      C   ,  wL  r  wL  R  w�  R  w�  r  wL  r      C   ,  y�  r  y�  R  zD  R  zD  r  y�  r      C   ,  {�  r  {�  R  |�  R  |�  r  {�  r      C   ,  ~6  r  ~6  R  ~�  R  ~�  r  ~6  r      C   ,  ��  r  ��  R  �.  R  �.  r  ��  r      C   ,  ��  r  ��  R  �|  R  �|  r  ��  r      C   ,  �   r  �   R  ��  R  ��  r  �   r      C   ,  �n  r  �n  R  �  R  �  r  �n  r      C   ,  ��  r  ��  R  �f  R  �f  r  ��  r      C   ,  �n���  �n  �  �  �  ����  �n���      C   ,  �����  ��  �  �F  �  �F���  �����      C   ,  �����  ��  �  ��  �  �����  �����      C   ,  �8���  �8  �  ��  �  �����  �8���      C   ,  �����  ��  �  �0  �  �0���  �����      C   ,  �����  ��  �  �~  �  �~���  �����      C   ,  �"���  �"  �  ��  �  �����  �"���      C   ,  ��  	�  ��  
�  �+  
�  �+  	�  ��  	�      C   ,  �/  	�  �/  
�  �y  
�  �y  	�  �/  	�      C   ,  �}  	�  �}  
�  ��  
�  ��  	�  �}  	�      C   ,  ��  	�  ��  
�  �  
�  �  	�  ��  	�      C   ,  �  	�  �  
�  �c  
�  �c  	�  �  	�      C   ,  �g  	�  �g  
�  ��  
�  ��  	�  �g  	�      C   ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C   ,  �  	�  �  
�  �M  
�  �M  	�  �  	�      C   ,  �Q  	�  �Q  
�  ��  
�  ��  	�  �Q  	�      C   ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C   ,  ��  	�  ��  
�  �7  
�  �7  	�  ��  	�      C   ,  �;  	�  �;  
�  ��  
�  ��  	�  �;  	�      C   ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C   ,  ��  	�  ��  
�  �!  
�  �!  	�  ��  	�      C   ,  �%  	�  �%  
�  �o  
�  �o  	�  �%  	�      C   ,  �s  	�  �s  
�  ��  
�  ��  	�  �s  	�      C   ,  ��  	�  ��  
�  �  
�  �  	�  ��  	�      C   ,  �  	�  �  
�  �Y  
�  �Y  	�  �  	�      C   ,  �]  	�  �]  
�  ��  
�  ��  	�  �]  	�      C   ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C   ,  �
���  �
  �  ��  �  �����  �
���      C   ,  ��  �  ��    �+    �+  �  ��  �      C   ,  �/  �  �/    �y    �y  �  �/  �      C   ,  �}  �  �}    ��    ��  �  �}  �      C   ,  ��  �  ��    �    �  �  ��  �      C   ,  �  �  �    �c    �c  �  �  �      C   ,  �g  �  �g    ��    ��  �  �g  �      C   ,  ��  �  ��    ��    ��  �  ��  �      C   ,  �  �  �    �M    �M  �  �  �      C   ,  �Q  �  �Q    ��    ��  �  �Q  �      C   ,  ��  �  ��    ��    ��  �  ��  �      C   ,  ��  �  ��    �7    �7  �  ��  �      C   ,  �;  �  �;    ��    ��  �  �;  �      C   ,  ��  �  ��    ��    ��  �  ��  �      C   ,  ��  �  ��    �!    �!  �  ��  �      C   ,  �%  �  �%    �o    �o  �  �%  �      C   ,  �s  �  �s    ��    ��  �  �s  �      C   ,  ��  �  ��    �    �  �  ��  �      C   ,  �  �  �    �Y    �Y  �  �  �      C   ,  �]  �  �]    ��    ��  �  �]  �      C   ,  ��  �  ��    ��    ��  �  ��  �      C   ,  �X���  �X  �  �  �  ����  �X���      C   ,  �����  ��  �  �P  �  �P���  �����      C   ,  �����  ��  �  ��  �  �����  �����      C   ,  �B���  �B  �  ��  �  �����  �B���      C   ,  �����  ��  �  �:  �  �:���  �����      C   ,  �����  ��  �  ��  �  �����  �����      C   ,  �,���  �,  �  ��  �  �����  �,���      C   ,  �z���  �z  �  �$  �  �$���  �z���      C   ,  �����  ��  �  �r  �  �r���  �����      C   ,  ����  �  �  ��  �  �����  ����      C   ,  �d���  �d  �  �  �  ����  �d���      C   ,  �����  ��  �  �\  �  �\���  �����      C   ,  � ���  �   �  ��  �  �����  � ���      C   ,  �
  r  �
  R  ��  R  ��  r  �
  r      C   ,  �X  r  �X  R  �  R  �  r  �X  r      C   ,  ��  r  ��  R  �P  R  �P  r  ��  r      C   ,  ��  r  ��  R  ��  R  ��  r  ��  r      C   ,  �B  r  �B  R  ��  R  ��  r  �B  r      C   ,  ��  r  ��  R  �:  R  �:  r  ��  r      C   ,  ��  r  ��  R  ��  R  ��  r  ��  r      C   ,  �,  r  �,  R  ��  R  ��  r  �,  r      C   ,  �z  r  �z  R  �$  R  �$  r  �z  r      C   ,  ��  r  ��  R  �r  R  �r  r  ��  r      C   ,  �  r  �  R  ��  R  ��  r  �  r      C   ,  �d  r  �d  R  �  R  �  r  �d  r      C   ,  ��  r  ��  R  �\  R  �\  r  ��  r      C   ,  �   r  �   R  ��  R  ��  r  �   r      C   ,  �N  r  �N  R  ��  R  ��  r  �N  r      C   ,  ��  r  ��  R  �F  R  �F  r  ��  r      C   ,  ��  r  ��  R  ��  R  ��  r  ��  r      C   ,  �8  r  �8  R  ��  R  ��  r  �8  r      C   ,  ��  r  ��  R  �0  R  �0  r  ��  r      C   ,  ��  r  ��  R  �~  R  �~  r  ��  r      C   ,  �"  r  �"  R  ��  R  ��  r  �"  r      C   ,  �N���  �N  �  ��  �  �����  �N���      C   ,  ������  �����  �����  ������  ������      C   ,  [����?  [����  \b���  \b���?  [����?      C   ,  ������  �����u  �����u  ������  ������      C   ,  ]����  ]�����  ^�����  ^����  ]����      C   ,  `@���  `@����  `�����  `����  `@���      C   ,  b����  b�����  c8����  c8���  b����      C   ,  d����  d�����  e�����  e����  d����      C   ,  g*���  g*����  g�����  g����  g*���      C   ,  ix���  ix����  j"����  j"���  ix���      C   ,  k����  k�����  lp����  lp���  k����      C   ,  n���  n����  n�����  n����  n���      C   ,  pb���  pb����  q����  q���  pb���      C   ,  r����  r�����  sZ����  sZ���  r����      C   ,  t����  t�����  u�����  u����  t����      C   ,  wL���  wL����  w�����  w����  wL���      C   ,  y����  y�����  zD����  zD���  y����      C   ,  {����  {�����  |�����  |����  {����      C   ,  ~6���  ~6����  ~�����  ~����  ~6���      C   ,  �����  ������  �.����  �.���  �����      C   ,  �����  ������  �|����  �|���  �����      C   ,  � ���  � ����  ������  �����  � ���      C   ,  �n���  �n����  �����  ����  �n���      C   ,  �����  ������  �f����  �f���  �����      C   ,  �
���  �
����  ������  �����  �
���      C   ,  �X���  �X����  �����  ����  �X���      C   ,  �����  ������  �P����  �P���  �����      C   ,  �����  ������  ������  �����  �����      C   ,  �B���  �B����  ������  �����  �B���      C   ,  �����  ������  �:����  �:���  �����      C   ,  �����  ������  ������  �����  �����      C   ,  �,���  �,����  ������  �����  �,���      C   ,  �z���  �z����  �$����  �$���  �z���      C   ,  �����  ������  �r����  �r���  �����      C   ,  ����  �����  ������  �����  ����      C   ,  �d���  �d����  �����  ����  �d���      C   ,  �����  ������  �\����  �\���  �����      C   ,  � ���  � ����  ������  �����  � ���      C   ,  �N���  �N����  ������  �����  �N���      C   ,  �����  ������  �F����  �F���  �����      C   ,  �����  ������  ������  �����  �����      C   ,  �8���  �8����  ������  �����  �8���      C   ,  �����  ������  �0����  �0���  �����      C   ,  �����  ������  �~����  �~���  �����      C   ,  �"���  �"����  ������  �����  �"���      C   ,  ������  �����  ����  �����  ������      C   ,  �����  ����  �c���  �c����  �����      C   ,  �g����  �g���  �����  ������  �g����      C   ,  ������  �����  �����  ������  ������      C   ,  �����  ����  �M���  �M����  �����      C   ,  �Q����  �Q���  �����  ������  �Q����      C   ,  ������  �����  �����  ������  ������      C   ,  ������  �����  �7���  �7����  ������      C   ,  �;����  �;���  �����  ������  �;����      C   ,  ������  �����  �����  ������  ������      C   ,  ������  �����  �!���  �!����  ������      C   ,  �%����  �%���  �o���  �o����  �%����      C   ,  �s����  �s���  �����  ������  �s����      C   ,  ������  �����  ����  �����  ������      C   ,  �����  ����  �Y���  �Y����  �����      C   ,  �]����  �]���  �����  ������  �]����      C   ,  ������  �����  �����  ������  ������      C   ,  ������  �����  �+���  �+����  ������      C   ,  �/����  �/���  �y���  �y����  �/����      C   ,  ������  �����u  �+���u  �+����  ������      C   ,  �/����  �/���u  �y���u  �y����  �/����      C   ,  �}����  �}���u  �����u  ������  �}����      C   ,  ������  �����u  ����u  �����  ������      C   ,  �����  ����u  �c���u  �c����  �����      C   ,  �g����  �g���u  �����u  ������  �g����      C   ,  ������  �����u  �����u  ������  ������      C   ,  �����  ����u  �M���u  �M����  �����      C   ,  �Q����  �Q���u  �����u  ������  �Q����      C   ,  ������  �����u  �����u  ������  ������      C   ,  ������  �����u  �7���u  �7����  ������      C   ,  �;����  �;���u  �����u  ������  �;����      C   ,  ������  �����u  �����u  ������  ������      C   ,  ������  �����u  �!���u  �!����  ������      C   ,  �%����  �%���u  �o���u  �o����  �%����      C   ,  �s����  �s���u  �����u  ������  �s����      C   ,  ������  �����u  ����u  �����  ������      C   ,  �����  ����u  �Y���u  �Y����  �����      C   ,  �]����  �]���u  �����u  ������  �]����      C   ,  ������  �����u  �����u  ������  ������      C   ,  �}����  �}���  �����  ������  �}����      C   ,  �
���h  �
���H  �����H  �����h  �
���h      C   ,  �X���h  �X���H  ����H  ����h  �X���h      C   ,  �����h  �����H  �P���H  �P���h  �����h      C   ,  �����h  �����H  �����H  �����h  �����h      C   ,  �B���h  �B���H  �����H  �����h  �B���h      C   ,  �����h  �����H  �:���H  �:���h  �����h      C   ,  �����h  �����H  �����H  �����h  �����h      C   ,  �,���h  �,���H  �����H  �����h  �,���h      C   ,  �z���h  �z���H  �$���H  �$���h  �z���h      C   ,  �����h  �����H  �r���H  �r���h  �����h      C   ,  ����h  ����H  �����H  �����h  ����h      C   ,  �d���h  �d���H  ����H  ����h  �d���h      C   ,  �����h  �����H  �\���H  �\���h  �����h      C   ,  � ���h  � ���H  �����H  �����h  � ���h      C   ,  �N���h  �N���H  �����H  �����h  �N���h      C   ,  �����h  �����H  �F���H  �F���h  �����h      C   ,  �����h  �����H  �����H  �����h  �����h      C   ,  �8���h  �8���H  �����H  �����h  �8���h      C   ,  �����h  �����H  �0���H  �0���h  �����h      C   ,  �����h  �����H  �~���H  �~���h  �����h      C   ,  �"���h  �"���H  �����H  �����h  �"���h      C   ,  b����h  b����H  c8���H  c8���h  b����h      C   ,  d����h  d����H  e����H  e����h  d����h      C   ,  g*���h  g*���H  g����H  g����h  g*���h      C   ,  ix���h  ix���H  j"���H  j"���h  ix���h      C   ,  k����h  k����H  lp���H  lp���h  k����h      C   ,  n���h  n���H  n����H  n����h  n���h      C   ,  pb���h  pb���H  q���H  q���h  pb���h      C   ,  r����h  r����H  sZ���H  sZ���h  r����h      C   ,  t����h  t����H  u����H  u����h  t����h      C   ,  wL���h  wL���H  w����H  w����h  wL���h      C   ,  y����h  y����H  zD���H  zD���h  y����h      C   ,  {����h  {����H  |����H  |����h  {����h      C   ,  ~6���h  ~6���H  ~����H  ~����h  ~6���h      C   ,  �����h  �����H  �.���H  �.���h  �����h      C   ,  �����h  �����H  �|���H  �|���h  �����h      C   ,  � ���h  � ���H  �����H  �����h  � ���h      C   ,  �n���h  �n���H  ����H  ����h  �n���h      C   ,  �����h  �����H  �f���H  �f���h  �����h      C   ,  e�����  e����u  f����u  f�����  e�����      C   ,  h����  h���u  iK���u  iK����  h����      C   ,  jO����  jO���u  k����u  k�����  jO����      C   ,  l�����  l����u  m����u  m�����  l�����      C   ,  n�����  n����u  p5���u  p5����  n�����      C   ,  q9����  q9���u  r����u  r�����  q9����      C   ,  s�����  s����u  t����u  t�����  s�����      C   ,  u�����  u����u  w���u  w����  u�����      C   ,  x#����  x#���u  ym���u  ym����  x#����      C   ,  zq����  zq���u  {����u  {�����  zq����      C   ,  |�����  |����u  ~	���u  ~	����  |�����      C   ,  ����  ���u  �W���u  �W����  ����      C   ,  �[����  �[���u  �����u  ������  �[����      C   ,  ������  �����u  �����u  ������  ������      C   ,  ������  �����u  �A���u  �A����  ������      C   ,  �E����  �E���u  �����u  ������  �E����      C   ,  ^�����  ^����u  `���u  `����  ^�����      C   ,  a����  a���u  ba���u  ba����  a����      C   ,  ]����h  ]����H  ^����H  ^����h  ]����h      C   ,  ce����  ce���u  d����u  d�����  ce����      C   ,  `@���h  `@���H  `����H  `����h  `@���h      C   ,  ^�����  ^����  `���  `����  ^�����      C   ,  a����  a���  ba���  ba����  a����      C   ,  ce����  ce���  d����  d�����  ce����      C   ,  e�����  e����  f����  f�����  e�����      C   ,  h����  h���  iK���  iK����  h����      C   ,  jO����  jO���  k����  k�����  jO����      C   ,  l�����  l����  m����  m�����  l�����      C   ,  n�����  n����  p5���  p5����  n�����      C   ,  q9����  q9���  r����  r�����  q9����      C   ,  s�����  s����  t����  t�����  s�����      C   ,  u�����  u����  w���  w����  u�����      C   ,  x#����  x#���  ym���  ym����  x#����      C   ,  zq����  zq���  {����  {�����  zq����      C   ,  |�����  |����  ~	���  ~	����  |�����      C   ,  ����  ���  �W���  �W����  ����      C   ,  �[����  �[���  �����  ������  �[����      C   ,  ������  �����  �����  ������  ������      C   ,  ������  �����  �A���  �A����  ������      C   ,  �E����  �E���  �����  ������  �E����      C   ,  �.���h  �.���H  �����H  �����h  �.���h      C   ,  �p���h  �p���H  ����H  ����h  �p���h      C   ,  �G����  �G���  �����  ������  �G����      C   ,  ������  �����  �����  ������  ������      C   ,  ������  �����  �-���  �-����  ������      C   ,  �1����  �1���  �{���  �{����  �1����      C   ,  �����  ����  �����  ������  �����      C   ,  ������  �����  ����  �����  ������      C   ,  �p���  �p����  �����  ����  �p���      C   ,  �����  ������  �h����  �h���  �����      C   ,  ����  �����  ������  �����  ����      C   ,  �Z���  �Z����  �����  ����  �Z���      C   ,  Ũ���  Ũ����  �R����  �R���  Ũ���      C   ,  �����  ������  Ƞ����  Ƞ���  �����      C   ,  �D���  �D����  ������  �����  �D���      C   ,  ̒���  ̒����  �<����  �<���  ̒���      C   ,  �����  ������  ϊ����  ϊ���  �����      C   ,  �.���  �.����  ������  �����  �.���      C   ,  �h���?  �h���  ����  ����?  �h���?      C   ,  �����  ����  �e���  �e����  �����      C   ,  �i����  �i���  γ���  γ����  �i����      C   ,  Ϸ����  Ϸ���  ����  �����  Ϸ����      C   ,  �����h  �����H  �h���H  �h���h  �����h      C   ,  ����h  ����H  �����H  �����h  ����h      C   ,  �Z���h  �Z���H  ����H  ����h  �Z���h      C   ,  �G����  �G���u  �����u  ������  �G����      C   ,  ������  �����u  �����u  ������  ������      C   ,  ������  �����u  �-���u  �-����  ������      C   ,  �1����  �1���u  �{���u  �{����  �1����      C   ,  �����  ����u  �����u  ������  �����      C   ,  ������  �����u  ����u  �����  ������      C   ,  �����  ����u  �e���u  �e����  �����      C   ,  �i����  �i���u  γ���u  γ����  �i����      C   ,  Ϸ����  Ϸ���u  ����u  �����  Ϸ����      C   ,  Ũ���h  Ũ���H  �R���H  �R���h  Ũ���h      C   ,  �����h  �����H  Ƞ���H  Ƞ���h  �����h      C   ,  �D���h  �D���H  �����H  �����h  �D���h      C   ,  ̒���h  ̒���H  �<���H  �<���h  ̒���h      C   ,  �����h  �����H  ϊ���H  ϊ���h  �����h      C   ,  ������  ������  �C����  �C����  ������      C   ,  ������  �����k  �C���k  �C����  ������      C   ,  [�����  [����5  ����5  �����  [�����      C   ,  \�����  \����}  ����}  �����  \�����      C   ,  \����  \�����  �����  ����  \����      C   ,  ������  �����}  �C���}  �C����  ������      C   ,  ������  �����a  �C���a  �C����  ������      C   ,  ]����P  ]�����  ^�����  ^����P  ]����P      C   ,  `@���P  `@����  `�����  `����P  `@���P      C   ,  b����P  b�����  c8����  c8���P  b����P      C   ,  d����P  d�����  e�����  e����P  d����P      C   ,  g*���P  g*����  g�����  g����P  g*���P      C   ,  ix���P  ix����  j"����  j"���P  ix���P      C   ,  k����P  k�����  lp����  lp���P  k����P      C   ,  n���P  n����  n�����  n����P  n���P      C   ,  pb���P  pb����  q����  q���P  pb���P      C   ,  r����P  r�����  sZ����  sZ���P  r����P      C   ,  t����P  t�����  u�����  u����P  t����P      C   ,  wL���P  wL����  w�����  w����P  wL���P      C   ,  y����P  y�����  zD����  zD���P  y����P      C   ,  {����P  {�����  |�����  |����P  {����P      C   ,  ~6���P  ~6����  ~�����  ~����P  ~6���P      C   ,  �����P  ������  �.����  �.���P  �����P      C   ,  �����P  ������  �|����  �|���P  �����P      C   ,  � ���P  � ����  ������  �����P  � ���P      C   ,  �n���P  �n����  �����  ����P  �n���P      C   ,  �����P  ������  �f����  �f���P  �����P      C   ,  �
���P  �
����  ������  �����P  �
���P      C   ,  �X���P  �X����  �����  ����P  �X���P      C   ,  �����P  ������  �P����  �P���P  �����P      C   ,  �����P  ������  ������  �����P  �����P      C   ,  �B���P  �B����  ������  �����P  �B���P      C   ,  �����P  ������  �:����  �:���P  �����P      C   ,  �����P  ������  ������  �����P  �����P      C   ,  �,���P  �,����  ������  �����P  �,���P      C   ,  �z���P  �z����  �$����  �$���P  �z���P      C   ,  �����P  ������  �r����  �r���P  �����P      C   ,  ����P  �����  ������  �����P  ����P      C   ,  �d���P  �d����  �����  ����P  �d���P      C   ,  �����P  ������  �\����  �\���P  �����P      C   ,  � ���P  � ����  ������  �����P  � ���P      C   ,  �N���P  �N����  ������  �����P  �N���P      C   ,  �����P  ������  �F����  �F���P  �����P      C   ,  �����P  ������  ������  �����P  �����P      C   ,  �8���P  �8����  ������  �����P  �8���P      C   ,  �����P  ������  �0����  �0���P  �����P      C   ,  �����P  ������  �~����  �~���P  �����P      C   ,  �"���P  �"����  ������  �����P  �"���P      C   ,  �p���P  �p����  �����  ����P  �p���P      C   ,  �����P  ������  �h����  �h���P  �����P      C   ,  ����P  �����  ������  �����P  ����P      C   ,  �Z���P  �Z����  �����  ����P  �Z���P      C   ,  Ũ���P  Ũ����  �R����  �R���P  Ũ���P      C   ,  �����P  ������  Ƞ����  Ƞ���P  �����P      C   ,  �D���P  �D����  ������  �����P  �D���P      C   ,  ̒���P  ̒����  �<����  �<���P  ̒���P      C   ,  �����P  ������  ϊ����  ϊ���P  �����P      C   ,  �.���P  �.����  ������  �����P  �.���P      C   ,  ]H��}�  ]H��~s  ҂��~s  ҂��}�  ]H��}�      C   ,  ]H��|  ]H��|�  ҂��|�  ҂��|  ]H��|      C   ,  ����f1  ����f�  �/��f�  �/��f1  ����f1      C   ,  ����d  ����d�  �/��d�  �/��d  ����d      C   ,  Ϸ����  Ϸ���a  ����a  �����  Ϸ����      C   ,  �����  �����  �e����  �e����  �����      C   ,  �i����  �i����  γ����  γ����  �i����      C   ,  Ϸ����  Ϸ����  �����  �����  Ϸ����      C   ,  �G����  �G����  ������  ������  �G����      C   ,  �G����  �G���k  �����k  ������  �G����      C   ,  ������  �����k  �����k  ������  ������      C   ,  ������  �����k  �-���k  �-����  ������      C   ,  �1����  �1���k  �{���k  �{����  �1����      C   ,  �����  ����k  �����k  ������  �����      C   ,  ������  �����k  ����k  �����  ������      C   ,  �����  ����k  �e���k  �e����  �����      C   ,  �i����  �i���k  γ���k  γ����  �i����      C   ,  Ϸ����  Ϸ���k  ����k  �����  Ϸ����      C   ,  �p���
  �p����  �����  ����
  �p���
      C   ,  �����
  ������  �h����  �h���
  �����
      C   ,  ����
  �����  ������  �����
  ����
      C   ,  �Z���
  �Z����  �����  ����
  �Z���
      C   ,  Ũ���
  Ũ����  �R����  �R���
  Ũ���
      C   ,  �����
  ������  Ƞ����  Ƞ���
  �����
      C   ,  �D���
  �D����  ������  �����
  �D���
      C   ,  ̒���
  ̒����  �<����  �<���
  ̒���
      C   ,  �����
  ������  ϊ����  ϊ���
  �����
      C   ,  �.���
  �.����  ������  �����
  �.���
      C   ,  ������  ������  ������  ������  ������      C   ,  ������  ������  �-����  �-����  ������      C   ,  �1����  �1����  �{����  �{����  �1����      C   ,  �p����  �p����  �����  �����  �p����      C   ,  ������  ������  �h����  �h����  ������      C   ,  �����  �����  ������  ������  �����      C   ,  �Z����  �Z����  �����  �����  �Z����      C   ,  Ũ����  Ũ����  �R����  �R����  Ũ����      C   ,  ������  ������  Ƞ����  Ƞ����  ������      C   ,  �D����  �D����  ������  ������  �D����      C   ,  ̒����  ̒����  �<����  �<����  ̒����      C   ,  ������  ������  ϊ����  ϊ����  ������      C   ,  �.����  �.����  ������  ������  �.����      C   ,  �����  �����  ������  ������  �����      C   ,  �G����  �G���}  �����}  ������  �G����      C   ,  ������  �����}  �����}  ������  ������      C   ,  ������  �����}  �-���}  �-����  ������      C   ,  �1����  �1���}  �{���}  �{����  �1����      C   ,  �����  ����}  �����}  ������  �����      C   ,  ������  �����}  ����}  �����  ������      C   ,  �����  ����}  �e���}  �e����  �����      C   ,  �i����  �i���}  γ���}  γ����  �i����      C   ,  Ϸ����  Ϸ���}  ����}  �����  Ϸ����      C   ,  ������  ������  �����  �����  ������      C   ,  �G����  �G���a  �����a  ������  �G����      C   ,  ������  �����a  �����a  ������  ������      C   ,  ������  �����a  �-���a  �-����  ������      C   ,  �1����  �1���a  �{���a  �{����  �1����      C   ,  �����  ����a  �����a  ������  �����      C   ,  ������  �����a  ����a  �����  ������      C   ,  �����  ����a  �e���a  �e����  �����      C   ,  �i����  �i���a  γ���a  γ����  �i����      C   ,  ������  �����}  �����}  ������  ������      C   ,  ������  �����a  �����a  ������  ������      C   ,  ������  �����k  �����k  ������  ������      C   ,  ������  ������  ������  ������  ������      C   ,  �����
  ������  �:����  �:���
  �����
      C   ,  �����
  ������  ������  �����
  �����
      C   ,  �,���
  �,����  ������  �����
  �,���
      C   ,  �z���
  �z����  �$����  �$���
  �z���
      C   ,  �����
  ������  �r����  �r���
  �����
      C   ,  ����
  �����  ������  �����
  ����
      C   ,  �d���
  �d����  �����  ����
  �d���
      C   ,  �����
  ������  �\����  �\���
  �����
      C   ,  � ���
  � ����  ������  �����
  � ���
      C   ,  �N���
  �N����  ������  �����
  �N���
      C   ,  �����
  ������  �F����  �F���
  �����
      C   ,  �����
  ������  ������  �����
  �����
      C   ,  �8���
  �8����  ������  �����
  �8���
      C   ,  �����
  ������  �0����  �0���
  �����
      C   ,  �����
  ������  �~����  �~���
  �����
      C   ,  �"���
  �"����  ������  �����
  �"���
      C   ,  ������  ������  �����  �����  ������      C   ,  �����  �����  �c����  �c����  �����      C   ,  �g����  �g����  ������  ������  �g����      C   ,  ������  ������  ������  ������  ������      C   ,  �����  �����  �M����  �M����  �����      C   ,  �Q����  �Q����  ������  ������  �Q����      C   ,  ������  ������  ������  ������  ������      C   ,  ������  ������  �7����  �7����  ������      C   ,  �;����  �;����  ������  ������  �;����      C   ,  ������  ������  ������  ������  ������      C   ,  ������  ������  �!����  �!����  ������      C   ,  �%����  �%����  �o����  �o����  �%����      C   ,  �s����  �s����  ������  ������  �s����      C   ,  ������  ������  �����  �����  ������      C   ,  �����  �����  �Y����  �Y����  �����      C   ,  �]����  �]����  ������  ������  �]����      C   ,  ������  ������  ������  ������  ������      C   ,  �X���
  �X����  �����  ����
  �X���
      C   ,  �����
  ������  �P����  �P���
  �����
      C   ,  �����
  ������  ������  �����
  �����
      C   ,  ������  �����k  �+���k  �+����  ������      C   ,  �/����  �/���k  �y���k  �y����  �/����      C   ,  �}����  �}���k  �����k  ������  �}����      C   ,  ������  �����k  ����k  �����  ������      C   ,  �����  ����k  �c���k  �c����  �����      C   ,  �g����  �g���k  �����k  ������  �g����      C   ,  ������  �����k  �����k  ������  ������      C   ,  �����  ����k  �M���k  �M����  �����      C   ,  �Q����  �Q���k  �����k  ������  �Q����      C   ,  ������  �����k  �����k  ������  ������      C   ,  ������  �����k  �7���k  �7����  ������      C   ,  �;����  �;���k  �����k  ������  �;����      C   ,  ������  �����k  �����k  ������  ������      C   ,  ������  �����k  �!���k  �!����  ������      C   ,  �%����  �%���k  �o���k  �o����  �%����      C   ,  �s����  �s���k  �����k  ������  �s����      C   ,  ������  �����k  ����k  �����  ������      C   ,  �����  ����k  �Y���k  �Y����  �����      C   ,  �]����  �]���k  �����k  ������  �]����      C   ,  ������  �����k  �����k  ������  ������      C   ,  �B���
  �B����  ������  �����
  �B���
      C   ,  ������  ������  �+����  �+����  ������      C   ,  �/����  �/����  �y����  �y����  �/����      C   ,  �}����  �}����  ������  ������  �}����      C   ,  �
���
  �
����  ������  �����
  �
���
      C   ,  �[����  �[���k  �����k  ������  �[����      C   ,  ������  �����k  �����k  ������  ������      C   ,  ������  �����k  �A���k  �A����  ������      C   ,  �E����  �E���k  �����k  ������  �E����      C   ,  h����  h����  iK����  iK����  h����      C   ,  jO����  jO����  k�����  k�����  jO����      C   ,  l�����  l�����  m�����  m�����  l�����      C   ,  n�����  n�����  p5����  p5����  n�����      C   ,  q9����  q9����  r�����  r�����  q9����      C   ,  ^�����  ^�����  `����  `����  ^�����      C   ,  s�����  s�����  t�����  t�����  s�����      C   ,  u�����  u�����  w����  w����  u�����      C   ,  x#����  x#����  ym����  ym����  x#����      C   ,  zq����  zq����  {�����  {�����  zq����      C   ,  ^�����  ^����k  `���k  `����  ^�����      C   ,  a����  a���k  ba���k  ba����  a����      C   ,  ce����  ce���k  d����k  d�����  ce����      C   ,  e�����  e����k  f����k  f�����  e�����      C   ,  h����  h���k  iK���k  iK����  h����      C   ,  jO����  jO���k  k����k  k�����  jO����      C   ,  e�����  e�����  f�����  f�����  e�����      C   ,  l�����  l����k  m����k  m�����  l�����      C   ,  n�����  n����k  p5���k  p5����  n�����      C   ,  q9����  q9���k  r����k  r�����  q9����      C   ,  s�����  s����k  t����k  t�����  s�����      C   ,  |�����  |�����  ~	����  ~	����  |�����      C   ,  ����  ����  �W����  �W����  ����      C   ,  �[����  �[����  ������  ������  �[����      C   ,  ������  ������  ������  ������  ������      C   ,  ������  ������  �A����  �A����  ������      C   ,  �E����  �E����  ������  ������  �E����      C   ,  u�����  u����k  w���k  w����  u�����      C   ,  x#����  x#���k  ym���k  ym����  x#����      C   ,  zq����  zq���k  {����k  {�����  zq����      C   ,  |�����  |����k  ~	���k  ~	����  |�����      C   ,  ]����
  ]�����  ^�����  ^����
  ]����
      C   ,  `@���
  `@����  `�����  `����
  `@���
      C   ,  b����
  b�����  c8����  c8���
  b����
      C   ,  d����
  d�����  e�����  e����
  d����
      C   ,  g*���
  g*����  g�����  g����
  g*���
      C   ,  ix���
  ix����  j"����  j"���
  ix���
      C   ,  k����
  k�����  lp����  lp���
  k����
      C   ,  n���
  n����  n�����  n����
  n���
      C   ,  pb���
  pb����  q����  q���
  pb���
      C   ,  r����
  r�����  sZ����  sZ���
  r����
      C   ,  t����
  t�����  u�����  u����
  t����
      C   ,  wL���
  wL����  w�����  w����
  wL���
      C   ,  y����
  y�����  zD����  zD���
  y����
      C   ,  {����
  {�����  |�����  |����
  {����
      C   ,  ~6���
  ~6����  ~�����  ~����
  ~6���
      C   ,  �����
  ������  �.����  �.���
  �����
      C   ,  �����
  ������  �|����  �|���
  �����
      C   ,  � ���
  � ����  ������  �����
  � ���
      C   ,  �n���
  �n����  �����  ����
  �n���
      C   ,  �����
  ������  �f����  �f���
  �����
      C   ,  ����  ���k  �W���k  �W����  ����      C   ,  a����  a����  ba����  ba����  a����      C   ,  ce����  ce����  d�����  d�����  ce����      C   ,  jO����  jO���}  k����}  k�����  jO����      C   ,  l�����  l����}  m����}  m�����  l�����      C   ,  n�����  n����}  p5���}  p5����  n�����      C   ,  q9����  q9���}  r����}  r�����  q9����      C   ,  s�����  s����}  t����}  t�����  s�����      C   ,  u�����  u����}  w���}  w����  u�����      C   ,  x#����  x#���}  ym���}  ym����  x#����      C   ,  zq����  zq���}  {����}  {�����  zq����      C   ,  |�����  |����}  ~	���}  ~	����  |�����      C   ,  ����  ���}  �W���}  �W����  ����      C   ,  �[����  �[���}  �����}  ������  �[����      C   ,  ������  �����}  �����}  ������  ������      C   ,  ������  �����}  �A���}  �A����  ������      C   ,  �E����  �E���}  �����}  ������  �E����      C   ,  y�����  y�����  zD����  zD����  y�����      C   ,  {�����  {�����  |�����  |�����  {�����      C   ,  ~6����  ~6����  ~�����  ~�����  ~6����      C   ,  ������  ������  �.����  �.����  ������      C   ,  ������  ������  �|����  �|����  ������      C   ,  � ����  � ����  ������  ������  � ����      C   ,  �n����  �n����  �����  �����  �n����      C   ,  ������  ������  �f����  �f����  ������      C   ,  b�����  b�����  c8����  c8����  b�����      C   ,  d�����  d�����  e�����  e�����  d�����      C   ,  g*����  g*����  g�����  g�����  g*����      C   ,  ^�����  ^����a  `���a  `����  ^�����      C   ,  a����  a���a  ba���a  ba����  a����      C   ,  ce����  ce���a  d����a  d�����  ce����      C   ,  e�����  e����a  f����a  f�����  e�����      C   ,  h����  h���a  iK���a  iK����  h����      C   ,  jO����  jO���a  k����a  k�����  jO����      C   ,  l�����  l����a  m����a  m�����  l�����      C   ,  n�����  n����a  p5���a  p5����  n�����      C   ,  q9����  q9���a  r����a  r�����  q9����      C   ,  s�����  s����a  t����a  t�����  s�����      C   ,  u�����  u����a  w���a  w����  u�����      C   ,  x#����  x#���a  ym���a  ym����  x#����      C   ,  zq����  zq���a  {����a  {�����  zq����      C   ,  |�����  |����a  ~	���a  ~	����  |�����      C   ,  ����  ���a  �W���a  �W����  ����      C   ,  �[����  �[���a  �����a  ������  �[����      C   ,  ������  �����a  �����a  ������  ������      C   ,  ������  �����a  �A���a  �A����  ������      C   ,  �E����  �E���a  �����a  ������  �E����      C   ,  ix����  ix����  j"����  j"����  ix����      C   ,  k�����  k�����  lp����  lp����  k�����      C   ,  n����  n����  n�����  n�����  n����      C   ,  pb����  pb����  q����  q����  pb����      C   ,  r�����  r�����  sZ����  sZ����  r�����      C   ,  t�����  t�����  u�����  u�����  t�����      C   ,  wL����  wL����  w�����  w�����  wL����      C   ,  ^�����  ^����}  `���}  `����  ^�����      C   ,  a����  a���}  ba���}  ba����  a����      C   ,  ce����  ce���}  d����}  d�����  ce����      C   ,  e�����  e����}  f����}  f�����  e�����      C   ,  h����  h���}  iK���}  iK����  h����      C   ,  �s����  �s���}  �����}  ������  �s����      C   ,  ������  �����}  ����}  �����  ������      C   ,  �����  ����}  �Y���}  �Y����  �����      C   ,  �]����  �]���}  �����}  ������  �]����      C   ,  ������  �����}  �����}  ������  ������      C   ,  ������  ������  �r����  �r����  ������      C   ,  �����  �����  ������  ������  �����      C   ,  �d����  �d����  �����  �����  �d����      C   ,  ������  ������  �\����  �\����  ������      C   ,  � ����  � ����  ������  ������  � ����      C   ,  �N����  �N����  ������  ������  �N����      C   ,  ������  ������  �F����  �F����  ������      C   ,  ������  ������  ������  ������  ������      C   ,  �8����  �8����  ������  ������  �8����      C   ,  ������  ������  �0����  �0����  ������      C   ,  ������  ������  �~����  �~����  ������      C   ,  �"����  �"����  ������  ������  �"����      C   ,  �
����  �
����  ������  ������  �
����      C   ,  �X����  �X����  �����  �����  �X����      C   ,  ������  ������  �P����  �P����  ������      C   ,  ������  ������  ������  ������  ������      C   ,  �B����  �B����  ������  ������  �B����      C   ,  ������  ������  �:����  �:����  ������      C   ,  ������  ������  ������  ������  ������      C   ,  �,����  �,����  ������  ������  �,����      C   ,  �z����  �z����  �$����  �$����  �z����      C   ,  ������  �����}  �+���}  �+����  ������      C   ,  �/����  �/���}  �y���}  �y����  �/����      C   ,  �}����  �}���}  �����}  ������  �}����      C   ,  ������  �����}  ����}  �����  ������      C   ,  �����  ����}  �c���}  �c����  �����      C   ,  �g����  �g���}  �����}  ������  �g����      C   ,  ������  �����}  �����}  ������  ������      C   ,  �����  ����}  �M���}  �M����  �����      C   ,  �Q����  �Q���}  �����}  ������  �Q����      C   ,  ������  �����a  �+���a  �+����  ������      C   ,  �/����  �/���a  �y���a  �y����  �/����      C   ,  �}����  �}���a  �����a  ������  �}����      C   ,  ������  �����a  ����a  �����  ������      C   ,  �����  ����a  �c���a  �c����  �����      C   ,  �g����  �g���a  �����a  ������  �g����      C   ,  ������  �����a  �����a  ������  ������      C   ,  �����  ����a  �M���a  �M����  �����      C   ,  �Q����  �Q���a  �����a  ������  �Q����      C   ,  ������  �����a  �����a  ������  ������      C   ,  ������  �����a  �7���a  �7����  ������      C   ,  �;����  �;���a  �����a  ������  �;����      C   ,  ������  �����a  �����a  ������  ������      C   ,  ������  �����a  �!���a  �!����  ������      C   ,  �%����  �%���a  �o���a  �o����  �%����      C   ,  �s����  �s���a  �����a  ������  �s����      C   ,  ������  �����a  ����a  �����  ������      C   ,  �����  ����a  �Y���a  �Y����  �����      C   ,  �]����  �]���a  �����a  ������  �]����      C   ,  ������  �����a  �����a  ������  ������      C   ,  ������  �����}  �����}  ������  ������      C   ,  ������  �����}  �7���}  �7����  ������      C   ,  �;����  �;���}  �����}  ������  �;����      C   ,  ������  �����}  �����}  ������  ������      C   ,  ������  �����}  �!���}  �!����  ������      C   ,  �%����  �%���}  �o���}  �o����  �%����      C   ,  ����g�  ����s  �B��s  �B��g�  ����g�      C   ,  ����g�  ����s  ����s  ����g�  ����g�      C   ,  �4��g�  �4��s  ����s  ����g�  �4��g�      C   ,  ����g�  ����s  �,��s  �,��g�  ����g�      C   ,  ����g�  ����s  �z��s  �z��g�  ����g�      C   ,  ���g�  ���s  ����s  ����g�  ���g�      C   ,  �l��g�  �l��s  ���s  ���g�  �l��g�      C   ,  ����g�  ����s  �d��s  �d��g�  ����g�      C   ,  ���g�  ���s  ����s  ����g�  ���g�      C   ,  �V��g�  �V��s  � ��s  � ��g�  �V��g�      C   ,  ����g�  ����s  �t��s  �t��g�  ����g�      C   ,  ���g�  ���s  ����s  ����g�  ���g�      C   ,  �f��g�  �f��s  ���s  ���g�  �f��g�      C   ,  ����g�  ����s  �^��s  �^��g�  ����g�      C   ,  ���g�  ���s  ����s  ����g�  ���g�      C   ,  �P��g�  �P��s  ����s  ����g�  �P��g�      C   ,  ����g�  ����s  �H��s  �H��g�  ����g�      C   ,  ����g�  ����s  ����s  ����g�  ����g�      C   ,  �:��g�  �:��s  ����s  ����g�  �:��g�      C   ,  ����g�  ����s  �2��s  �2��g�  ����g�      C   ,  ����g�  ����s  ����s  ����g�  ����g�      C   ,  �$��g�  �$��s  ����s  ����g�  �$��g�      C   ,  �r��g�  �r��s  ���s  ���g�  �r��g�      C   ,  ����g�  ����s  �j��s  �j��g�  ����g�      C   ,  ���g�  ���s  ����s  ����g�  ���g�      C   ,  ����f1  ����f�  ����f�  ����f1  ����f1      C   ,  w`��g�  w`��s  x
��s  x
��g�  w`��g�      C   ,  ����d  ����d�  ����d�  ����d  ����d      C   ,  y���g�  y���s  zX��s  zX��g�  y���g�      C   ,  {���g�  {���s  |���s  |���g�  {���g�      C   ,  ~J��g�  ~J��s  ~���s  ~���g�  ~J��g�      C   ,  �o��f1  �o��f�  ����f�  ����f1  �o��f1      C   ,  ����f1  ����f�  ���f�  ���f1  ����f1      C   ,  ���f1  ���f�  �U��f�  �U��f1  ���f1      C   ,  �Y��f1  �Y��f�  ����f�  ����f1  �Y��f1      C   ,  s���f1  s���f�  t���f�  t���f1  s���f1      C   ,  u���f1  u���f�  w3��f�  w3��f1  u���f1      C   ,  s���d  s���d�  t���d�  t���d  s���d      C   ,  u���d  u���d�  w3��d�  w3��d  u���d      C   ,  x7��d  x7��d�  y���d�  y���d  x7��d      C   ,  z���d  z���d�  {���d�  {���d  z���d      C   ,  |���d  |���d�  ~��d�  ~��d  |���d      C   ,  !��d  !��d�  �k��d�  �k��d  !��d      C   ,  �o��d  �o��d�  ����d�  ����d  �o��d      C   ,  ����d  ����d�  ���d�  ���d  ����d      C   ,  ���d  ���d�  �U��d�  �U��d  ���d      C   ,  �Y��d  �Y��d�  ����d�  ����d  �Y��d      C   ,  x7��f1  x7��f�  y���f�  y���f1  x7��f1      C   ,  z���f1  z���f�  {���f�  {���f1  z���f1      C   ,  r���W�  r���c  sn��c  sn��W�  r���W�      C   ,  u��W�  u��c  u���c  u���W�  u��W�      C   ,  w`��W�  w`��c  x
��c  x
��W�  w`��W�      C   ,  y���W�  y���c  zX��c  zX��W�  y���W�      C   ,  {���W�  {���c  |���c  |���W�  {���W�      C   ,  ~J��W�  ~J��c  ~���c  ~���W�  ~J��W�      C   ,  ����W�  ����c  �B��c  �B��W�  ����W�      C   ,  ����W�  ����c  ����c  ����W�  ����W�      C   ,  �4��W�  �4��c  ����c  ����W�  �4��W�      C   ,  ����W�  ����c  �,��c  �,��W�  ����W�      C   ,  ����W�  ����c  �z��c  �z��W�  ����W�      C   ,  |���f1  |���f�  ~��f�  ~��f1  |���f1      C   ,  !��f1  !��f�  �k��f�  �k��f1  !��f1      C   ,  ����f1  ����f�  �#��f�  �#��f1  ����f1      C   ,  �'��f1  �'��f�  �q��f�  �q��f1  �'��f1      C   ,  �u��f1  �u��f�  ����f�  ����f1  �u��f1      C   ,  ����f1  ����f�  ���f�  ���f1  ����f1      C   ,  ����d  ����d�  �?��d�  �?��d  ����d      C   ,  �C��d  �C��d�  ����d�  ����d  �C��d      C   ,  ����d  ����d�  ����d�  ����d  ����d      C   ,  ����d  ����d�  �)��d�  �)��d  ����d      C   ,  ����d  ����d�  ����d�  ����d  ����d      C   ,  ����d  ����d�  �9��d�  �9��d  ����d      C   ,  �=��d  �=��d�  ����d�  ����d  �=��d      C   ,  ����d  ����d�  ����d�  ����d  ����d      C   ,  ����d  ����d�  �#��d�  �#��d  ����d      C   ,  �'��d  �'��d�  �q��d�  �q��d  �'��d      C   ,  �u��d  �u��d�  ����d�  ����d  �u��d      C   ,  ����d  ����d�  ���d�  ���d  ����d      C   ,  ���d  ���d�  �[��d�  �[��d  ���d      C   ,  �_��d  �_��d�  ����d�  ����d  �_��d      C   ,  ����d  ����d�  ����d�  ����d  ����d      C   ,  ����d  ����d�  �E��d�  �E��d  ����d      C   ,  �I��d  �I��d�  ����d�  ����d  �I��d      C   ,  ����d  ����d�  ����d�  ����d  ����d      C   ,  ���f1  ���f�  �[��f�  �[��f1  ���f1      C   ,  �_��f1  �_��f�  ����f�  ����f1  �_��f1      C   ,  ����f1  ����f�  ����f�  ����f1  ����f1      C   ,  ����f1  ����f�  �E��f�  �E��f1  ����f1      C   ,  �I��f1  �I��f�  ����f�  ����f1  �I��f1      C   ,  ����f1  ����f�  ����f�  ����f1  ����f1      C   ,  ����f1  ����f�  �?��f�  �?��f1  ����f1      C   ,  �C��f1  �C��f�  ����f�  ����f1  �C��f1      C   ,  ����f1  ����f�  ����f�  ����f1  ����f1      C   ,  ����f1  ����f�  �)��f�  �)��f1  ����f1      C   ,  ����f1  ����f�  ����f�  ����f1  ����f1      C   ,  ����f1  ����f�  �9��f�  �9��f1  ����f1      C   ,  ���W�  ���c  ����c  ����W�  ���W�      C   ,  �l��W�  �l��c  ���c  ���W�  �l��W�      C   ,  ����W�  ����c  �d��c  �d��W�  ����W�      C   ,  ���W�  ���c  ����c  ����W�  ���W�      C   ,  �V��W�  �V��c  � ��c  � ��W�  �V��W�      C   ,  ����W�  ����c  �t��c  �t��W�  ����W�      C   ,  ���W�  ���c  ����c  ����W�  ���W�      C   ,  �f��W�  �f��c  ���c  ���W�  �f��W�      C   ,  ����W�  ����c  �^��c  �^��W�  ����W�      C   ,  ���W�  ���c  ����c  ����W�  ���W�      C   ,  �P��W�  �P��c  ����c  ����W�  �P��W�      C   ,  ����W�  ����c  �H��c  �H��W�  ����W�      C   ,  ����W�  ����c  ����c  ����W�  ����W�      C   ,  �:��W�  �:��c  ����c  ����W�  �:��W�      C   ,  ����W�  ����c  �2��c  �2��W�  ����W�      C   ,  ����W�  ����c  ����c  ����W�  ����W�      C   ,  �$��W�  �$��c  ����c  ����W�  �$��W�      C   ,  �r��W�  �r��c  ���c  ���W�  �r��W�      C   ,  ����W�  ����c  �j��c  �j��W�  ����W�      C   ,  ���W�  ���c  ����c  ����W�  ���W�      C   ,  �=��f1  �=��f�  ����f�  ����f1  �=��f1      C   ,  ����f1  ����f�  ����f�  ����f1  ����f1      C   ,  �Z��f  �Z��f�  ���f�  ���f  �Z��f      C   ,  �Z��d�  �Z��eF  ���eF  ���d�  �Z��d�      C   ,  �Z��c*  �Z��c�  ���c�  ���c*  �Z��c*      C   ,  �Z��n�  �Z��od  ���od  ���n�  �Z��n�      C   ,  �Z��mH  �Z��m�  ���m�  ���mH  �Z��mH      C   ,  �Z��k�  �Z��l�  ���l�  ���k�  �Z��k�      C   ,  �Z��jd  �Z��k  ���k  ���jd  �Z��jd      C   ,  �Z��h�  �Z��i�  ���i�  ���h�  �Z��h�      C   ,  �Z��g�  �Z��h*  ���h*  ���g�  �Z��g�      C   ,  �\��g�  �\��s  ���s  ���g�  �\��g�      C   ,  �\��W�  �\��c  ���c  ���W�  �\��W�      C   ,  �Z��a�  �Z��bb  ���bb  ���a�  �Z��a�      C   ,  ����a�  ����s  �x��s  �x��a�  ����a�      C   ,  ����a�  ����s  �\��s  �\��a�  ����a�      C   ,  ����a�  ����s  �@��s  �@��a�  ����a�      C   ,  �z��a�  �z��s  �$��s  �$��a�  �z��a�      C   ,  ^��a�  ^��s ��s ��a�  ^��a�      C   , B��a� B��s ���s ���a� B��a�      C   , &��a� &��s ���s ���a� &��a�      C   , 	
��a� 	
��s 	���s 	���a� 	
��a�      C   , ���a� ���s ���s ���a� ���a�      C   , ���a� ���s |��s |��a� ���a�      C   , ���a� ���s `��s `��a� ���a�      C   , ���a� ���s D��s D��a� ���a�      C   , ~��a� ~��s (��s (��a� ~��a�      C   , b��a� b��s ��s ��a� b��a�      C   ,  �Z��q�  �Z��rH  ���rH  ���q�  �Z��q�      C   ,  �Z��`F  �Z��`�  ���`�  ���`F  �Z��`F      C   ,  ����`U  ����`�  �Z��`�  �Z��`U  ����`U      C   ,  �|��`U  �|��`�  �>��`�  �>��`U  �|��`U      C   ,  �`��`U  �`��`�  "��`�  "��`U  �`��`U      C   , D��`U D��`� ��`� ��`U D��`U      C   , (��`U (��`� ���`� ���`U (��`U      C   , ��`U ��`� ���`� ���`U ��`U      C   , 	���`U 	���`� ���`� ���`U 	���`U      C   , ���`U ���`� ���`� ���`U ���`U      C   , ���`U ���`� z��`� z��`U ���`U      C   , ���`U ���`� ^��`� ^��`U ���`U      C   , ���`U ���`� B��`� B��`U ���`U      C   , d��`U d��`� &��`� &��`U d��`U      C   , H��`U H��`� 
��`� 
��`U H��`U      C   ,  �Z��^�  �Z��_~  ���_~  ���^�  �Z��^�      C   ,  ����^9  ����^�  �Z��^�  �Z��^9  ����^9      C   ,  �|��^9  �|��^�  �>��^�  �>��^9  �|��^9      C   ,  �`��^9  �`��^�  "��^�  "��^9  �`��^9      C   , D��^9 D��^� ��^� ��^9 D��^9      C   , (��^9 (��^� ���^� ���^9 (��^9      C   , ��^9 ��^� ���^� ���^9 ��^9      C   , 	���^9 	���^� ���^� ���^9 	���^9      C   , ���^9 ���^� ���^� ���^9 ���^9      C   , ���^9 ���^� z��^� z��^9 ���^9      C   , ���^9 ���^� ^��^� ^��^9 ���^9      C   , ���^9 ���^� B��^� B��^9 ���^9      C   , d��^9 d��^� &��^� &��^9 d��^9      C   , H��^9 H��^� 
��^� 
��^9 H��^9      C   ,  �Z��]b  �Z��^  ���^  ���]b  �Z��]b      C   ,  �Z��[�  �Z��\�  ���\�  ���[�  �Z��[�      C   ,  �Z��Z~  �Z��[(  ���[(  ���Z~  �Z��Z~      C   ,  �Z��Y  �Z��Y�  ���Y�  ���Y  �Z��Y      C   ,  �Z��W�  �Z��XD  ���XD  ���W�  �Z��W�      C   ,  �Z��V(  �Z��V�  ���V�  ���V(  �Z��V(      C   ,  ����L#  ����]?  �x��]?  �x��L#  ����L#      C   ,  ����L#  ����]?  �\��]?  �\��L#  ����L#      C   ,  ����L#  ����]?  �@��]?  �@��L#  ����L#      C   ,  �z��L#  �z��]?  �$��]?  �$��L#  �z��L#      C   ,  ^��L#  ^��]? ��]? ��L#  ^��L#      C   , B��L# B��]? ���]? ���L# B��L#      C   , &��L# &��]? ���]? ���L# &��L#      C   , 	
��L# 	
��]? 	���]? 	���L# 	
��L#      C   , ���L# ���]? ���]? ���L# ���L#      C   , ���L# ���]? |��]? |��L# ���L#      C   , ���L# ���]? `��]? `��L# ���L#      C   , ���L# ���]? D��]? D��L# ���L#      C   , ~��L# ~��]? (��]? (��L# ~��L#      C   , b��L# b��]? ��]? ��L# b��L#      C   ,  �Z��p,  �Z��p�  ���p�  ���p,  �Z��p,      C   , ���a� ���s �8��s �8��a� ���a�      C   , ���L# ���]? �8��]? �8��L# ���L#      C   , %���a� %���s &���s &���a� %���a�      C   , (���a� (���s )���s )���a� (���a�      C   , +���a� +���s ,d��s ,d��a� +���a�      C   , .���a� .���s /H��s /H��a� .���a�      C   , 1���a� 1���s 2,��s 2,��a� 1���a�      C   , 4f��a� 4f��s 5��s 5��a� 4f��a�      C   , 7J��a� 7J��s 7���s 7���a� 7J��a�      C   , :.��a� :.��s :���s :���a� :.��a�      C   , =��a� =��s =���s =���a� =��a�      C   , ?���a� ?���s @���s @���a� ?���a�      C   , B���a� B���s C���s C���a� B���a�      C   , E���a� E���s Fh��s Fh��a� E���a�      C   , H���a� H���s IL��s IL��a� H���a�      C   , K���a� K���s L0��s L0��a� K���a�      C   , Nj��a� Nj��s O��s O��a� Nj��a�      C   , QN��a� QN��s Q���s Q���a� QN��a�      C   , T2��a� T2��s T���s T���a� T2��a�      C   , W��a� W��s W���s W���a� W��a�      C   , Y���a� Y���s Z���s Z���a� Y���a�      C   , \���a� \���s ]���s ]���a� \���a�      C   , _���a� _���s `l��s `l��a� _���a�      C   , b���a� b���s cP��s cP��a� b���a�      C   , e���a� e���s f4��s f4��a� e���a�      C   , hn��a� hn��s i��s i��a� hn��a�      C   , kR��a� kR��s k���s k���a� kR��a�      C   , n6��a� n6��s n���s n���a� n6��a�      C   , q��a� q��s q���s q���a� q��a�      C   , s���a� s���s t���s t���a� s���a�      C   , v���a� v���s w���s w���a� v���a�      C   , y���a� y���s zp��s zp��a� y���a�      C   , |���a� |���s }T��s }T��a� |���a�      C   ,  *��a�  *��s  ���s  ���a�  *��a�      C   , Nj��L# Nj��]? O��]? O��L# Nj��L#      C   , #��a� #��s #���s #���a� #��a�      C   , ,���`U ,���`� .b��`� .b��`U ,���`U      C   , /���`U /���`� 1F��`� 1F��`U /���`U      C   , 2h��`U 2h��`� 4*��`� 4*��`U 2h��`U      C   , 5L��`U 5L��`� 7��`� 7��`U 5L��`U      C   , 80��`U 80��`� 9���`� 9���`U 80��`U      C   , ;��`U ;��`� <���`� <���`U ;��`U      C   , =���`U =���`� ?���`� ?���`U =���`U      C   , @���`U @���`� B���`� B���`U @���`U      C   , C���`U C���`� E���`� E���`U C���`U      C   , ,��^9 ,��^� ���^� ���^9 ,��^9      C   , !��^9 !��^� "���^� "���^9 !��^9      C   , #���^9 #���^� %���^� %���^9 #���^9      C   , &���^9 &���^� (���^� (���^9 &���^9      C   , )���^9 )���^� +~��^� +~��^9 )���^9      C   , ,���^9 ,���^� .b��^� .b��^9 ,���^9      C   , /���^9 /���^� 1F��^� 1F��^9 /���^9      C   , 2h��^9 2h��^� 4*��^� 4*��^9 2h��^9      C   , 5L��^9 5L��^� 7��^� 7��^9 5L��^9      C   , 80��^9 80��^� 9���^� 9���^9 80��^9      C   , ;��^9 ;��^� <���^� <���^9 ;��^9      C   , =���^9 =���^� ?���^� ?���^9 =���^9      C   , @���^9 @���^� B���^� B���^9 @���^9      C   , C���^9 C���^� E���^� E���^9 C���^9      C   , F���^9 F���^� Hf��^� Hf��^9 F���^9      C   , I���^9 I���^� KJ��^� KJ��^9 I���^9      C   , Ll��^9 Ll��^� N.��^� N.��^9 Ll��^9      C   , F���`U F���`� Hf��`� Hf��`U F���`U      C   , I���`U I���`� KJ��`� KJ��`U I���`U      C   , Ll��`U Ll��`� N.��`� N.��`U Ll��`U      C   , ,��`U ,��`� ���`� ���`U ,��`U      C   , !��`U !��`� "���`� "���`U !��`U      C   , #���`U #���`� %���`� %���`U #���`U      C   ,  *��L#  *��]?  ���]?  ���L#  *��L#      C   , #��L# #��]? #���]? #���L# #��L#      C   , %���L# %���]? &���]? &���L# %���L#      C   , (���L# (���]? )���]? )���L# (���L#      C   , +���L# +���]? ,d��]? ,d��L# +���L#      C   , .���L# .���]? /H��]? /H��L# .���L#      C   , 1���L# 1���]? 2,��]? 2,��L# 1���L#      C   , 4f��L# 4f��]? 5��]? 5��L# 4f��L#      C   , 7J��L# 7J��]? 7���]? 7���L# 7J��L#      C   , :.��L# :.��]? :���]? :���L# :.��L#      C   , =��L# =��]? =���]? =���L# =��L#      C   , ?���L# ?���]? @���]? @���L# ?���L#      C   , B���L# B���]? C���]? C���L# B���L#      C   , E���L# E���]? Fh��]? Fh��L# E���L#      C   , H���L# H���]? IL��]? IL��L# H���L#      C   , K���L# K���]? L0��]? L0��L# K���L#      C   , &���`U &���`� (���`� (���`U &���`U      C   , )���`U )���`� +~��`� +~��`U )���`U      C   , c���^9 c���^� eN��^� eN��^9 c���^9      C   , fp��^9 fp��^� h2��^� h2��^9 fp��^9      C   , iT��^9 iT��^� k��^� k��^9 iT��^9      C   , l8��^9 l8��^� m���^� m���^9 l8��^9      C   , o��^9 o��^� p���^� p���^9 o��^9      C   , r ��^9 r ��^� s���^� s���^9 r ��^9      C   , t���^9 t���^� v���^� v���^9 t���^9      C   , w���^9 w���^� y���^� y���^9 w���^9      C   , z���^9 z���^� |n��^� |n��^9 z���^9      C   , }���^9 }���^� R��^� R��^9 }���^9      C   , w���`U w���`� y���`� y���`U w���`U      C   , z���`U z���`� |n��`� |n��`U z���`U      C   , }���`U }���`� R��`� R��`U }���`U      C   , OP��`U OP��`� Q��`� Q��`U OP��`U      C   , R4��`U R4��`� S���`� S���`U R4��`U      C   , U��`U U��`� V���`� V���`U U��`U      C   , W���`U W���`� Y���`� Y���`U W���`U      C   , Z���`U Z���`� \���`� \���`U Z���`U      C   , ]���`U ]���`� _���`� _���`U ]���`U      C   , `���`U `���`� bj��`� bj��`U `���`U      C   , c���`U c���`� eN��`� eN��`U c���`U      C   , fp��`U fp��`� h2��`� h2��`U fp��`U      C   , iT��`U iT��`� k��`� k��`U iT��`U      C   , l8��`U l8��`� m���`� m���`U l8��`U      C   , o��`U o��`� p���`� p���`U o��`U      C   , r ��`U r ��`� s���`� s���`U r ��`U      C   , t���`U t���`� v���`� v���`U t���`U      C   , OP��^9 OP��^� Q��^� Q��^9 OP��^9      C   , R4��^9 R4��^� S���^� S���^9 R4��^9      C   , U��^9 U��^� V���^� V���^9 U��^9      C   , W���^9 W���^� Y���^� Y���^9 W���^9      C   , Z���^9 Z���^� \���^� \���^9 Z���^9      C   , ]���^9 ]���^� _���^� _���^9 ]���^9      C   , QN��L# QN��]? Q���]? Q���L# QN��L#      C   , T2��L# T2��]? T���]? T���L# T2��L#      C   , W��L# W��]? W���]? W���L# W��L#      C   , Y���L# Y���]? Z���]? Z���L# Y���L#      C   , \���L# \���]? ]���]? ]���L# \���L#      C   , _���L# _���]? `l��]? `l��L# _���L#      C   , b���L# b���]? cP��]? cP��L# b���L#      C   , e���L# e���]? f4��]? f4��L# e���L#      C   , hn��L# hn��]? i��]? i��L# hn��L#      C   , kR��L# kR��]? k���]? k���L# kR��L#      C   , n6��L# n6��]? n���]? n���L# n6��L#      C   , q��L# q��]? q���]? q���L# q��L#      C   , s���L# s���]? t���]? t���L# s���L#      C   , v���L# v���]? w���]? w���L# v���L#      C   , y���L# y���]? zp��]? zp��L# y���L#      C   , |���L# |���]? }T��]? }T��L# |���L#      C   , `���^9 `���^� bj��^� bj��^9 `���^9      C   , �z��a� �z��s �$��s �$��a� �z��a�      C   , �r��a� �r��s ���s ���a� �r��a�      C   , �V��a� �V��s � ��s � ��a� �V��a�      C   , �:��a� �:��s ����s ����a� �:��a�      C   , ���a� ���s ����s ����a� ���a�      C   , ���a� ���s ����s ����a� ���a�      C   , ����a� ����s ����s ����a� ����a�      C   , ����a� ����s �t��s �t��a� ����a�      C   , ����a� ����s �X��s �X��a� ����a�      C   , ����a� ����s �<��s �<��a� ����a�      C   , �v��a� �v��s � ��s � ��a� �v��a�      C   , �Z��a� �Z��s ���s ���a� �Z��a�      C   , �>��a� �>��s ����s ����a� �>��a�      C   , �"��a� �"��s ����s ����a� �"��a�      C   , ���a� ���s ����s ����a� ���a�      C   , ����a� ����s ����s ����a� ����a�      C   , �^��a� �^��s ���s ���a� �^��a�      C   , �B��a� �B��s ����s ����a� �B��a�      C   , �&��a� �&��s ����s ����a� �&��a�      C   , �
��a� �
��s ´��s ´��a� �
��a�      C   , ����a� ����s Ř��s Ř��a� ����a�      C   , ����a� ����s �|��s �|��a� ����a�      C   , ͚��a� ͚��s �D��s �D��a� ͚��a�      C   , ����a� ����s �x��s �x��a� ����a�      C   , ����a� ����s �\��s �\��a� ����a�      C   , ����a� ����s �@��s �@��a� ����a�      C   , ����^9 ����^� �V��^� �V��^9 ����^9      C   , �x��^9 �x��^� �:��^� �:��^9 �x��^9      C   , �\��^9 �\��^� ���^� ���^9 �\��^9      C   , �@��^9 �@��^� ���^� ���^9 �@��^9      C   , �$��^9 �$��^� ����^� ����^9 �$��^9      C   , ���^9 ���^� ����^� ����^9 ���^9      C   , ����^9 ����^� ����^� ����^9 ����^9      C   , ����^9 ����^� ����^� ����^9 ����^9      C   , ����^9 ����^� �v��^� �v��^9 ����^9      C   , �<��^9 �<��^� ����^� ����^9 �<��^9      C   , ����`U ����`� ����`� ����`U ����`U      C   , ����`U ����`� ����`� ����`U ����`U      C   , ����`U ����`� �r��`� �r��`U ����`U      C   , ����`U ����`� �V��`� �V��`U ����`U      C   , �x��`U �x��`� �:��`� �:��`U �x��`U      C   , �\��`U �\��`� ���`� ���`U �\��`U      C   , �@��`U �@��`� ���`� ���`U �@��`U      C   , �$��`U �$��`� ����`� ����`U �$��`U      C   , ���`U ���`� ����`� ����`U ���`U      C   , ����`U ����`� ����`� ����`U ����`U      C   , ����`U ����`� ����`� ����`U ����`U      C   , ����`U ����`� �v��`� �v��`U ����`U      C   , �t��`U �t��`� �6��`� �6��`U �t��`U      C   , �X��`U �X��`� ���`� ���`U �X��`U      C   , �<��`U �<��`� ����`� ����`U �<��`U      C   , � ��`U � ��`� ����`� ����`U � ��`U      C   , ���`U ���`� ����`� ����`U ���`U      C   , � ��^9 � ��^� ����^� ����^9 � ��^9      C   , ���^9 ���^� ����^� ����^9 ���^9      C   , ����^9 ����^� ����^� ����^9 ����^9      C   , ����^9 ����^� ����^� ����^9 ����^9      C   , ����^9 ����^� �r��^� �r��^9 ����^9      C   , �t��^9 �t��^� �6��^� �6��^9 �t��^9      C   , �X��^9 �X��^� ���^� ���^9 �X��^9      C   , �r��L# �r��]? ���]? ���L# �r��L#      C   , �V��L# �V��]? � ��]? � ��L# �V��L#      C   , �:��L# �:��]? ����]? ����L# �:��L#      C   , ���L# ���]? ����]? ����L# ���L#      C   , ���L# ���]? ����]? ����L# ���L#      C   , ����L# ����]? ����]? ����L# ����L#      C   , ����L# ����]? �t��]? �t��L# ����L#      C   , ����L# ����]? �X��]? �X��L# ����L#      C   , ����L# ����]? �<��]? �<��L# ����L#      C   , �v��L# �v��]? � ��]? � ��L# �v��L#      C   , �Z��L# �Z��]? ���]? ���L# �Z��L#      C   , �>��L# �>��]? ����]? ����L# �>��L#      C   , �"��L# �"��]? ����]? ����L# �"��L#      C   , ���L# ���]? ����]? ����L# ���L#      C   , ����L# ����]? ����]? ����L# ����L#      C   , ����L# ����]? �x��]? �x��L# ����L#      C   , �|��^9 �|��^� �>��^� �>��^9 �|��^9      C   , �`��^9 �`��^� �"��^� �"��^9 �`��^9      C   , ����`U ����`� �Z��`� �Z��`U ����`U      C   , �|��`U �|��`� �>��`� �>��`U �|��`U      C   , �`��`U �`��`� �"��`� �"��`U �`��`U      C   , �D��`U �D��`� ���`� ���`U �D��`U      C   , �(��`U �(��`� ����`� ����`U �(��`U      C   , ���`U ���`� ����`� ����`U ���`U      C   , ����`U ����`� Ĳ��`� Ĳ��`U ����`U      C   , ����`U ����`� ǖ��`� ǖ��`U ����`U      C   , ȸ��`U ȸ��`� �z��`� �z��`U ȸ��`U      C   , ˜��`U ˜��`� �^��`� �^��`U ˜��`U      C   , �D��^9 �D��^� ���^� ���^9 �D��^9      C   , �(��^9 �(��^� ����^� ����^9 �(��^9      C   , ���^9 ���^� ����^� ����^9 ���^9      C   , ����^9 ����^� Ĳ��^� Ĳ��^9 ����^9      C   , ����^9 ����^� ǖ��^� ǖ��^9 ����^9      C   , ȸ��^9 ȸ��^� �z��^� �z��^9 ȸ��^9      C   , ˜��^9 ˜��^� �^��^� �^��^9 ˜��^9      C   , ����^9 ����^� �Z��^� �Z��^9 ����^9      C   , ����L# ����]? �\��]? �\��L# ����L#      C   , ����L# ����]? �@��]? �@��L# ����L#      C   , �z��L# �z��]? �$��]? �$��L# �z��L#      C   , �^��L# �^��]? ���]? ���L# �^��L#      C   , �B��L# �B��]? ����]? ����L# �B��L#      C   , �&��L# �&��]? ����]? ����L# �&��L#      C   , �
��L# �
��]? ´��]? ´��L# �
��L#      C   , ����L# ����]? Ř��]? Ř��L# ����L#      C   , ����L# ����]? �|��]? �|��L# ����L#      C  , , �  31 �  3� J  3� J  31 �  31      C  , , �  1� �  2s J  2s J  1� �  1�      C  , , �  0a �  1 J  1 J  0a �  0a      C  , , �  .� �  /� J  /� J  .� �  .�      C  , , �  -� �  .; J  .; J  -� �  -�      C  , , �  ,) �  ,� J  ,� J  ,) �  ,)      C  , , �  *� �  +k J  +k J  *� �  *�      C  , , �  )Y �  * J  * J  )Y �  )Y      C  , , �  "� �  #� J  #� J  "� �  "�      C  , , �  !u �  " J  " J  !u �  !u      C  , , �    �   � J   � J    �         C  , , �  � �  O J  O J  � �  �      C  , , �  = �  � J  � J  = �  =      C  , , �  � �   J   J  � �  �      C  , , �  m �   J   J  m �  m      C  , , �   �  � J  � J   �        C  , ,  ]����E  ]�����  ^�����  ^����E  ]����E      C  , ,  `@���E  `@����  `�����  `����E  `@���E      C  , ,  b����E  b�����  c8����  c8���E  b����E      C  , ,  d����E  d�����  e�����  e����E  d����E      C  , ,  g*���E  g*����  g�����  g����E  g*���E      C  , ,  ix���E  ix����  j"����  j"���E  ix���E      C  , ,  k����E  k�����  lp����  lp���E  k����E      C  , ,  n���E  n����  n�����  n����E  n���E      C  , ,  pb���E  pb����  q����  q���E  pb���E      C  , ,  r����E  r�����  sZ����  sZ���E  r����E      C  , ,  t����E  t�����  u�����  u����E  t����E      C  , ,  wL���E  wL����  w�����  w����E  wL���E      C  , ,  y����E  y�����  zD����  zD���E  y����E      C  , ,  {����E  {�����  |�����  |����E  {����E      C  , ,  ~6���E  ~6����  ~�����  ~����E  ~6���E      C  , ,  �����E  ������  �.����  �.���E  �����E      C  , ,  �����E  ������  �|����  �|���E  �����E      C  , ,  � ���E  � ����  ������  �����E  � ���E      C  , ,  �n���E  �n����  �����  ����E  �n���E      C  , ,  �����E  ������  �f����  �f���E  �����E      C  , ,  �
���E  �
����  ������  �����E  �
���E      C  , ,  �X���E  �X����  �����  ����E  �X���E      C  , ,  �����E  ������  �P����  �P���E  �����E      C  , ,  �����E  ������  ������  �����E  �����E      C  , ,  �B���E  �B����  ������  �����E  �B���E      C  , ,  �����E  ������  �:����  �:���E  �����E      C  , ,  �����E  ������  ������  �����E  �����E      C  , ,  �,���E  �,����  ������  �����E  �,���E      C  , ,  �z���E  �z����  �$����  �$���E  �z���E      C  , ,  �����E  ������  �r����  �r���E  �����E      C  , ,  ����E  �����  ������  �����E  ����E      C  , ,  �d���E  �d����  �����  ����E  �d���E      C  , ,  �����E  ������  �\����  �\���E  �����E      C  , ,  � ���E  � ����  ������  �����E  � ���E      C  , ,  �N���E  �N����  ������  �����E  �N���E      C  , ,  �����E  ������  �F����  �F���E  �����E      C  , ,  �����E  ������  ������  �����E  �����E      C  , ,  �8���E  �8����  ������  �����E  �8���E      C  , ,  �����E  ������  �0����  �0���E  �����E      C  , ,  �����E  ������  �~����  �~���E  �����E      C  , ,  �"���E  �"����  ������  �����E  �"���E      C  , ,  �p���E  �p����  �����  ����E  �p���E      C  , ,  �����E  ������  �h����  �h���E  �����E      C  , ,  ����E  �����  ������  �����E  ����E      C  , ,  �Z���E  �Z����  �����  ����E  �Z���E      C  , ,  Ũ���E  Ũ����  �R����  �R���E  Ũ���E      C  , ,  �����E  ������  Ƞ����  Ƞ���E  �����E      C  , ,  �D���E  �D����  ������  �����E  �D���E      C  , ,  ̒���E  ̒����  �<����  �<���E  ̒���E      C  , ,  �����E  ������  ϊ����  ϊ���E  �����E      C  , ,  �.���E  �.����  ������  �����E  �.���E      C  , , F��q� F��r� ���r� ���q� F��q�      C  , , F��p� F��q0 ���q0 ���p� F��p�      C  , , F��o F��o� ���o� ���o F��o      C  , , F��m� F��n` ���n` ���m� F��m�      C  , , F��lN F��l� ���l� ���lN F��lN      C  , , F��j� F��k� ���k� ���j� F��j�      C  , , F��i~ F��j( ���j( ���i~ F��i~      C  , , F��h F��h� ���h� ���h F��h      C  , , F��f� F��gX ���gX ���f� F��f�      C  , , F��eF F��e� ���e� ���eF F��eF      C  , , F��c� F��d� ���d� ���c� F��c�      C  , , F��bv F��c  ���c  ���bv F��bv      C  , , F��\ F��\� ���\� ���\ F��\      C  , , F��Z� F��[Z ���[Z ���Z� F��Z�      C  , , F��YH F��Y� ���Y� ���YH F��YH      C  , , F��W� F��X� ���X� ���W� F��W�      C  , , F��Vx F��W" ���W" ���Vx F��Vx      C  , , F��U F��U� ���U� ���U F��U      C  , , F��S� F��TR ���TR ���S� F��S�      C  , , F��R@ F��R� ���R� ���R@ F��R@      C  , , F��P� F��Q� ���Q� ���P� F��P�      C  , , F��Op F��P ���P ���Op F��Op      C  , , F��N F��N� ���N� ���N F��N      C  , , F��L� F��MJ ���MJ ���L� F��L�      C  , , �  ') �  '� ɷ  '� ɷ  ') �  ')      C  , , �  % �  %� ɷ  %� ɷ  % �  %      C  , , ��  %] ��  & ӏ  & ӏ  %] ��  %]      C  , , �M  %] �M  & ��  & ��  %] �M  %]      C  , , յ  %] յ  & �_  & �_  %] յ  %]      C  , , �  %] �  & ��  & ��  %] �  %]      C  , , ؅  %] ؅  & �/  & �/  %] ؅  %]      C  , , ��  %] ��  & ڗ  & ڗ  %] ��  %]      C  , , �U  %] �U  & ��  & ��  %] �U  %]      C  , , ܽ  %] ܽ  & �g  & �g  %] ܽ  %]      C  , , �%  %] �%  & ��  & ��  %] �%  %]      C  , , ߍ  %] ߍ  & �7  & �7  %] ߍ  %]      C  , , ��  %] ��  & �  & �  %] ��  %]      C  , , ��  ,� ��  -A ӏ  -A ӏ  ,� ��  ,�      C  , , �M  ,� �M  -A ��  -A ��  ,� �M  ,�      C  , , յ  ,� յ  -A �_  -A �_  ,� յ  ,�      C  , , �  ,� �  -A ��  -A ��  ,� �  ,�      C  , , ؅  ,� ؅  -A �/  -A �/  ,� ؅  ,�      C  , , ��  ,� ��  -A ڗ  -A ڗ  ,� ��  ,�      C  , , �U  ,� �U  -A ��  -A ��  ,� �U  ,�      C  , , ܽ  ,� ܽ  -A �g  -A �g  ,� ܽ  ,�      C  , , �%  ,� �%  -A ��  -A ��  ,� �%  ,�      C  , , ߍ  ,� ߍ  -A �7  -A �7  ,� ߍ  ,�      C  , , ��  ,� ��  -A �  -A �  ,� ��  ,�      C  , , �  /{ �  0% ��  0% ��  /{ �  /{      C  , , ؅  /{ ؅  0% �/  0% �/  /{ ؅  /{      C  , , ��  /{ ��  0% ڗ  0% ڗ  /{ ��  /{      C  , , �U  /{ �U  0% ��  0% ��  /{ �U  /{      C  , , ܽ  /{ ܽ  0% �g  0% �g  /{ ܽ  /{      C  , , �%  /{ �%  0% ��  0% ��  /{ �%  /{      C  , , ߍ  /{ ߍ  0% �7  0% �7  /{ ߍ  /{      C  , , ��  /{ ��  0% �  0% �  /{ ��  /{      C  , , յ  .	 յ  .� �_  .� �_  .	 յ  .	      C  , , �  .	 �  .� ��  .� ��  .	 �  .	      C  , , ؅  .	 ؅  .� �/  .� �/  .	 ؅  .	      C  , , ��  .	 ��  .� ڗ  .� ڗ  .	 ��  .	      C  , , �U  .	 �U  .� ��  .� ��  .	 �U  .	      C  , , ܽ  .	 ܽ  .� �g  .� �g  .	 ܽ  .	      C  , , �%  .	 �%  .� ��  .� ��  .	 �%  .	      C  , , ߍ  .	 ߍ  .� �7  .� �7  .	 ߍ  .	      C  , , ��  .	 ��  .� �  .� �  .	 ��  .	      C  , , ��  2_ ��  3	 �  3	 �  2_ ��  2_      C  , , յ  0� յ  1� �_  1� �_  0� յ  0�      C  , , �  0� �  1� ��  1� ��  0� �  0�      C  , , ؅  0� ؅  1� �/  1� �/  0� ؅  0�      C  , , ��  0� ��  1� ڗ  1� ڗ  0� ��  0�      C  , , �U  0� �U  1� ��  1� ��  0� �U  0�      C  , , ܽ  0� ܽ  1� �g  1� �g  0� ܽ  0�      C  , , �%  0� �%  1� ��  1� ��  0� �%  0�      C  , , ߍ  0� ߍ  1� �7  1� �7  0� ߍ  0�      C  , , ��  0� ��  1� �  1� �  0� ��  0�      C  , , յ  /{ յ  0% �_  0% �_  /{ յ  /{      C  , , յ  2_ յ  3	 �_  3	 �_  2_ յ  2_      C  , , �  2_ �  3	 ��  3	 ��  2_ �  2_      C  , , ؅  2_ ؅  3	 �/  3	 �/  2_ ؅  2_      C  , , ��  2_ ��  3	 ڗ  3	 ڗ  2_ ��  2_      C  , , �U  2_ �U  3	 ��  3	 ��  2_ �U  2_      C  , , ܽ  2_ ܽ  3	 �g  3	 �g  2_ ܽ  2_      C  , , �%  2_ �%  3	 ��  3	 ��  2_ �%  2_      C  , , ߍ  2_ ߍ  3	 �7  3	 �7  2_ ߍ  2_      C  , , յ  3� յ  4{ �_  4{ �_  3� յ  3�      C  , , �  3� �  4{ ��  4{ ��  3� �  3�      C  , , ؅  3� ؅  4{ �/  4{ �/  3� ؅  3�      C  , , ��  3� ��  4{ ڗ  4{ ڗ  3� ��  3�      C  , , �U  3� �U  4{ ��  4{ ��  3� �U  3�      C  , , ܽ  3� ܽ  4{ �g  4{ �g  3� ܽ  3�      C  , , �%  3� �%  4{ ��  4{ ��  3� �%  3�      C  , , ߍ  3� ߍ  4{ �7  4{ �7  3� ߍ  3�      C  , , ��  3� ��  4{ �  4{ �  3� ��  3�      C  , , ��  1� ��  2s �z  2s �z  1� ��  1�      C  , , ��  2_ ��  3	 ӏ  3	 ӏ  2_ ��  2_      C  , , �M  2_ �M  3	 ��  3	 ��  2_ �M  2_      C  , , ��  0� ��  1� ӏ  1� ӏ  0� ��  0�      C  , , �4  .� �4  /� ��  /� ��  .� �4  .�      C  , , ̂  .� ̂  /� �,  /� �,  .� ̂  .�      C  , , ��  .� ��  /� �z  /� �z  .� ��  .�      C  , , ��  /{ ��  0% ӏ  0% ӏ  /{ ��  /{      C  , , �4  -� �4  .; ��  .; ��  -� �4  -�      C  , , ̂  -� ̂  .; �,  .; �,  -� ̂  -�      C  , , ��  -� ��  .; �z  .; �z  -� ��  -�      C  , , �4  31 �4  3� ��  3� ��  31 �4  31      C  , , ̂  31 ̂  3� �,  3� �,  31 ̂  31      C  , , ��  31 ��  3� �z  3� �z  31 ��  31      C  , , ��  3� ��  4{ ӏ  4{ ӏ  3� ��  3�      C  , , �M  3� �M  4{ ��  4{ ��  3� �M  3�      C  , , ��  .	 ��  .� ӏ  .� ӏ  .	 ��  .	      C  , , �M  .	 �M  .� ��  .� ��  .	 �M  .	      C  , , �M  /{ �M  0% ��  0% ��  /{ �M  /{      C  , , �M  0� �M  1� ��  1� ��  0� �M  0�      C  , , �4  0a �4  1 ��  1 ��  0a �4  0a      C  , , ̂  0a ̂  1 �,  1 �,  0a ̂  0a      C  , , ��  0a ��  1 �z  1 �z  0a ��  0a      C  , , �4  1� �4  2s ��  2s ��  1� �4  1�      C  , , ̂  1� ̂  2s �,  2s �,  1� ̂  1�      C  , , �4  )Y �4  * ��  * ��  )Y �4  )Y      C  , , ̂  )Y ̂  * �,  * �,  )Y ̂  )Y      C  , , ��  )Y ��  * �z  * �z  )Y ��  )Y      C  , , ��  )� ��  *] ӏ  *] ӏ  )� ��  )�      C  , , �M  )� �M  *] ��  *] ��  )� �M  )�      C  , , ��  (A ��  (� ӏ  (� ӏ  (A ��  (A      C  , , �M  (A �M  (� ��  (� ��  (A �M  (A      C  , , ��  ,) ��  ,� �z  ,� �z  ,) ��  ,)      C  , , �[  ') �[  '� �  '� �  ') �[  ')      C  , , ͩ  ') ͩ  '� �S  '� �S  ') ͩ  ')      C  , , ��  &� ��  'y ӏ  'y ӏ  &� ��  &�      C  , , �M  &� �M  'y ��  'y ��  &� �M  &�      C  , , �4  ,) �4  ,� ��  ,� ��  ,) �4  ,)      C  , , ̂  ,) ̂  ,� �,  ,� �,  ,) ̂  ,)      C  , , �4  *� �4  +k ��  +k ��  *� �4  *�      C  , , ̂  *� ̂  +k �,  +k �,  *� ̂  *�      C  , , ��  *� ��  +k �z  +k �z  *� ��  *�      C  , , ��  +% ��  +� ӏ  +� ӏ  +% ��  +%      C  , , �M  +% �M  +� ��  +� ��  +% �M  +%      C  , , ؅  +% ؅  +� �/  +� �/  +% ؅  +%      C  , , յ  &� յ  'y �_  'y �_  &� յ  &�      C  , , �  &� �  'y ��  'y ��  &� �  &�      C  , , ؅  &� ؅  'y �/  'y �/  &� ؅  &�      C  , , ��  &� ��  'y ڗ  'y ڗ  &� ��  &�      C  , , �U  &� �U  'y ��  'y ��  &� �U  &�      C  , , ܽ  &� ܽ  'y �g  'y �g  &� ܽ  &�      C  , , �%  &� �%  'y ��  'y ��  &� �%  &�      C  , , ߍ  &� ߍ  'y �7  'y �7  &� ߍ  &�      C  , , ��  &� ��  'y �  'y �  &� ��  &�      C  , , ��  +% ��  +� ڗ  +� ڗ  +% ��  +%      C  , , �U  +% �U  +� ��  +� ��  +% �U  +%      C  , , յ  )� յ  *] �_  *] �_  )� յ  )�      C  , , �  )� �  *] ��  *] ��  )� �  )�      C  , , ؅  )� ؅  *] �/  *] �/  )� ؅  )�      C  , , ��  )� ��  *] ڗ  *] ڗ  )� ��  )�      C  , , �U  )� �U  *] ��  *] ��  )� �U  )�      C  , , ܽ  )� ܽ  *] �g  *] �g  )� ܽ  )�      C  , , �%  )� �%  *] ��  *] ��  )� �%  )�      C  , , ߍ  )� ߍ  *] �7  *] �7  )� ߍ  )�      C  , , ��  )� ��  *] �  *] �  )� ��  )�      C  , , ܽ  +% ܽ  +� �g  +� �g  +% ܽ  +%      C  , , �%  +% �%  +� ��  +� ��  +% �%  +%      C  , , յ  (A յ  (� �_  (� �_  (A յ  (A      C  , , �  (A �  (� ��  (� ��  (A �  (A      C  , , ؅  (A ؅  (� �/  (� �/  (A ؅  (A      C  , , ��  (A ��  (� ڗ  (� ڗ  (A ��  (A      C  , , �U  (A �U  (� ��  (� ��  (A �U  (A      C  , , ܽ  (A ܽ  (� �g  (� �g  (A ܽ  (A      C  , , �%  (A �%  (� ��  (� ��  (A �%  (A      C  , , ߍ  (A ߍ  (� �7  (� �7  (A ߍ  (A      C  , , ��  (A ��  (� �  (� �  (A ��  (A      C  , , ߍ  +% ߍ  +� �7  +� �7  +% ߍ  +%      C  , , ��  +% ��  +� �  +� �  +% ��  +%      C  , , յ  +% յ  +� �_  +� �_  +% յ  +%      C  , , �  +% �  +� ��  +� ��  +% �  +%      C  , , �J  -� �J  .; ��  .; ��  -� �J  -�      C  , , ��  )Y ��  * ��  * ��  )Y ��  )Y      C  , , �(  )Y �(  * ��  * ��  )Y �(  )Y      C  , , �v  )Y �v  * �   * �   )Y �v  )Y      C  , , ��  )Y ��  * �n  * �n  )Y ��  )Y      C  , , �  )Y �  * ��  * ��  )Y �  )Y      C  , , �`  )Y �`  * �
  * �
  )Y �`  )Y      C  , , ��  )Y ��  * �X  * �X  )Y ��  )Y      C  , , ��  )Y ��  * ��  * ��  )Y ��  )Y      C  , , �J  )Y �J  * ��  * ��  )Y �J  )Y      C  , , Ř  )Y Ř  * �B  * �B  )Y Ř  )Y      C  , , ��  )Y ��  * Ȑ  * Ȑ  )Y ��  )Y      C  , , Ř  -� Ř  .; �B  .; �B  -� Ř  -�      C  , , ��  -� ��  .; Ȑ  .; Ȑ  -� ��  -�      C  , , Ř  1� Ř  2s �B  2s �B  1� Ř  1�      C  , , ��  1� ��  2s Ȑ  2s Ȑ  1� ��  1�      C  , , ��  1� ��  2s ��  2s ��  1� ��  1�      C  , , �(  1� �(  2s ��  2s ��  1� �(  1�      C  , , �v  1� �v  2s �   2s �   1� �v  1�      C  , , ��  0a ��  1 ��  1 ��  0a ��  0a      C  , , �(  0a �(  1 ��  1 ��  0a �(  0a      C  , , �v  0a �v  1 �   1 �   0a �v  0a      C  , , ��  .� ��  /� ��  /� ��  .� ��  .�      C  , , �(  .� �(  /� ��  /� ��  .� �(  .�      C  , , �v  .� �v  /� �   /� �   .� �v  .�      C  , , ��  .� ��  /� �n  /� �n  .� ��  .�      C  , , �  .� �  /� ��  /� ��  .� �  .�      C  , , �`  .� �`  /� �
  /� �
  .� �`  .�      C  , , ��  ,) ��  ,� ��  ,� ��  ,) ��  ,)      C  , , �(  ,) �(  ,� ��  ,� ��  ,) �(  ,)      C  , , �v  ,) �v  ,� �   ,� �   ,) �v  ,)      C  , , ��  ,) ��  ,� �n  ,� �n  ,) ��  ,)      C  , , �  ,) �  ,� ��  ,� ��  ,) �  ,)      C  , , �`  ,) �`  ,� �
  ,� �
  ,) �`  ,)      C  , , ��  ,) ��  ,� �X  ,� �X  ,) ��  ,)      C  , , ��  ,) ��  ,� ��  ,� ��  ,) ��  ,)      C  , , �J  ,) �J  ,� ��  ,� ��  ,) �J  ,)      C  , , �  ') �  '� ��  '� ��  ') �  ')      C  , , �O  ') �O  '� ��  '� ��  ') �O  ')      C  , , ��  ') ��  '� �G  '� �G  ') ��  ')      C  , , ��  ') ��  '� ��  '� ��  ') ��  ')      C  , , �9  ') �9  '� ��  '� ��  ') �9  ')      C  , , ��  ') ��  '� �1  '� �1  ') ��  ')      C  , , ��  ') ��  '� �  '� �  ') ��  ')      C  , , �#  ') �#  '� ��  '� ��  ') �#  ')      C  , , �q  ') �q  '� �  '� �  ') �q  ')      C  , , ƿ  ') ƿ  '� �i  '� �i  ') ƿ  ')      C  , , Ř  ,) Ř  ,� �B  ,� �B  ,) Ř  ,)      C  , , ��  ,) ��  ,� Ȑ  ,� Ȑ  ,) ��  ,)      C  , , ��  .� ��  /� �X  /� �X  .� ��  .�      C  , , ��  .� ��  /� ��  /� ��  .� ��  .�      C  , , �J  .� �J  /� ��  /� ��  .� �J  .�      C  , , Ř  .� Ř  /� �B  /� �B  .� Ř  .�      C  , , ��  .� ��  /� Ȑ  /� Ȑ  .� ��  .�      C  , , ��  0a ��  1 �n  1 �n  0a ��  0a      C  , , �  0a �  1 ��  1 ��  0a �  0a      C  , , �`  0a �`  1 �
  1 �
  0a �`  0a      C  , , ��  0a ��  1 �X  1 �X  0a ��  0a      C  , , ��  0a ��  1 ��  1 ��  0a ��  0a      C  , , �J  0a �J  1 ��  1 ��  0a �J  0a      C  , , Ř  0a Ř  1 �B  1 �B  0a Ř  0a      C  , , ��  0a ��  1 Ȑ  1 Ȑ  0a ��  0a      C  , , ��  1� ��  2s �n  2s �n  1� ��  1�      C  , , ��  *� ��  +k ��  +k ��  *� ��  *�      C  , , �(  *� �(  +k ��  +k ��  *� �(  *�      C  , , �v  *� �v  +k �   +k �   *� �v  *�      C  , , ��  *� ��  +k �n  +k �n  *� ��  *�      C  , , �  *� �  +k ��  +k ��  *� �  *�      C  , , �`  *� �`  +k �
  +k �
  *� �`  *�      C  , , ��  *� ��  +k �X  +k �X  *� ��  *�      C  , , ��  *� ��  +k ��  +k ��  *� ��  *�      C  , , �J  *� �J  +k ��  +k ��  *� �J  *�      C  , , Ř  *� Ř  +k �B  +k �B  *� Ř  *�      C  , , ��  31 ��  3� ��  3� ��  31 ��  31      C  , , �(  31 �(  3� ��  3� ��  31 �(  31      C  , , �v  31 �v  3� �   3� �   31 �v  31      C  , , ��  31 ��  3� �n  3� �n  31 ��  31      C  , , �  31 �  3� ��  3� ��  31 �  31      C  , , �`  31 �`  3� �
  3� �
  31 �`  31      C  , , ��  31 ��  3� �X  3� �X  31 ��  31      C  , , ��  31 ��  3� ��  3� ��  31 ��  31      C  , , �J  31 �J  3� ��  3� ��  31 �J  31      C  , , Ř  31 Ř  3� �B  3� �B  31 Ř  31      C  , , ��  31 ��  3� Ȑ  3� Ȑ  31 ��  31      C  , , ��  *� ��  +k Ȑ  +k Ȑ  *� ��  *�      C  , , �  1� �  2s ��  2s ��  1� �  1�      C  , , �`  1� �`  2s �
  2s �
  1� �`  1�      C  , , ��  1� ��  2s �X  2s �X  1� ��  1�      C  , , ��  1� ��  2s ��  2s ��  1� ��  1�      C  , , �J  1� �J  2s ��  2s ��  1� �J  1�      C  , , ��  -� ��  .; ��  .; ��  -� ��  -�      C  , , �(  -� �(  .; ��  .; ��  -� �(  -�      C  , , �v  -� �v  .; �   .; �   -� �v  -�      C  , , ��  -� ��  .; �n  .; �n  -� ��  -�      C  , , �  -� �  .; ��  .; ��  -� �  -�      C  , , �`  -� �`  .; �
  .; �
  -� �`  -�      C  , , ��  -� ��  .; �X  .; �X  -� ��  -�      C  , , ��  -� ��  .; ��  .; ��  -� ��  -�      C  , , �  !u �  " ��  " ��  !u �  !u      C  , , �`  !u �`  " �
  " �
  !u �`  !u      C  , , ��  !u ��  " �X  " �X  !u ��  !u      C  , , ��  !u ��  " ��  " ��  !u ��  !u      C  , , �J  !u �J  " ��  " ��  !u �J  !u      C  , , Ř  !u Ř  " �B  " �B  !u Ř  !u      C  , , ��  !u ��  " Ȑ  " Ȑ  !u ��  !u      C  , , ��    ��   � ��   � ��    ��         C  , , �(    �(   � ��   � ��    �(         C  , , �v    �v   � �    � �     �v         C  , , ��    ��   � �n   � �n    ��         C  , , �    �   � ��   � ��    �         C  , , �`    �`   � �
   � �
    �`         C  , , ��    ��   � �X   � �X    ��         C  , , ��    ��   � ��   � ��    ��         C  , , �J    �J   � ��   � ��    �J         C  , , Ř    Ř   � �B   � �B    Ř         C  , , ��    ��   � Ȑ   � Ȑ    ��         C  , , ��  � ��  O ��  O ��  � ��  �      C  , , �(  � �(  O ��  O ��  � �(  �      C  , , �v  � �v  O �   O �   � �v  �      C  , , ��  � ��  O �n  O �n  � ��  �      C  , , �  � �  O ��  O ��  � �  �      C  , , �`  � �`  O �
  O �
  � �`  �      C  , , ��  � ��  O �X  O �X  � ��  �      C  , , ��  � ��  O ��  O ��  � ��  �      C  , , �J  � �J  O ��  O ��  � �J  �      C  , , Ř  � Ř  O �B  O �B  � Ř  �      C  , , ��  � ��  O Ȑ  O Ȑ  � ��  �      C  , , ��  = ��  � ��  � ��  = ��  =      C  , , �(  = �(  � ��  � ��  = �(  =      C  , , �v  = �v  � �   � �   = �v  =      C  , , ��  = ��  � �n  � �n  = ��  =      C  , , �  = �  � ��  � ��  = �  =      C  , , �`  = �`  � �
  � �
  = �`  =      C  , , ��  = ��  � �X  � �X  = ��  =      C  , , ��  = ��  � ��  � ��  = ��  =      C  , , �J  = �J  � ��  � ��  = �J  =      C  , , Ř  = Ř  � �B  � �B  = Ř  =      C  , , ��  = ��  � Ȑ  � Ȑ  = ��  =      C  , , ��  � ��   ��   ��  � ��  �      C  , , �(  � �(   ��   ��  � �(  �      C  , , �v  � �v   �    �   � �v  �      C  , , ��  � ��   �n   �n  � ��  �      C  , , �  � �   ��   ��  � �  �      C  , , �`  � �`   �
   �
  � �`  �      C  , , ��  � ��   �X   �X  � ��  �      C  , , ��  � ��   ��   ��  � ��  �      C  , , �J  � �J   ��   ��  � �J  �      C  , , Ř  � Ř   �B   �B  � Ř  �      C  , , ��  � ��   Ȑ   Ȑ  � ��  �      C  , , ��  m ��   ��   ��  m ��  m      C  , , �(  m �(   ��   ��  m �(  m      C  , , �v  m �v   �    �   m �v  m      C  , , ��  m ��   �n   �n  m ��  m      C  , , �  m �   ��   ��  m �  m      C  , , �`  m �`   �
   �
  m �`  m      C  , , ��  m ��   �X   �X  m ��  m      C  , , ��  m ��   ��   ��  m ��  m      C  , , �J  m �J   ��   ��  m �J  m      C  , , Ř  m Ř   �B   �B  m Ř  m      C  , , ��  m ��   Ȑ   Ȑ  m ��  m      C  , , ��   ��  � ��  � ��   ��        C  , , �(   �(  � ��  � ��   �(        C  , , �v   �v  � �   � �    �v        C  , , ��   ��  � �n  � �n   ��        C  , , �   �  � ��  � ��   �        C  , , �`   �`  � �
  � �
   �`        C  , , ��   ��  � �X  � �X   ��        C  , , ��   ��  � ��  � ��   ��        C  , , �J   �J  � ��  � ��   �J        C  , , Ř   Ř  � �B  � �B   Ř        C  , , ��   ��  � Ȑ  � Ȑ   ��        C  , , ��  % ��  %� �G  %� �G  % ��  %      C  , , ��  % ��  %� ��  %� ��  % ��  %      C  , , �9  % �9  %� ��  %� ��  % �9  %      C  , , ��  % ��  %� �1  %� �1  % ��  %      C  , , ��  % ��  %� �  %� �  % ��  %      C  , , �#  % �#  %� ��  %� ��  % �#  %      C  , , �q  % �q  %� �  %� �  % �q  %      C  , , ƿ  % ƿ  %� �i  %� �i  % ƿ  %      C  , , �  % �  %� ��  %� ��  % �  %      C  , , �O  % �O  %� ��  %� ��  % �O  %      C  , , ��  "� ��  #� ��  #� ��  "� ��  "�      C  , , �(  "� �(  #� ��  #� ��  "� �(  "�      C  , , �v  "� �v  #� �   #� �   "� �v  "�      C  , , ��  "� ��  #� �n  #� �n  "� ��  "�      C  , , �  "� �  #� ��  #� ��  "� �  "�      C  , , �`  "� �`  #� �
  #� �
  "� �`  "�      C  , , ��  "� ��  #� �X  #� �X  "� ��  "�      C  , , ��  "� ��  #� ��  #� ��  "� ��  "�      C  , , �J  "� �J  #� ��  #� ��  "� �J  "�      C  , , Ř  "� Ř  #� �B  #� �B  "� Ř  "�      C  , , ��  "� ��  #� Ȑ  #� Ȑ  "� ��  "�      C  , , ��  !u ��  " ��  " ��  !u ��  !u      C  , , �(  !u �(  " ��  " ��  !u �(  !u      C  , , �v  !u �v  " �   " �   !u �v  !u      C  , , ��  !u ��  " �n  " �n  !u ��  !u      C  , , �4  � �4  O ��  O ��  � �4  �      C  , , ̂  � ̂  O �,  O �,  � ̂  �      C  , , ��  � ��  O �z  O �z  � ��  �      C  , , ��  # ��  � ӏ  � ӏ  # ��  #      C  , , �M  # �M  � ��  � ��  # �M  #      C  , , յ  # յ  � �_  � �_  # յ  #      C  , , �  # �  � ��  � ��  # �  #      C  , , ؅  # ؅  � �/  � �/  # ؅  #      C  , , ��  # ��  � ڗ  � ڗ  # ��  #      C  , , �U  # �U  � ��  � ��  # �U  #      C  , , ܽ  # ܽ  � �g  � �g  # ܽ  #      C  , , �%  # �%  � ��  � ��  # �%  #      C  , , ߍ  # ߍ  � �7  � �7  # ߍ  #      C  , , ��  # ��  � �  � �  # ��  #      C  , , ܽ  #� ܽ  $� �g  $� �g  #� ܽ  #�      C  , , �%  #� �%  $� ��  $� ��  #� �%  #�      C  , , յ  "y յ  ## �_  ## �_  "y յ  "y      C  , , �  "y �  ## ��  ## ��  "y �  "y      C  , , ؅  "y ؅  ## �/  ## �/  "y ؅  "y      C  , , ��  "y ��  ## ڗ  ## ڗ  "y ��  "y      C  , , յ  � յ   ? �_   ? �_  � յ  �      C  , , �  � �   ? ��   ? ��  � �  �      C  , , ؅  � ؅   ? �/   ? �/  � ؅  �      C  , , ��  � ��   ? ڗ   ? ڗ  � ��  �      C  , , �U  � �U   ? ��   ? ��  � �U  �      C  , , ܽ  � ܽ   ? �g   ? �g  � ܽ  �      C  , , �%  � �%   ? ��   ? ��  � �%  �      C  , , ߍ  � ߍ   ? �7   ? �7  � ߍ  �      C  , , ��  � ��   ? �   ? �  � ��  �      C  , , �U  "y �U  ## ��  ## ��  "y �U  "y      C  , , ܽ  "y ܽ  ## �g  ## �g  "y ܽ  "y      C  , , �%  "y �%  ## ��  ## ��  "y �%  "y      C  , , ߍ  "y ߍ  ## �7  ## �7  "y ߍ  "y      C  , , ��  "y ��  ## �  ## �  "y ��  "y      C  , , ߍ  #� ߍ  $� �7  $� �7  #� ߍ  #�      C  , , ��  #� ��  $� �  $� �  #� ��  #�      C  , , յ  #� յ  $� �_  $� �_  #� յ  #�      C  , , �  #� �  $� ��  $� ��  #� �  #�      C  , , ؅  #� ؅  $� �/  $� �/  #� ؅  #�      C  , , ��  #� ��  $� ڗ  $� ڗ  #� ��  #�      C  , , �U  #� �U  $� ��  $� ��  #� �U  #�      C  , , յ  ! յ  !� �_  !� �_  ! յ  !      C  , , �  ! �  !� ��  !� ��  ! �  !      C  , , ؅  ! ؅  !� �/  !� �/  ! ؅  !      C  , , ��  ! ��  !� ڗ  !� ڗ  ! ��  !      C  , , �U  ! �U  !� ��  !� ��  ! �U  !      C  , , ܽ  ! ܽ  !� �g  !� �g  ! ܽ  !      C  , , �%  ! �%  !� ��  !� ��  ! �%  !      C  , , ߍ  ! ߍ  !� �7  !� �7  ! ߍ  !      C  , , ��  ! ��  !� �  !� �  ! ��  !      C  , , �4  !u �4  " ��  " ��  !u �4  !u      C  , , ͩ  % ͩ  %� �S  %� �S  % ͩ  %      C  , , �[  % �[  %� �  %� �  % �[  %      C  , , ��  #� ��  $� ӏ  $� ӏ  #� ��  #�      C  , , �M  #� �M  $� ��  $� ��  #� �M  #�      C  , , �4  "� �4  #� ��  #� ��  "� �4  "�      C  , , ̂  "� ̂  #� �,  #� �,  "� ̂  "�      C  , , ��  "� ��  #� �z  #� �z  "� ��  "�      C  , , ��  "y ��  ## ӏ  ## ӏ  "y ��  "y      C  , , �M  "y �M  ## ��  ## ��  "y �M  "y      C  , , ̂  !u ̂  " �,  " �,  !u ̂  !u      C  , , ��  !u ��  " �z  " �z  !u ��  !u      C  , , ��  ! ��  !� ӏ  !� ӏ  ! ��  !      C  , , �M  ! �M  !� ��  !� ��  ! �M  !      C  , , �4    �4   � ��   � ��    �4         C  , , ̂    ̂   � �,   � �,    ̂         C  , , ��    ��   � �z   � �z    ��         C  , , ��  � ��   ? ӏ   ? ӏ  � ��  �      C  , , �M  � �M   ? ��   ? ��  � �M  �      C  , , ��  � ��  [ ӏ  [ ӏ  � ��  �      C  , , �M  � �M  [ ��  [ ��  � �M  �      C  , , �4  = �4  � ��  � ��  = �4  =      C  , , �4  � �4   ��   ��  � �4  �      C  , , ̂  � ̂   �,   �,  � ̂  �      C  , , ��  � ��   �z   �z  � ��  �      C  , , ��  ? ��  � ӏ  � ӏ  ? ��  ?      C  , , �M  ? �M  � ��  � ��  ? �M  ?      C  , , ̂  = ̂  � �,  � �,  = ̂  =      C  , , �4  m �4   ��   ��  m �4  m      C  , , �4   �4  � ��  � ��   �4        C  , , ̂   ̂  � �,  � �,   ̂        C  , , ��   ��  � �z  � �z   ��        C  , , ��  [ ��   ӏ   ӏ  [ ��  [      C  , , �M  [ �M   ��   ��  [ �M  [      C  , , ̂  m ̂   �,   �,  m ̂  m      C  , , ��  m ��   �z   �z  m ��  m      C  , , ��  � ��  w ӏ  w ӏ  � ��  �      C  , , �M  � �M  w ��  w ��  � �M  �      C  , , ��  = ��  � �z  � �z  = ��  =      C  , , ��  ? ��  � ڗ  � ڗ  ? ��  ?      C  , , �U  ? �U  � ��  � ��  ? �U  ?      C  , , յ  [ յ   �_   �_  [ յ  [      C  , , �  [ �   ��   ��  [ �  [      C  , , ؅  [ ؅   �/   �/  [ ؅  [      C  , , ��  [ ��   ڗ   ڗ  [ ��  [      C  , , �U  [ �U   ��   ��  [ �U  [      C  , , ܽ  [ ܽ   �g   �g  [ ܽ  [      C  , , �%  [ �%   ��   ��  [ �%  [      C  , , ߍ  [ ߍ   �7   �7  [ ߍ  [      C  , , ��  [ ��   �   �  [ ��  [      C  , , ܽ  ? ܽ  � �g  � �g  ? ܽ  ?      C  , , �%  ? �%  � ��  � ��  ? �%  ?      C  , , յ  � յ  w �_  w �_  � յ  �      C  , , �  � �  w ��  w ��  � �  �      C  , , ؅  � ؅  w �/  w �/  � ؅  �      C  , , ��  � ��  w ڗ  w ڗ  � ��  �      C  , , �U  � �U  w ��  w ��  � �U  �      C  , , ܽ  � ܽ  w �g  w �g  � ܽ  �      C  , , �%  � �%  w ��  w ��  � �%  �      C  , , ߍ  � ߍ  w �7  w �7  � ߍ  �      C  , , ��  � ��  w �  w �  � ��  �      C  , , ߍ  ? ߍ  � �7  � �7  ? ߍ  ?      C  , , ��  ? ��  � �  � �  ? ��  ?      C  , , ߍ  � ߍ  [ �7  [ �7  � ߍ  �      C  , , ��  � ��  [ �  [ �  � ��  �      C  , , յ  � յ  [ �_  [ �_  � յ  �      C  , , �  � �  [ ��  [ ��  � �  �      C  , , ؅  � ؅  [ �/  [ �/  � ؅  �      C  , , ��  � ��  [ ڗ  [ ڗ  � ��  �      C  , , �U  � �U  [ ��  [ ��  � �U  �      C  , , ܽ  � ܽ  [ �g  [ �g  � ܽ  �      C  , , �%  � �%  [ ��  [ ��  � �%  �      C  , , յ  ? յ  � �_  � �_  ? յ  ?      C  , , �  ? �  � ��  � ��  ? �  ?      C  , , ؅  ? ؅  � �/  � �/  ? ؅  ?      C  , , �^  %] �^  & �  & �  %] �^  %]      C  , , ��  %] ��  & �p  & �p  %] ��  %]      C  , , �.  %] �.  & ��  & ��  %] �.  %]      C  , , ��  %] ��  & �@  & �@  %] ��  %]      C  , , ��  %] ��  & ��  & ��  %] ��  %]      C  , , �f  %] �f  & �  & �  %] �f  %]      C  , , ��  %] ��  & �x  & �x  %] ��  %]      C  , , �6  %] �6  & ��  & ��  %] �6  %]      C  , , ��  %] ��  & �H  & �H  %] ��  %]      C  , , �  %] �  & ��  & ��  %] �  %]      C  , , �n  %] �n  & �  & �  %] �n  %]      C  , , ��  1� ��  2s �x  2s �x  1� ��  1�      C  , , ��  -� ��  .; �x  .; �x  -� ��  -�      C  , , ��  )Y ��  * �x  * �x  )Y ��  )Y      C  , , �  )Y �  * ��  * ��  )Y �  )Y      C  , , �j  )Y �j  * �  * �  )Y �j  )Y      C  , , ��  )Y ��  * �b  * �b  )Y ��  )Y      C  , , �  )Y �  * ��  * ��  )Y �  )Y      C  , , �T  )Y �T  * ��  * ��  )Y �T  )Y      C  , , ��  )Y ��  * �L  * �L  )Y ��  )Y      C  , , ��  )Y ��  * ��  * ��  )Y ��  )Y      C  , , �>  )Y �>  * ��  * ��  )Y �>  )Y      C  , , ��  )Y ��  * �6  * �6  )Y ��  )Y      C  , , �  -� �  .; ��  .; ��  -� �  -�      C  , , �j  -� �j  .; �  .; �  -� �j  -�      C  , , ��  -� ��  .; �b  .; �b  -� ��  -�      C  , , �  -� �  .; ��  .; ��  -� �  -�      C  , , �T  -� �T  .; ��  .; ��  -� �T  -�      C  , , ��  -� ��  .; �L  .; �L  -� ��  -�      C  , , ��  -� ��  .; ��  .; ��  -� ��  -�      C  , , �>  -� �>  .; ��  .; ��  -� �>  -�      C  , , ��  -� ��  .; �6  .; �6  -� ��  -�      C  , , �  1� �  2s ��  2s ��  1� �  1�      C  , , �j  1� �j  2s �  2s �  1� �j  1�      C  , , ��  1� ��  2s �b  2s �b  1� ��  1�      C  , , �  1� �  2s ��  2s ��  1� �  1�      C  , , �T  1� �T  2s ��  2s ��  1� �T  1�      C  , , ��  1� ��  2s �L  2s �L  1� ��  1�      C  , , ��  1� ��  2s ��  2s ��  1� ��  1�      C  , , �>  1� �>  2s ��  2s ��  1� �>  1�      C  , , ��  1� ��  2s �6  2s �6  1� ��  1�      C  , , ��  ') ��  '� �Q  '� �Q  ') ��  ')      C  , , ��  ') ��  '� ��  '� ��  ') ��  ')      C  , , �C  ') �C  '� ��  '� ��  ') �C  ')      C  , , ��  ') ��  '� �;  '� �;  ') ��  ')      C  , , ��  ') ��  '� ��  '� ��  ') ��  ')      C  , , �-  ') �-  '� ��  '� ��  ') �-  ')      C  , , �{  ') �{  '� �%  '� �%  ') �{  ')      C  , , ��  ') ��  '� �s  '� �s  ') ��  ')      C  , , �  ') �  '� ��  '� ��  ') �  ')      C  , , �e  ') �e  '� �  '� �  ') �e  ')      C  , , ��  ') ��  '� �]  '� �]  ') ��  ')      C  , , ��  ,) ��  ,� �x  ,� �x  ,) ��  ,)      C  , , �  ,) �  ,� ��  ,� ��  ,) �  ,)      C  , , �j  ,) �j  ,� �  ,� �  ,) �j  ,)      C  , , ��  ,) ��  ,� �b  ,� �b  ,) ��  ,)      C  , , �  ,) �  ,� ��  ,� ��  ,) �  ,)      C  , , �T  ,) �T  ,� ��  ,� ��  ,) �T  ,)      C  , , ��  ,) ��  ,� �L  ,� �L  ,) ��  ,)      C  , , ��  ,) ��  ,� ��  ,� ��  ,) ��  ,)      C  , , �>  ,) �>  ,� ��  ,� ��  ,) �>  ,)      C  , , ��  ,) ��  ,� �6  ,� �6  ,) ��  ,)      C  , , ��  .� ��  /� �x  /� �x  .� ��  .�      C  , , �  .� �  /� ��  /� ��  .� �  .�      C  , , �  *� �  +k ��  +k ��  *� �  *�      C  , , �T  *� �T  +k ��  +k ��  *� �T  *�      C  , , ��  *� ��  +k �L  +k �L  *� ��  *�      C  , , ��  *� ��  +k ��  +k ��  *� ��  *�      C  , , �>  *� �>  +k ��  +k ��  *� �>  *�      C  , , ��  *� ��  +k �6  +k �6  *� ��  *�      C  , , �T  0a �T  1 ��  1 ��  0a �T  0a      C  , , ��  0a ��  1 �L  1 �L  0a ��  0a      C  , , ��  0a ��  1 ��  1 ��  0a ��  0a      C  , , �>  0a �>  1 ��  1 ��  0a �>  0a      C  , , ��  0a ��  1 �6  1 �6  0a ��  0a      C  , , �j  .� �j  /� �  /� �  .� �j  .�      C  , , ��  .� ��  /� �b  /� �b  .� ��  .�      C  , , �  .� �  /� ��  /� ��  .� �  .�      C  , , �T  .� �T  /� ��  /� ��  .� �T  .�      C  , , ��  .� ��  /� �L  /� �L  .� ��  .�      C  , , ��  .� ��  /� ��  /� ��  .� ��  .�      C  , , �>  .� �>  /� ��  /� ��  .� �>  .�      C  , , ��  .� ��  /� �6  /� �6  .� ��  .�      C  , , ��  0a ��  1 �x  1 �x  0a ��  0a      C  , , �  0a �  1 ��  1 ��  0a �  0a      C  , , �j  0a �j  1 �  1 �  0a �j  0a      C  , , ��  0a ��  1 �b  1 �b  0a ��  0a      C  , , �  0a �  1 ��  1 ��  0a �  0a      C  , , ��  31 ��  3� �x  3� �x  31 ��  31      C  , , �  31 �  3� ��  3� ��  31 �  31      C  , , �j  31 �j  3� �  3� �  31 �j  31      C  , , ��  31 ��  3� �b  3� �b  31 ��  31      C  , , �  31 �  3� ��  3� ��  31 �  31      C  , , �T  31 �T  3� ��  3� ��  31 �T  31      C  , , ��  31 ��  3� �L  3� �L  31 ��  31      C  , , ��  31 ��  3� ��  3� ��  31 ��  31      C  , , �>  31 �>  3� ��  3� ��  31 �>  31      C  , , ��  31 ��  3� �6  3� �6  31 ��  31      C  , , ��  *� ��  +k �x  +k �x  *� ��  *�      C  , , �  *� �  +k ��  +k ��  *� �  *�      C  , , �j  *� �j  +k �  +k �  *� �j  *�      C  , , ��  *� ��  +k �b  +k �b  *� ��  *�      C  , , �.  ,� �.  -A ��  -A ��  ,� �.  ,�      C  , , ��  ,� ��  -A �@  -A �@  ,� ��  ,�      C  , , ��  ,� ��  -A ��  -A ��  ,� ��  ,�      C  , , �f  ,� �f  -A �  -A �  ,� �f  ,�      C  , , ��  ,� ��  -A �x  -A �x  ,� ��  ,�      C  , , �6  ,� �6  -A ��  -A ��  ,� �6  ,�      C  , , ��  ,� ��  -A �H  -A �H  ,� ��  ,�      C  , , �  ,� �  -A ��  -A ��  ,� �  ,�      C  , , �n  ,� �n  -A �  -A �  ,� �n  ,�      C  , , �^  ,� �^  -A �  -A �  ,� �^  ,�      C  , , ��  ,� ��  -A �p  -A �p  ,� ��  ,�      C  , , �n  2_ �n  3	 �  3	 �  2_ �n  2_      C  , , �6  2_ �6  3	 ��  3	 ��  2_ �6  2_      C  , , �6  .	 �6  .� ��  .� ��  .	 �6  .	      C  , , ��  .	 ��  .� �H  .� �H  .	 ��  .	      C  , , �  .	 �  .� ��  .� ��  .	 �  .	      C  , , �n  .	 �n  .� �  .� �  .	 �n  .	      C  , , ��  /{ ��  0% �H  0% �H  /{ ��  /{      C  , , �  /{ �  0% ��  0% ��  /{ �  /{      C  , , �n  /{ �n  0% �  0% �  /{ �n  /{      C  , , �6  0� �6  1� ��  1� ��  0� �6  0�      C  , , ��  0� ��  1� �H  1� �H  0� ��  0�      C  , , �  0� �  1� ��  1� ��  0� �  0�      C  , , �n  0� �n  1� �  1� �  0� �n  0�      C  , , �6  3� �6  4{ ��  4{ ��  3� �6  3�      C  , , ��  3� ��  4{ �H  4{ �H  3� ��  3�      C  , , �  3� �  4{ ��  4{ ��  3� �  3�      C  , , �n  3� �n  4{ �  4{ �  3� �n  3�      C  , , �6  /{ �6  0% ��  0% ��  /{ �6  /{      C  , , ��  2_ ��  3	 �H  3	 �H  2_ ��  2_      C  , , �  2_ �  3	 ��  3	 ��  2_ �  2_      C  , , ��  2_ ��  3	 �p  3	 �p  2_ ��  2_      C  , , �.  2_ �.  3	 ��  3	 ��  2_ �.  2_      C  , , ��  2_ ��  3	 �@  3	 �@  2_ ��  2_      C  , , �^  0� �^  1� �  1� �  0� �^  0�      C  , , ��  0� ��  1� �p  1� �p  0� ��  0�      C  , , �.  0� �.  1� ��  1� ��  0� �.  0�      C  , , ��  0� ��  1� ��  1� ��  0� ��  0�      C  , , �f  0� �f  1� �  1� �  0� �f  0�      C  , , ��  0� ��  1� �x  1� �x  0� ��  0�      C  , , �f  .	 �f  .� �  .� �  .	 �f  .	      C  , , ��  .	 ��  .� �x  .� �x  .	 ��  .	      C  , , ��  .	 ��  .� �p  .� �p  .	 ��  .	      C  , , �.  .	 �.  .� ��  .� ��  .	 �.  .	      C  , , �^  3� �^  4{ �  4{ �  3� �^  3�      C  , , ��  3� ��  4{ �p  4{ �p  3� ��  3�      C  , , �.  3� �.  4{ ��  4{ ��  3� �.  3�      C  , , ��  3� ��  4{ �@  4{ �@  3� ��  3�      C  , , ��  3� ��  4{ ��  4{ ��  3� ��  3�      C  , , �f  3� �f  4{ �  4{ �  3� �f  3�      C  , , ��  3� ��  4{ �x  4{ �x  3� ��  3�      C  , , ��  .	 ��  .� �@  .� �@  .	 ��  .	      C  , , ��  2_ ��  3	 �x  3	 �x  2_ ��  2_      C  , , �f  2_ �f  3	 �  3	 �  2_ �f  2_      C  , , ��  2_ ��  3	 ��  3	 ��  2_ ��  2_      C  , , ��  0� ��  1� �@  1� �@  0� ��  0�      C  , , �^  /{ �^  0% �  0% �  /{ �^  /{      C  , , ��  /{ ��  0% �p  0% �p  /{ ��  /{      C  , , �.  /{ �.  0% ��  0% ��  /{ �.  /{      C  , , ��  /{ ��  0% �@  0% �@  /{ ��  /{      C  , , ��  /{ ��  0% ��  0% ��  /{ ��  /{      C  , , �f  /{ �f  0% �  0% �  /{ �f  /{      C  , , ��  /{ ��  0% �x  0% �x  /{ ��  /{      C  , , �^  .	 �^  .� �  .� �  .	 �^  .	      C  , , ��  .	 ��  .� ��  .� ��  .	 ��  .	      C  , , �^  2_ �^  3	 �  3	 �  2_ �^  2_      C  , , ��  &� ��  'y �x  'y �x  &� ��  &�      C  , , ��  &� ��  'y �@  'y �@  &� ��  &�      C  , , ��  &� ��  'y ��  'y ��  &� ��  &�      C  , , �.  )� �.  *] ��  *] ��  )� �.  )�      C  , , �^  (A �^  (� �  (� �  (A �^  (A      C  , , ��  (A ��  (� �p  (� �p  (A ��  (A      C  , , �.  (A �.  (� ��  (� ��  (A �.  (A      C  , , ��  (A ��  (� �@  (� �@  (A ��  (A      C  , , ��  (A ��  (� ��  (� ��  (A ��  (A      C  , , �f  (A �f  (� �  (� �  (A �f  (A      C  , , ��  )� ��  *] �@  *] �@  )� ��  )�      C  , , ��  )� ��  *] ��  *] ��  )� ��  )�      C  , , �f  )� �f  *] �  *] �  )� �f  )�      C  , , ��  )� ��  *] �x  *] �x  )� ��  )�      C  , , �f  &� �f  'y �  'y �  &� �f  &�      C  , , �^  )� �^  *] �  *] �  )� �^  )�      C  , , ��  )� ��  *] �p  *] �p  )� ��  )�      C  , , ��  (A ��  (� �x  (� �x  (A ��  (A      C  , , �^  +% �^  +� �  +� �  +% �^  +%      C  , , ��  +% ��  +� �p  +� �p  +% ��  +%      C  , , �.  +% �.  +� ��  +� ��  +% �.  +%      C  , , ��  +% ��  +� ��  +� ��  +% ��  +%      C  , , �f  +% �f  +� �  +� �  +% �f  +%      C  , , ��  +% ��  +� �x  +� �x  +% ��  +%      C  , , ��  +% ��  +� �@  +� �@  +% ��  +%      C  , , �^  &� �^  'y �  'y �  &� �^  &�      C  , , ��  &� ��  'y �p  'y �p  &� ��  &�      C  , , �.  &� �.  'y ��  'y ��  &� �.  &�      C  , , �6  (A �6  (� ��  (� ��  (A �6  (A      C  , , ��  (A ��  (� �H  (� �H  (A ��  (A      C  , , �  (A �  (� ��  (� ��  (A �  (A      C  , , �n  (A �n  (� �  (� �  (A �n  (A      C  , , �6  )� �6  *] ��  *] ��  )� �6  )�      C  , , ��  )� ��  *] �H  *] �H  )� ��  )�      C  , , �  )� �  *] ��  *] ��  )� �  )�      C  , , �  &� �  'y ��  'y ��  &� �  &�      C  , , �6  +% �6  +� ��  +� ��  +% �6  +%      C  , , ��  +% ��  +� �H  +� �H  +% ��  +%      C  , , �  +% �  +� ��  +� ��  +% �  +%      C  , , �n  +% �n  +� �  +� �  +% �n  +%      C  , , �n  &� �n  'y �  'y �  &� �n  &�      C  , , �n  )� �n  *] �  *] �  )� �n  )�      C  , , �6  &� �6  'y ��  'y ��  &� �6  &�      C  , , ��  &� ��  'y �H  'y �H  &� ��  &�      C  , , �^  # �^  � �  � �  # �^  #      C  , , ��  # ��  � �p  � �p  # ��  #      C  , , �.  # �.  � ��  � ��  # �.  #      C  , , ��  # ��  � �@  � �@  # ��  #      C  , , ��  # ��  � ��  � ��  # ��  #      C  , , �f  # �f  � �  � �  # �f  #      C  , , ��  # ��  � �x  � �x  # ��  #      C  , , �6  # �6  � ��  � ��  # �6  #      C  , , ��  # ��  � �H  � �H  # ��  #      C  , , �  # �  � ��  � ��  # �  #      C  , , �n  # �n  � �  � �  # �n  #      C  , , �2  � �2  O ��  O ��  � �2  �      C  , , ��  � ��  O �*  O �*  � ��  �      C  , , �n  � �n   ? �   ? �  � �n  �      C  , , �  � �   ? ��   ? ��  � �  �      C  , , �2    �2   � ��   � ��    �2         C  , , ��    ��   � �*   � �*    ��         C  , , �n  ! �n  !� �  !� �  ! �n  !      C  , , �2  !u �2  " ��  " ��  !u �2  !u      C  , , ��  !u ��  " �*  " �*  !u ��  !u      C  , , ��  "� ��  #� �*  #� �*  "� ��  "�      C  , , �6  #� �6  $� ��  $� ��  #� �6  #�      C  , , ��  #� ��  $� �H  $� �H  #� ��  #�      C  , , �6  ! �6  !� ��  !� ��  ! �6  !      C  , , ��  ! ��  !� �H  !� �H  ! ��  !      C  , , �  ! �  !� ��  !� ��  ! �  !      C  , , �  #� �  $� ��  $� ��  #� �  #�      C  , , �n  #� �n  $� �  $� �  #� �n  #�      C  , , �6  � �6   ? ��   ? ��  � �6  �      C  , , ��  � ��   ? �H   ? �H  � ��  �      C  , , �6  "y �6  ## ��  ## ��  "y �6  "y      C  , , ��  "y ��  ## �H  ## �H  "y ��  "y      C  , , �  "y �  ## ��  ## ��  "y �  "y      C  , , �n  "y �n  ## �  ## �  "y �n  "y      C  , , �2  "� �2  #� ��  #� ��  "� �2  "�      C  , , �f  ! �f  !� �  !� �  ! �f  !      C  , , ��  ! ��  !� �x  !� �x  ! ��  !      C  , , �.  ! �.  !� ��  !� ��  ! �.  !      C  , , ��  ! ��  !� �@  !� �@  ! ��  !      C  , , �^  #� �^  $� �  $� �  #� �^  #�      C  , , �^  � �^   ? �   ? �  � �^  �      C  , , ��  � ��   ? �p   ? �p  � ��  �      C  , , �.  � �.   ? ��   ? ��  � �.  �      C  , , ��  � ��   ? �@   ? �@  � ��  �      C  , , ��  #� ��  $� �p  $� �p  #� ��  #�      C  , , �.  #� �.  $� ��  $� ��  #� �.  #�      C  , , ��  � ��   ? ��   ? ��  � ��  �      C  , , �f  � �f   ? �   ? �  � �f  �      C  , , ��  � ��   ? �x   ? �x  � ��  �      C  , , ��  #� ��  $� �@  $� �@  #� ��  #�      C  , , ��  #� ��  $� ��  $� ��  #� ��  #�      C  , , �^  "y �^  ## �  ## �  "y �^  "y      C  , , ��  "y ��  ## �p  ## �p  "y ��  "y      C  , , �.  "y �.  ## ��  ## ��  "y �.  "y      C  , , ��  "y ��  ## �@  ## �@  "y ��  "y      C  , , ��  "y ��  ## ��  ## ��  "y ��  "y      C  , , �f  "y �f  ## �  ## �  "y �f  "y      C  , , ��  "y ��  ## �x  ## �x  "y ��  "y      C  , , �f  #� �f  $� �  $� �  #� �f  #�      C  , , ��  #� ��  $� �x  $� �x  #� ��  #�      C  , , �^  ! �^  !� �  !� �  ! �^  !      C  , , ��  ! ��  !� �p  !� �p  ! ��  !      C  , , ��  ! ��  !� ��  !� ��  ! ��  !      C  , , ��  ? ��  � �p  � �p  ? ��  ?      C  , , �^  � �^  w �  w �  � �^  �      C  , , ��  � ��  w �p  w �p  � ��  �      C  , , �.  � �.  w ��  w ��  � �.  �      C  , , ��  � ��  w �@  w �@  � ��  �      C  , , ��  � ��  w ��  w ��  � ��  �      C  , , �f  � �f  w �  w �  � �f  �      C  , , ��  � ��  w �x  w �x  � ��  �      C  , , ��  � ��  [ �x  [ �x  � ��  �      C  , , �^  [ �^   �   �  [ �^  [      C  , , �^  � �^  [ �  [ �  � �^  �      C  , , ��  � ��  [ �p  [ �p  � ��  �      C  , , �.  � �.  [ ��  [ ��  � �.  �      C  , , ��  � ��  [ �@  [ �@  � ��  �      C  , , ��  � ��  [ ��  [ ��  � ��  �      C  , , �f  � �f  [ �  [ �  � �f  �      C  , , �.  ? �.  � ��  � ��  ? �.  ?      C  , , ��  ? ��  � �@  � �@  ? ��  ?      C  , , ��  ? ��  � ��  � ��  ? ��  ?      C  , , �f  ? �f  � �  � �  ? �f  ?      C  , , ��  ? ��  � �x  � �x  ? ��  ?      C  , , ��  [ ��   �p   �p  [ ��  [      C  , , �.  [ �.   ��   ��  [ �.  [      C  , , ��  [ ��   �@   �@  [ ��  [      C  , , ��  [ ��   ��   ��  [ ��  [      C  , , �f  [ �f   �   �  [ �f  [      C  , , ��  [ ��   �x   �x  [ ��  [      C  , , �^  ? �^  � �  � �  ? �^  ?      C  , , �  � �  [ ��  [ ��  � �  �      C  , , �6  � �6  [ ��  [ ��  � �6  �      C  , , �6  � �6  w ��  w ��  � �6  �      C  , , ��  � ��  w �H  w �H  � ��  �      C  , , �  � �  w ��  w ��  � �  �      C  , , �6  [ �6   ��   ��  [ �6  [      C  , , ��  [ ��   �H   �H  [ ��  [      C  , , �6  ? �6  � ��  � ��  ? �6  ?      C  , , ��  ? ��  � �H  � �H  ? ��  ?      C  , , �  ? �  � ��  � ��  ? �  ?      C  , , �n  ? �n  � �  � �  ? �n  ?      C  , , �2  � �2   ��   ��  � �2  �      C  , , ��  � ��   �*   �*  � ��  �      C  , , �  [ �   ��   ��  [ �  [      C  , , �n  [ �n   �   �  [ �n  [      C  , , �n  � �n  w �  w �  � �n  �      C  , , �2  m �2   ��   ��  m �2  m      C  , , ��  m ��   �*   �*  m ��  m      C  , , �n  � �n  [ �  [ �  � �n  �      C  , , �2  = �2  � ��  � ��  = �2  =      C  , , �2   �2  � ��  � ��   �2        C  , , ��   ��  � �*  � �*   ��        C  , , ��  = ��  � �*  � �*  = ��  =      C  , , ��  � ��  [ �H  [ �H  � ��  �      C  , , �   �  � ��  � ��   �        C  , , �j   �j  � �  � �   �j        C  , , ��   ��  � �b  � �b   ��        C  , , �   �  � ��  � ��   �        C  , , �T   �T  � ��  � ��   �T        C  , , ��   ��  � �L  � �L   ��        C  , , ��   ��  � ��  � ��   ��        C  , , �>   �>  � ��  � ��   �>        C  , , ��   ��  � �6  � �6   ��        C  , , �  � �   ��   ��  � �  �      C  , , �T  � �T   ��   ��  � �T  �      C  , , ��  � ��   �L   �L  � ��  �      C  , , ��  � ��   ��   ��  � ��  �      C  , , �>  � �>   ��   ��  � �>  �      C  , , ��  � ��   �6   �6  � ��  �      C  , , ��  � ��  O �L  O �L  � ��  �      C  , , ��  � ��  O ��  O ��  � ��  �      C  , , ��  = ��  � �x  � �x  = ��  =      C  , , �  = �  � ��  � ��  = �  =      C  , , �j  = �j  � �  � �  = �j  =      C  , , ��  = ��  � �b  � �b  = ��  =      C  , , �  = �  � ��  � ��  = �  =      C  , , �T  = �T  � ��  � ��  = �T  =      C  , , ��  = ��  � �L  � �L  = ��  =      C  , , ��  = ��  � ��  � ��  = ��  =      C  , , �>  = �>  � ��  � ��  = �>  =      C  , , ��  = ��  � �6  � �6  = ��  =      C  , , �>  � �>  O ��  O ��  � �>  �      C  , , ��  � ��  O �6  O �6  � ��  �      C  , , �  "� �  #� ��  #� ��  "� �  "�      C  , , �T  "� �T  #� ��  #� ��  "� �T  "�      C  , , ��  "� ��  #� �L  #� �L  "� ��  "�      C  , , ��  "� ��  #� ��  #� ��  "� ��  "�      C  , , ��  !u ��  " �x  " �x  !u ��  !u      C  , , �  !u �  " ��  " ��  !u �  !u      C  , , �j  !u �j  " �  " �  !u �j  !u      C  , , ��  !u ��  " �b  " �b  !u ��  !u      C  , , �  !u �  " ��  " ��  !u �  !u      C  , , �T  !u �T  " ��  " ��  !u �T  !u      C  , , ��  !u ��  " �L  " �L  !u ��  !u      C  , , ��  !u ��  " ��  " ��  !u ��  !u      C  , , ��    ��   � �x   � �x    ��         C  , , �    �   � ��   � ��    �         C  , , �j    �j   � �   � �    �j         C  , , ��    ��   � �b   � �b    ��         C  , , �    �   � ��   � ��    �         C  , , �T    �T   � ��   � ��    �T         C  , , ��    ��   � �L   � �L    ��         C  , , ��    ��   � ��   � ��    ��         C  , , �>    �>   � ��   � ��    �>         C  , , ��    ��   � �6   � �6    ��         C  , , �>  !u �>  " ��  " ��  !u �>  !u      C  , , ��  !u ��  " �6  " �6  !u ��  !u      C  , , ��  m ��   �x   �x  m ��  m      C  , , �  m �   ��   ��  m �  m      C  , , �j  m �j   �   �  m �j  m      C  , , ��  m ��   �b   �b  m ��  m      C  , , �  m �   ��   ��  m �  m      C  , , �T  m �T   ��   ��  m �T  m      C  , , ��  m ��   �L   �L  m ��  m      C  , , ��  m ��   ��   ��  m ��  m      C  , , �>  m �>   ��   ��  m �>  m      C  , , ��  m ��   �6   �6  m ��  m      C  , , �>  "� �>  #� ��  #� ��  "� �>  "�      C  , , ��  "� ��  #� �6  #� �6  "� ��  "�      C  , , ��  "� ��  #� �x  #� �x  "� ��  "�      C  , , �  "� �  #� ��  #� ��  "� �  "�      C  , , �j  "� �j  #� �  #� �  "� �j  "�      C  , , ��  "� ��  #� �b  #� �b  "� ��  "�      C  , , ��  % ��  %� �Q  %� �Q  % ��  %      C  , , ��  % ��  %� ��  %� ��  % ��  %      C  , , �C  % �C  %� ��  %� ��  % �C  %      C  , , ��  % ��  %� �;  %� �;  % ��  %      C  , , ��  % ��  %� ��  %� ��  % ��  %      C  , , �-  % �-  %� ��  %� ��  % �-  %      C  , , �{  % �{  %� �%  %� �%  % �{  %      C  , , ��  % ��  %� �s  %� �s  % ��  %      C  , , �  % �  %� ��  %� ��  % �  %      C  , , �e  % �e  %� �  %� �  % �e  %      C  , , ��  % ��  %� �]  %� �]  % ��  %      C  , , ��  � ��  O �x  O �x  � ��  �      C  , , �  � �  O ��  O ��  � �  �      C  , , �j  � �j  O �  O �  � �j  �      C  , , ��  � ��  O �b  O �b  � ��  �      C  , , �  � �  O ��  O ��  � �  �      C  , , �T  � �T  O ��  O ��  � �T  �      C  , , ��  � ��   �x   �x  � ��  �      C  , , �  � �   ��   ��  � �  �      C  , , �j  � �j   �   �  � �j  �      C  , , ��  � ��   �b   �b  � ��  �      C  , , ��   ��  � �x  � �x   ��        C  , , g=  "� g=  #� g�  #� g�  "� g=  "�      C  , , g=  *� g=  +k g�  +k g�  *� g=  *�      C  , , g=  0a g=  1 g�  1 g�  0a g=  0a      C  , , g=  !u g=  " g�  " g�  !u g=  !u      C  , , g=    g=   � g�   � g�    g=         C  , , g=  )Y g=  * g�  * g�  )Y g=  )Y      C  , , g=  -� g=  .; g�  .; g�  -� g=  -�      C  , , g=  � g=  O g�  O g�  � g=  �      C  , , g=  1� g=  2s g�  2s g�  1� g=  1�      C  , , g=  = g=  � g�  � g�  = g=  =      C  , , g=  � g=   g�   g�  � g=  �      C  , , g=  ,) g=  ,� g�  ,� g�  ,) g=  ,)      C  , , g=  m g=   g�   g�  m g=  m      C  , , g=   g=  � g�  � g�   g=        C  , , g=  .� g=  /� g�  /� g�  .� g=  .�      C  , , g=  31 g=  3� g�  3� g�  31 g=  31      C  , , k�  *� k�  +k l�  +k l�  *� k�  *�      C  , , pu  0a pu  1 q  1 q  0a pu  0a      C  , , r�  0a r�  1 sm  1 sm  0a r�  0a      C  , , u  0a u  1 u�  1 u�  0a u  0a      C  , , w_  0a w_  1 x	  1 x	  0a w_  0a      C  , , y�  0a y�  1 zW  1 zW  0a y�  0a      C  , , {�  0a {�  1 |�  1 |�  0a {�  0a      C  , , ~I  0a ~I  1 ~�  1 ~�  0a ~I  0a      C  , , n'  *� n'  +k n�  +k n�  *� n'  *�      C  , , pu  *� pu  +k q  +k q  *� pu  *�      C  , , i�  )Y i�  * j5  * j5  )Y i�  )Y      C  , , k�  )Y k�  * l�  * l�  )Y k�  )Y      C  , , n'  )Y n'  * n�  * n�  )Y n'  )Y      C  , , pu  )Y pu  * q  * q  )Y pu  )Y      C  , , r�  )Y r�  * sm  * sm  )Y r�  )Y      C  , , u  )Y u  * u�  * u�  )Y u  )Y      C  , , w_  )Y w_  * x	  * x	  )Y w_  )Y      C  , , y�  )Y y�  * zW  * zW  )Y y�  )Y      C  , , {�  )Y {�  * |�  * |�  )Y {�  )Y      C  , , ~I  )Y ~I  * ~�  * ~�  )Y ~I  )Y      C  , , r�  *� r�  +k sm  +k sm  *� r�  *�      C  , , i�  -� i�  .; j5  .; j5  -� i�  -�      C  , , k�  -� k�  .; l�  .; l�  -� k�  -�      C  , , n'  -� n'  .; n�  .; n�  -� n'  -�      C  , , pu  -� pu  .; q  .; q  -� pu  -�      C  , , r�  -� r�  .; sm  .; sm  -� r�  -�      C  , , u  *� u  +k u�  +k u�  *� u  *�      C  , , u  -� u  .; u�  .; u�  -� u  -�      C  , , w_  -� w_  .; x	  .; x	  -� w_  -�      C  , , y�  -� y�  .; zW  .; zW  -� y�  -�      C  , , {�  -� {�  .; |�  .; |�  -� {�  -�      C  , , ~I  -� ~I  .; ~�  .; ~�  -� ~I  -�      C  , , w_  *� w_  +k x	  +k x	  *� w_  *�      C  , , i�  1� i�  2s j5  2s j5  1� i�  1�      C  , , k�  1� k�  2s l�  2s l�  1� k�  1�      C  , , n'  1� n'  2s n�  2s n�  1� n'  1�      C  , , pu  1� pu  2s q  2s q  1� pu  1�      C  , , r�  1� r�  2s sm  2s sm  1� r�  1�      C  , , u  1� u  2s u�  2s u�  1� u  1�      C  , , w_  1� w_  2s x	  2s x	  1� w_  1�      C  , , y�  1� y�  2s zW  2s zW  1� y�  1�      C  , , {�  1� {�  2s |�  2s |�  1� {�  1�      C  , , ~I  1� ~I  2s ~�  2s ~�  1� ~I  1�      C  , , y�  *� y�  +k zW  +k zW  *� y�  *�      C  , , hd  ') hd  '� i  '� i  ') hd  ')      C  , , j�  ') j�  '� k\  '� k\  ') j�  ')      C  , , m   ') m   '� m�  '� m�  ') m   ')      C  , , oN  ') oN  '� o�  '� o�  ') oN  ')      C  , , q�  ') q�  '� rF  '� rF  ') q�  ')      C  , , s�  ') s�  '� t�  '� t�  ') s�  ')      C  , , v8  ') v8  '� v�  '� v�  ') v8  ')      C  , , x�  ') x�  '� y0  '� y0  ') x�  ')      C  , , z�  ') z�  '� {~  '� {~  ') z�  ')      C  , , }"  ') }"  '� }�  '� }�  ') }"  ')      C  , , {�  *� {�  +k |�  +k |�  *� {�  *�      C  , , ~I  *� ~I  +k ~�  +k ~�  *� ~I  *�      C  , , i�  ,) i�  ,� j5  ,� j5  ,) i�  ,)      C  , , k�  ,) k�  ,� l�  ,� l�  ,) k�  ,)      C  , , n'  ,) n'  ,� n�  ,� n�  ,) n'  ,)      C  , , i�  *� i�  +k j5  +k j5  *� i�  *�      C  , , pu  ,) pu  ,� q  ,� q  ,) pu  ,)      C  , , r�  ,) r�  ,� sm  ,� sm  ,) r�  ,)      C  , , u  ,) u  ,� u�  ,� u�  ,) u  ,)      C  , , w_  ,) w_  ,� x	  ,� x	  ,) w_  ,)      C  , , y�  ,) y�  ,� zW  ,� zW  ,) y�  ,)      C  , , {�  ,) {�  ,� |�  ,� |�  ,) {�  ,)      C  , , ~I  ,) ~I  ,� ~�  ,� ~�  ,) ~I  ,)      C  , , i�  0a i�  1 j5  1 j5  0a i�  0a      C  , , k�  0a k�  1 l�  1 l�  0a k�  0a      C  , , i�  .� i�  /� j5  /� j5  .� i�  .�      C  , , k�  .� k�  /� l�  /� l�  .� k�  .�      C  , , n'  .� n'  /� n�  /� n�  .� n'  .�      C  , , pu  .� pu  /� q  /� q  .� pu  .�      C  , , r�  .� r�  /� sm  /� sm  .� r�  .�      C  , , u  .� u  /� u�  /� u�  .� u  .�      C  , , w_  .� w_  /� x	  /� x	  .� w_  .�      C  , , y�  .� y�  /� zW  /� zW  .� y�  .�      C  , , {�  .� {�  /� |�  /� |�  .� {�  .�      C  , , ~I  .� ~I  /� ~�  /� ~�  .� ~I  .�      C  , , n'  0a n'  1 n�  1 n�  0a n'  0a      C  , , i�  31 i�  3� j5  3� j5  31 i�  31      C  , , k�  31 k�  3� l�  3� l�  31 k�  31      C  , , n'  31 n'  3� n�  3� n�  31 n'  31      C  , , pu  31 pu  3� q  3� q  31 pu  31      C  , , r�  31 r�  3� sm  3� sm  31 r�  31      C  , , u  31 u  3� u�  3� u�  31 u  31      C  , , w_  31 w_  3� x	  3� x	  31 w_  31      C  , , y�  31 y�  3� zW  3� zW  31 y�  31      C  , , {�  31 {�  3� |�  3� |�  31 {�  31      C  , , ~I  31 ~I  3� ~�  3� ~�  31 ~I  31      C  , , Yi  0a Yi  1 Z  1 Z  0a Yi  0a      C  , , [�  0a [�  1 \a  1 \a  0a [�  0a      C  , , ^  0a ^  1 ^�  1 ^�  0a ^  0a      C  , , `S  0a `S  1 `�  1 `�  0a `S  0a      C  , , O
  ') O
  '� O�  '� O�  ') O
  ')      C  , , QX  ') QX  '� R  '� R  ') QX  ')      C  , , S�  ') S�  '� TP  '� TP  ') S�  ')      C  , , U�  ') U�  '� V�  '� V�  ') U�  ')      C  , , XB  ') XB  '� X�  '� X�  ') XB  ')      C  , , Z�  ') Z�  '� [:  '� [:  ') Z�  ')      C  , , \�  ') \�  '� ]�  '� ]�  ') \�  ')      C  , , _,  ') _,  '� _�  '� _�  ') _,  ')      C  , , az  ') az  '� b$  '� b$  ') az  ')      C  , , c�  ') c�  '� dr  '� dr  ') c�  ')      C  , , f  ') f  '� f�  '� f�  ') f  ')      C  , , b�  0a b�  1 cK  1 cK  0a b�  0a      C  , , d�  0a d�  1 e�  1 e�  0a d�  0a      C  , , R  *� R  +k S)  +k S)  *� R  *�      C  , , T�  *� T�  +k Uw  +k Uw  *� T�  *�      C  , , W  *� W  +k W�  +k W�  *� W  *�      C  , , Yi  *� Yi  +k Z  +k Z  *� Yi  *�      C  , , P1  -� P1  .; P�  .; P�  -� P1  -�      C  , , R  -� R  .; S)  .; S)  -� R  -�      C  , , T�  -� T�  .; Uw  .; Uw  -� T�  -�      C  , , W  -� W  .; W�  .; W�  -� W  -�      C  , , Yi  -� Yi  .; Z  .; Z  -� Yi  -�      C  , , P1  ,) P1  ,� P�  ,� P�  ,) P1  ,)      C  , , R  ,) R  ,� S)  ,� S)  ,) R  ,)      C  , , T�  ,) T�  ,� Uw  ,� Uw  ,) T�  ,)      C  , , W  ,) W  ,� W�  ,� W�  ,) W  ,)      C  , , Yi  ,) Yi  ,� Z  ,� Z  ,) Yi  ,)      C  , , [�  ,) [�  ,� \a  ,� \a  ,) [�  ,)      C  , , ^  ,) ^  ,� ^�  ,� ^�  ,) ^  ,)      C  , , `S  ,) `S  ,� `�  ,� `�  ,) `S  ,)      C  , , b�  ,) b�  ,� cK  ,� cK  ,) b�  ,)      C  , , d�  ,) d�  ,� e�  ,� e�  ,) d�  ,)      C  , , [�  -� [�  .; \a  .; \a  -� [�  -�      C  , , ^  -� ^  .; ^�  .; ^�  -� ^  -�      C  , , `S  -� `S  .; `�  .; `�  -� `S  -�      C  , , b�  -� b�  .; cK  .; cK  -� b�  -�      C  , , d�  -� d�  .; e�  .; e�  -� d�  -�      C  , , [�  *� [�  +k \a  +k \a  *� [�  *�      C  , , ^  *� ^  +k ^�  +k ^�  *� ^  *�      C  , , `S  *� `S  +k `�  +k `�  *� `S  *�      C  , , b�  *� b�  +k cK  +k cK  *� b�  *�      C  , , d�  *� d�  +k e�  +k e�  *� d�  *�      C  , , P1  *� P1  +k P�  +k P�  *� P1  *�      C  , , P1  0a P1  1 P�  1 P�  0a P1  0a      C  , , R  0a R  1 S)  1 S)  0a R  0a      C  , , P1  .� P1  /� P�  /� P�  .� P1  .�      C  , , R  .� R  /� S)  /� S)  .� R  .�      C  , , T�  .� T�  /� Uw  /� Uw  .� T�  .�      C  , , W  .� W  /� W�  /� W�  .� W  .�      C  , , Yi  .� Yi  /� Z  /� Z  .� Yi  .�      C  , , [�  .� [�  /� \a  /� \a  .� [�  .�      C  , , ^  .� ^  /� ^�  /� ^�  .� ^  .�      C  , , `S  .� `S  /� `�  /� `�  .� `S  .�      C  , , b�  .� b�  /� cK  /� cK  .� b�  .�      C  , , d�  .� d�  /� e�  /� e�  .� d�  .�      C  , , T�  0a T�  1 Uw  1 Uw  0a T�  0a      C  , , P1  )Y P1  * P�  * P�  )Y P1  )Y      C  , , R  )Y R  * S)  * S)  )Y R  )Y      C  , , T�  )Y T�  * Uw  * Uw  )Y T�  )Y      C  , , P1  1� P1  2s P�  2s P�  1� P1  1�      C  , , R  1� R  2s S)  2s S)  1� R  1�      C  , , T�  1� T�  2s Uw  2s Uw  1� T�  1�      C  , , W  1� W  2s W�  2s W�  1� W  1�      C  , , Yi  1� Yi  2s Z  2s Z  1� Yi  1�      C  , , [�  1� [�  2s \a  2s \a  1� [�  1�      C  , , ^  1� ^  2s ^�  2s ^�  1� ^  1�      C  , , P1  31 P1  3� P�  3� P�  31 P1  31      C  , , R  31 R  3� S)  3� S)  31 R  31      C  , , T�  31 T�  3� Uw  3� Uw  31 T�  31      C  , , W  31 W  3� W�  3� W�  31 W  31      C  , , Yi  31 Yi  3� Z  3� Z  31 Yi  31      C  , , [�  31 [�  3� \a  3� \a  31 [�  31      C  , , ^  31 ^  3� ^�  3� ^�  31 ^  31      C  , , `S  31 `S  3� `�  3� `�  31 `S  31      C  , , b�  31 b�  3� cK  3� cK  31 b�  31      C  , , d�  31 d�  3� e�  3� e�  31 d�  31      C  , , `S  1� `S  2s `�  2s `�  1� `S  1�      C  , , b�  1� b�  2s cK  2s cK  1� b�  1�      C  , , d�  1� d�  2s e�  2s e�  1� d�  1�      C  , , W  )Y W  * W�  * W�  )Y W  )Y      C  , , Yi  )Y Yi  * Z  * Z  )Y Yi  )Y      C  , , [�  )Y [�  * \a  * \a  )Y [�  )Y      C  , , ^  )Y ^  * ^�  * ^�  )Y ^  )Y      C  , , `S  )Y `S  * `�  * `�  )Y `S  )Y      C  , , b�  )Y b�  * cK  * cK  )Y b�  )Y      C  , , d�  )Y d�  * e�  * e�  )Y d�  )Y      C  , , W  0a W  1 W�  1 W�  0a W  0a      C  , , `S    `S   � `�   � `�    `S         C  , , b�    b�   � cK   � cK    b�         C  , , d�    d�   � e�   � e�    d�         C  , , d�  "� d�  #� e�  #� e�  "� d�  "�      C  , , P1  !u P1  " P�  " P�  !u P1  !u      C  , , R  !u R  " S)  " S)  !u R  !u      C  , , T�  !u T�  " Uw  " Uw  !u T�  !u      C  , , W  !u W  " W�  " W�  !u W  !u      C  , , P1  m P1   P�   P�  m P1  m      C  , , R  m R   S)   S)  m R  m      C  , , T�  m T�   Uw   Uw  m T�  m      C  , , W  m W   W�   W�  m W  m      C  , , Yi  m Yi   Z   Z  m Yi  m      C  , , [�  m [�   \a   \a  m [�  m      C  , , ^  m ^   ^�   ^�  m ^  m      C  , , `S  m `S   `�   `�  m `S  m      C  , , b�  m b�   cK   cK  m b�  m      C  , , d�  m d�   e�   e�  m d�  m      C  , , Yi  !u Yi  " Z  " Z  !u Yi  !u      C  , , O
  % O
  %� O�  %� O�  % O
  %      C  , , QX  % QX  %� R  %� R  % QX  %      C  , , S�  % S�  %� TP  %� TP  % S�  %      C  , , U�  % U�  %� V�  %� V�  % U�  %      C  , , XB  % XB  %� X�  %� X�  % XB  %      C  , , Z�  % Z�  %� [:  %� [:  % Z�  %      C  , , \�  % \�  %� ]�  %� ]�  % \�  %      C  , , _,  % _,  %� _�  %� _�  % _,  %      C  , , az  % az  %� b$  %� b$  % az  %      C  , , c�  % c�  %� dr  %� dr  % c�  %      C  , , f  % f  %� f�  %� f�  % f  %      C  , , [�  !u [�  " \a  " \a  !u [�  !u      C  , , P1  = P1  � P�  � P�  = P1  =      C  , , R  = R  � S)  � S)  = R  =      C  , , T�  = T�  � Uw  � Uw  = T�  =      C  , , W  = W  � W�  � W�  = W  =      C  , , Yi  = Yi  � Z  � Z  = Yi  =      C  , , [�  = [�  � \a  � \a  = [�  =      C  , , P1   P1  � P�  � P�   P1        C  , , R   R  � S)  � S)   R        C  , , T�   T�  � Uw  � Uw   T�        C  , , W   W  � W�  � W�   W        C  , , Yi   Yi  � Z  � Z   Yi        C  , , [�   [�  � \a  � \a   [�        C  , , ^   ^  � ^�  � ^�   ^        C  , , `S   `S  � `�  � `�   `S        C  , , b�   b�  � cK  � cK   b�        C  , , d�   d�  � e�  � e�   d�        C  , , ^  = ^  � ^�  � ^�  = ^  =      C  , , `S  = `S  � `�  � `�  = `S  =      C  , , b�  = b�  � cK  � cK  = b�  =      C  , , d�  = d�  � e�  � e�  = d�  =      C  , , ^  !u ^  " ^�  " ^�  !u ^  !u      C  , , `S  !u `S  " `�  " `�  !u `S  !u      C  , , P1  � P1  O P�  O P�  � P1  �      C  , , R  � R  O S)  O S)  � R  �      C  , , T�  � T�  O Uw  O Uw  � T�  �      C  , , W  � W  O W�  O W�  � W  �      C  , , Yi  � Yi  O Z  O Z  � Yi  �      C  , , [�  � [�  O \a  O \a  � [�  �      C  , , ^  � ^  O ^�  O ^�  � ^  �      C  , , `S  � `S  O `�  O `�  � `S  �      C  , , b�  � b�  O cK  O cK  � b�  �      C  , , d�  � d�  O e�  O e�  � d�  �      C  , , b�  !u b�  " cK  " cK  !u b�  !u      C  , , d�  !u d�  " e�  " e�  !u d�  !u      C  , , R  "� R  #� S)  #� S)  "� R  "�      C  , , T�  "� T�  #� Uw  #� Uw  "� T�  "�      C  , , W  "� W  #� W�  #� W�  "� W  "�      C  , , Yi  "� Yi  #� Z  #� Z  "� Yi  "�      C  , , [�  "� [�  #� \a  #� \a  "� [�  "�      C  , , ^  "� ^  #� ^�  #� ^�  "� ^  "�      C  , , `S  "� `S  #� `�  #� `�  "� `S  "�      C  , , b�  "� b�  #� cK  #� cK  "� b�  "�      C  , , P1  � P1   P�   P�  � P1  �      C  , , R  � R   S)   S)  � R  �      C  , , T�  � T�   Uw   Uw  � T�  �      C  , , W  � W   W�   W�  � W  �      C  , , Yi  � Yi   Z   Z  � Yi  �      C  , , [�  � [�   \a   \a  � [�  �      C  , , ^  � ^   ^�   ^�  � ^  �      C  , , `S  � `S   `�   `�  � `S  �      C  , , b�  � b�   cK   cK  � b�  �      C  , , d�  � d�   e�   e�  � d�  �      C  , , P1    P1   � P�   � P�    P1         C  , , R    R   � S)   � S)    R         C  , , T�    T�   � Uw   � Uw    T�         C  , , W    W   � W�   � W�    W         C  , , Yi    Yi   � Z   � Z    Yi         C  , , [�    [�   � \a   � \a    [�         C  , , ^    ^   � ^�   � ^�    ^         C  , , P1  "� P1  #� P�  #� P�  "� P1  "�      C  , , r�    r�   � sm   � sm    r�         C  , , u    u   � u�   � u�    u         C  , , w_    w_   � x	   � x	    w_         C  , , y�    y�   � zW   � zW    y�         C  , , {�    {�   � |�   � |�    {�         C  , , ~I    ~I   � ~�   � ~�    ~I         C  , , {�  !u {�  " |�  " |�  !u {�  !u      C  , , ~I  !u ~I  " ~�  " ~�  !u ~I  !u      C  , , w_  "� w_  #� x	  #� x	  "� w_  "�      C  , , hd  % hd  %� i  %� i  % hd  %      C  , , j�  % j�  %� k\  %� k\  % j�  %      C  , , m   % m   %� m�  %� m�  % m   %      C  , , oN  % oN  %� o�  %� o�  % oN  %      C  , , q�  % q�  %� rF  %� rF  % q�  %      C  , , s�  % s�  %� t�  %� t�  % s�  %      C  , , v8  % v8  %� v�  %� v�  % v8  %      C  , , x�  % x�  %� y0  %� y0  % x�  %      C  , , z�  % z�  %� {~  %� {~  % z�  %      C  , , }"  % }"  %� }�  %� }�  % }"  %      C  , , y�  "� y�  #� zW  #� zW  "� y�  "�      C  , , {�  "� {�  #� |�  #� |�  "� {�  "�      C  , , ~I  "� ~I  #� ~�  #� ~�  "� ~I  "�      C  , , i�  "� i�  #� j5  #� j5  "� i�  "�      C  , , k�  "� k�  #� l�  #� l�  "� k�  "�      C  , , n'  "� n'  #� n�  #� n�  "� n'  "�      C  , , pu  "� pu  #� q  #� q  "� pu  "�      C  , , r�  "� r�  #� sm  #� sm  "� r�  "�      C  , , u  "� u  #� u�  #� u�  "� u  "�      C  , , i�  !u i�  " j5  " j5  !u i�  !u      C  , , k�  !u k�  " l�  " l�  !u k�  !u      C  , , n'  !u n'  " n�  " n�  !u n'  !u      C  , , pu  !u pu  " q  " q  !u pu  !u      C  , , r�  !u r�  " sm  " sm  !u r�  !u      C  , , i�  � i�   j5   j5  � i�  �      C  , , k�  � k�   l�   l�  � k�  �      C  , , n'  � n'   n�   n�  � n'  �      C  , , pu  � pu   q   q  � pu  �      C  , , i�   i�  � j5  � j5   i�        C  , , k�   k�  � l�  � l�   k�        C  , , n'   n'  � n�  � n�   n'        C  , , pu   pu  � q  � q   pu        C  , , r�   r�  � sm  � sm   r�        C  , , u   u  � u�  � u�   u        C  , , w_   w_  � x	  � x	   w_        C  , , y�   y�  � zW  � zW   y�        C  , , {�   {�  � |�  � |�   {�        C  , , ~I   ~I  � ~�  � ~�   ~I        C  , , r�  � r�   sm   sm  � r�  �      C  , , u  � u   u�   u�  � u  �      C  , , w_  � w_   x	   x	  � w_  �      C  , , y�  � y�   zW   zW  � y�  �      C  , , {�  � {�   |�   |�  � {�  �      C  , , ~I  � ~I   ~�   ~�  � ~I  �      C  , , u  !u u  " u�  " u�  !u u  !u      C  , , i�  � i�  O j5  O j5  � i�  �      C  , , k�  � k�  O l�  O l�  � k�  �      C  , , n'  � n'  O n�  O n�  � n'  �      C  , , pu  � pu  O q  O q  � pu  �      C  , , r�  � r�  O sm  O sm  � r�  �      C  , , u  � u  O u�  O u�  � u  �      C  , , w_  � w_  O x	  O x	  � w_  �      C  , , i�  = i�  � j5  � j5  = i�  =      C  , , k�  = k�  � l�  � l�  = k�  =      C  , , n'  = n'  � n�  � n�  = n'  =      C  , , pu  = pu  � q  � q  = pu  =      C  , , r�  = r�  � sm  � sm  = r�  =      C  , , u  = u  � u�  � u�  = u  =      C  , , w_  = w_  � x	  � x	  = w_  =      C  , , y�  = y�  � zW  � zW  = y�  =      C  , , {�  = {�  � |�  � |�  = {�  =      C  , , ~I  = ~I  � ~�  � ~�  = ~I  =      C  , , y�  � y�  O zW  O zW  � y�  �      C  , , {�  � {�  O |�  O |�  � {�  �      C  , , ~I  � ~I  O ~�  O ~�  � ~I  �      C  , , w_  !u w_  " x	  " x	  !u w_  !u      C  , , y�  !u y�  " zW  " zW  !u y�  !u      C  , , i�    i�   � j5   � j5    i�         C  , , k�    k�   � l�   � l�    k�         C  , , i�  m i�   j5   j5  m i�  m      C  , , k�  m k�   l�   l�  m k�  m      C  , , n'  m n'   n�   n�  m n'  m      C  , , pu  m pu   q   q  m pu  m      C  , , r�  m r�   sm   sm  m r�  m      C  , , u  m u   u�   u�  m u  m      C  , , w_  m w_   x	   x	  m w_  m      C  , , y�  m y�   zW   zW  m y�  m      C  , , {�  m {�   |�   |�  m {�  m      C  , , ~I  m ~I   ~�   ~�  m ~I  m      C  , , n'    n'   � n�   � n�    n'         C  , , pu    pu   � q   � q    pu         C  , , 6  &� 6  'y 6�  'y 6�  &� 6  &�      C  , , 6  ! 6  !� 6�  !� 6�  ! 6  !      C  , , 6  2_ 6  3	 6�  3	 6�  2_ 6  2_      C  , , 6  .	 6  .� 6�  .� 6�  .	 6  .	      C  , , 6  ? 6  � 6�  � 6�  ? 6  ?      C  , , 6  ,� 6  -A 6�  -A 6�  ,� 6  ,�      C  , , 6  3� 6  4{ 6�  4{ 6�  3� 6  3�      C  , , 6  � 6  w 6�  w 6�  � 6  �      C  , , 6  # 6  � 6�  � 6�  # 6  #      C  , , 1�  %] 1�  & 2�  & 2�  %] 1�  %]      C  , , 3?  %] 3?  & 3�  & 3�  %] 3?  %]      C  , , 4�  %] 4�  & 5Q  & 5Q  %] 4�  %]      C  , , 6  %] 6  & 6�  & 6�  %] 6  %]      C  , , 7w  %] 7w  & 8!  & 8!  %] 7w  %]      C  , , 8�  %] 8�  & 9�  & 9�  %] 8�  %]      C  , , :G  %] :G  & :�  & :�  %] :G  %]      C  , , ;�  %] ;�  & <Y  & <Y  %] ;�  %]      C  , , =  %] =  & =�  & =�  %] =  %]      C  , , >  %] >  & ?)  & ?)  %] >  %]      C  , , ?�  %] ?�  & @�  & @�  %] ?�  %]      C  , , 6  )� 6  *] 6�  *] 6�  )� 6  )�      C  , , 6  � 6   ? 6�   ? 6�  � 6  �      C  , , 6  (A 6  (� 6�  (� 6�  (A 6  (A      C  , , 6  /{ 6  0% 6�  0% 6�  /{ 6  /{      C  , , 6  [ 6   6�   6�  [ 6  [      C  , , 6  #� 6  $� 6�  $� 6�  #� 6  #�      C  , , 6  � 6  [ 6�  [ 6�  � 6  �      C  , , 6  0� 6  1� 6�  1� 6�  0� 6  0�      C  , , 6  +% 6  +� 6�  +� 6�  +% 6  +%      C  , , 6  "y 6  ## 6�  ## 6�  "y 6  "y      C  , , :G  .	 :G  .� :�  .� :�  .	 :G  .	      C  , , ;�  .	 ;�  .� <Y  .� <Y  .	 ;�  .	      C  , , =  .	 =  .� =�  .� =�  .	 =  .	      C  , , >  .	 >  .� ?)  .� ?)  .	 >  .	      C  , , ?�  .	 ?�  .� @�  .� @�  .	 ?�  .	      C  , , IG  -� IG  .; I�  .; I�  -� IG  -�      C  , , K�  -� K�  .; L?  .; L?  -� K�  -�      C  , , M�  -� M�  .; N�  .; N�  -� M�  -�      C  , , 7w  2_ 7w  3	 8!  3	 8!  2_ 7w  2_      C  , , 8�  2_ 8�  3	 9�  3	 9�  2_ 8�  2_      C  , , :G  2_ :G  3	 :�  3	 :�  2_ :G  2_      C  , , =  0� =  1� =�  1� =�  0� =  0�      C  , , 7w  ,� 7w  -A 8!  -A 8!  ,� 7w  ,�      C  , , 8�  ,� 8�  -A 9�  -A 9�  ,� 8�  ,�      C  , , :G  ,� :G  -A :�  -A :�  ,� :G  ,�      C  , , ;�  ,� ;�  -A <Y  -A <Y  ,� ;�  ,�      C  , , =  ,� =  -A =�  -A =�  ,� =  ,�      C  , , >  ,� >  -A ?)  -A ?)  ,� >  ,�      C  , , ?�  ,� ?�  -A @�  -A @�  ,� ?�  ,�      C  , , IG  ,) IG  ,� I�  ,� I�  ,) IG  ,)      C  , , K�  ,) K�  ,� L?  ,� L?  ,) K�  ,)      C  , , M�  ,) M�  ,� N�  ,� N�  ,) M�  ,)      C  , , >  0� >  1� ?)  1� ?)  0� >  0�      C  , , :G  3� :G  4{ :�  4{ :�  3� :G  3�      C  , , ?�  0� ?�  1� @�  1� @�  0� ?�  0�      C  , , IG  0a IG  1 I�  1 I�  0a IG  0a      C  , , K�  0a K�  1 L?  1 L?  0a K�  0a      C  , , M�  0a M�  1 N�  1 N�  0a M�  0a      C  , , ;�  +% ;�  +� <Y  +� <Y  +% ;�  +%      C  , , >  +% >  +� ?)  +� ?)  +% >  +%      C  , , 7w  &� 7w  'y 8!  'y 8!  &� 7w  &�      C  , , 8�  &� 8�  'y 9�  'y 9�  &� 8�  &�      C  , , :G  &� :G  'y :�  'y :�  &� :G  &�      C  , , ;�  &� ;�  'y <Y  'y <Y  &� ;�  &�      C  , , =  &� =  'y =�  'y =�  &� =  &�      C  , , >  &� >  'y ?)  'y ?)  &� >  &�      C  , , ?�  &� ?�  'y @�  'y @�  &� ?�  &�      C  , , H   ') H   '� H�  '� H�  ') H   ')      C  , , 7w  )� 7w  *] 8!  *] 8!  )� 7w  )�      C  , , 8�  )� 8�  *] 9�  *] 9�  )� 8�  )�      C  , , :G  )� :G  *] :�  *] :�  )� :G  )�      C  , , ;�  )� ;�  *] <Y  *] <Y  )� ;�  )�      C  , , =  )� =  *] =�  *] =�  )� =  )�      C  , , >  )� >  *] ?)  *] ?)  )� >  )�      C  , , ?�  )� ?�  *] @�  *] @�  )� ?�  )�      C  , , IG  )Y IG  * I�  * I�  )Y IG  )Y      C  , , K�  )Y K�  * L?  * L?  )Y K�  )Y      C  , , M�  )Y M�  * N�  * N�  )Y M�  )Y      C  , , ;�  2_ ;�  3	 <Y  3	 <Y  2_ ;�  2_      C  , , =  2_ =  3	 =�  3	 =�  2_ =  2_      C  , , >  2_ >  3	 ?)  3	 ?)  2_ >  2_      C  , , ?�  2_ ?�  3	 @�  3	 @�  2_ ?�  2_      C  , , IG  1� IG  2s I�  2s I�  1� IG  1�      C  , , K�  1� K�  2s L?  2s L?  1� K�  1�      C  , , M�  1� M�  2s N�  2s N�  1� M�  1�      C  , , ;�  3� ;�  4{ <Y  4{ <Y  3� ;�  3�      C  , , Jn  ') Jn  '� K  '� K  ') Jn  ')      C  , , L�  ') L�  '� Mf  '� Mf  ') L�  ')      C  , , 7w  (A 7w  (� 8!  (� 8!  (A 7w  (A      C  , , 8�  (A 8�  (� 9�  (� 9�  (A 8�  (A      C  , , :G  (A :G  (� :�  (� :�  (A :G  (A      C  , , ;�  (A ;�  (� <Y  (� <Y  (A ;�  (A      C  , , =  (A =  (� =�  (� =�  (A =  (A      C  , , >  (A >  (� ?)  (� ?)  (A >  (A      C  , , ?�  (A ?�  (� @�  (� @�  (A ?�  (A      C  , , ?�  +% ?�  +� @�  +� @�  +% ?�  +%      C  , , 7w  /{ 7w  0% 8!  0% 8!  /{ 7w  /{      C  , , 8�  /{ 8�  0% 9�  0% 9�  /{ 8�  /{      C  , , :G  /{ :G  0% :�  0% :�  /{ :G  /{      C  , , ;�  /{ ;�  0% <Y  0% <Y  /{ ;�  /{      C  , , =  /{ =  0% =�  0% =�  /{ =  /{      C  , , >  /{ >  0% ?)  0% ?)  /{ >  /{      C  , , ?�  /{ ?�  0% @�  0% @�  /{ ?�  /{      C  , , IG  .� IG  /� I�  /� I�  .� IG  .�      C  , , K�  .� K�  /� L?  /� L?  .� K�  .�      C  , , M�  .� M�  /� N�  /� N�  .� M�  .�      C  , , 7w  3� 7w  4{ 8!  4{ 8!  3� 7w  3�      C  , , IG  *� IG  +k I�  +k I�  *� IG  *�      C  , , K�  *� K�  +k L?  +k L?  *� K�  *�      C  , , =  3� =  4{ =�  4{ =�  3� =  3�      C  , , >  3� >  4{ ?)  4{ ?)  3� >  3�      C  , , ?�  3� ?�  4{ @�  4{ @�  3� ?�  3�      C  , , IG  31 IG  3� I�  3� I�  31 IG  31      C  , , K�  31 K�  3� L?  3� L?  31 K�  31      C  , , M�  31 M�  3� N�  3� N�  31 M�  31      C  , , 7w  .	 7w  .� 8!  .� 8!  .	 7w  .	      C  , , 8�  .	 8�  .� 9�  .� 9�  .	 8�  .	      C  , , 7w  0� 7w  1� 8!  1� 8!  0� 7w  0�      C  , , 8�  0� 8�  1� 9�  1� 9�  0� 8�  0�      C  , , :G  0� :G  1� :�  1� :�  0� :G  0�      C  , , ;�  0� ;�  1� <Y  1� <Y  0� ;�  0�      C  , , 8�  3� 8�  4{ 9�  4{ 9�  3� 8�  3�      C  , , 7w  +% 7w  +� 8!  +� 8!  +% 7w  +%      C  , , 8�  +% 8�  +� 9�  +� 9�  +% 8�  +%      C  , , :G  +% :G  +� :�  +� :�  +% :G  +%      C  , , M�  *� M�  +k N�  +k N�  *� M�  *�      C  , , =  +% =  +� =�  +� =�  +% =  +%      C  , , &�  -� &�  .; '�  .; '�  -� &�  -�      C  , , 4�  )� 4�  *] 5Q  *] 5Q  )� 4�  )�      C  , , )&  -� )&  .; )�  .; )�  -� )&  -�      C  , , +t  -� +t  .; ,  .; ,  -� +t  -�      C  , , -�  -� -�  .; .l  .; .l  -� -�  -�      C  , , 1�  .	 1�  .� 2�  .� 2�  .	 1�  .	      C  , , 3?  .	 3?  .� 3�  .� 3�  .	 3?  .	      C  , , $�  31 $�  3� %4  3� %4  31 $�  31      C  , , �  .� �  /�  �  /�  �  .� �  .�      C  , , "<  .� "<  /� "�  /� "�  .� "<  .�      C  , , $�  .� $�  /� %4  /� %4  .� $�  .�      C  , , &�  .� &�  /� '�  /� '�  .� &�  .�      C  , , )&  .� )&  /� )�  /� )�  .� )&  .�      C  , , 4�  3� 4�  4{ 5Q  4{ 5Q  3� 4�  3�      C  , , +t  .� +t  /� ,  /� ,  .� +t  .�      C  , , -�  .� -�  /� .l  /� .l  .� -�  .�      C  , , )&  31 )&  3� )�  3� )�  31 )&  31      C  , , �  ,) �  ,�  �  ,�  �  ,) �  ,)      C  , , "<  ,) "<  ,� "�  ,� "�  ,) "<  ,)      C  , , $�  ,) $�  ,� %4  ,� %4  ,) $�  ,)      C  , , &�  ,) &�  ,� '�  ,� '�  ,) &�  ,)      C  , , 1�  /{ 1�  0% 2�  0% 2�  /{ 1�  /{      C  , , 3?  /{ 3?  0% 3�  0% 3�  /{ 3?  /{      C  , , 4�  /{ 4�  0% 5Q  0% 5Q  /{ 4�  /{      C  , , )&  ,) )&  ,� )�  ,� )�  ,) )&  ,)      C  , , +t  ,) +t  ,� ,  ,� ,  ,) +t  ,)      C  , , 1�  (A 1�  (� 2�  (� 2�  (A 1�  (A      C  , , 3?  (A 3?  (� 3�  (� 3�  (A 3?  (A      C  , , 4�  (A 4�  (� 5Q  (� 5Q  (A 4�  (A      C  , , -�  ,) -�  ,� .l  ,� .l  ,) -�  ,)      C  , , 1�  ,� 1�  -A 2�  -A 2�  ,� 1�  ,�      C  , , 3?  ,� 3?  -A 3�  -A 3�  ,� 3?  ,�      C  , , 4�  ,� 4�  -A 5Q  -A 5Q  ,� 4�  ,�      C  , , 3?  2_ 3?  3	 3�  3	 3�  2_ 3?  2_      C  , , 4�  2_ 4�  3	 5Q  3	 5Q  2_ 4�  2_      C  , , 1�  &� 1�  'y 2�  'y 2�  &� 1�  &�      C  , , 3?  &� 3?  'y 3�  'y 3�  &� 3?  &�      C  , , 4�  &� 4�  'y 5Q  'y 5Q  &� 4�  &�      C  , , 3?  3� 3?  4{ 3�  4{ 3�  3� 3?  3�      C  , , $�  0a $�  1 %4  1 %4  0a $�  0a      C  , , &�  0a &�  1 '�  1 '�  0a &�  0a      C  , , +t  1� +t  2s ,  2s ,  1� +t  1�      C  , , "<  31 "<  3� "�  3� "�  31 "<  31      C  , , �  0a �  1  �  1  �  0a �  0a      C  , , 4�  .	 4�  .� 5Q  .� 5Q  .	 4�  .	      C  , , -�  31 -�  3� .l  3� .l  31 -�  31      C  , , �  )Y �  *  �  *  �  )Y �  )Y      C  , , "<  0a "<  1 "�  1 "�  0a "<  0a      C  , , "<  1� "<  2s "�  2s "�  1� "<  1�      C  , , $�  1� $�  2s %4  2s %4  1� $�  1�      C  , , &�  1� &�  2s '�  2s '�  1� &�  1�      C  , , )&  1� )&  2s )�  2s )�  1� )&  1�      C  , , �  ') �  '� q  '� q  ') �  ')      C  , , !  ') !  '� !�  '� !�  ') !  ')      C  , , )&  0a )&  1 )�  1 )�  0a )&  0a      C  , , +t  0a +t  1 ,  1 ,  0a +t  0a      C  , , -�  0a -�  1 .l  1 .l  0a -�  0a      C  , , 1�  0� 1�  1� 2�  1� 2�  0� 1�  0�      C  , , #c  ') #c  '� $  '� $  ') #c  ')      C  , , 3?  0� 3?  1� 3�  1� 3�  0� 3?  0�      C  , , "<  )Y "<  * "�  * "�  )Y "<  )Y      C  , , $�  )Y $�  * %4  * %4  )Y $�  )Y      C  , , &�  )Y &�  * '�  * '�  )Y &�  )Y      C  , , )&  )Y )&  * )�  * )�  )Y )&  )Y      C  , , +t  )Y +t  * ,  * ,  )Y +t  )Y      C  , , -�  )Y -�  * .l  * .l  )Y -�  )Y      C  , , 1�  )� 1�  *] 2�  *] 2�  )� 1�  )�      C  , , 4�  0� 4�  1� 5Q  1� 5Q  0� 4�  0�      C  , , 3?  )� 3?  *] 3�  *] 3�  )� 3?  )�      C  , , %�  ') %�  '� &[  '� &[  ') %�  ')      C  , , '�  ') '�  '� (�  '� (�  ') '�  ')      C  , , *M  ') *M  '� *�  '� *�  ') *M  ')      C  , , ,�  ') ,�  '� -E  '� -E  ') ,�  ')      C  , , +t  31 +t  3� ,  3� ,  31 +t  31      C  , , �  *� �  +k  �  +k  �  *� �  *�      C  , , "<  *� "<  +k "�  +k "�  *� "<  *�      C  , , $�  *� $�  +k %4  +k %4  *� $�  *�      C  , , &�  *� &�  +k '�  +k '�  *� &�  *�      C  , , )&  *� )&  +k )�  +k )�  *� )&  *�      C  , , +t  *� +t  +k ,  +k ,  *� +t  *�      C  , , -�  *� -�  +k .l  +k .l  *� -�  *�      C  , , 1�  +% 1�  +� 2�  +� 2�  +% 1�  +%      C  , , 3?  +% 3?  +� 3�  +� 3�  +% 3?  +%      C  , , 4�  +% 4�  +� 5Q  +� 5Q  +% 4�  +%      C  , , -�  1� -�  2s .l  2s .l  1� -�  1�      C  , , 1�  2_ 1�  3	 2�  3	 2�  2_ 1�  2_      C  , , &�  31 &�  3� '�  3� '�  31 &�  31      C  , , �  -� �  .;  �  .;  �  -� �  -�      C  , , 1�  3� 1�  4{ 2�  4{ 2�  3� 1�  3�      C  , , "<  -� "<  .; "�  .; "�  -� "<  -�      C  , , $�  -� $�  .; %4  .; %4  -� $�  -�      C  , , �  31 �  3�  �  3�  �  31 �  31      C  , , �  1� �  2s  �  2s  �  1� �  1�      C  , , )&  !u )&  " )�  " )�  !u )&  !u      C  , , +t  !u +t  " ,  " ,  !u +t  !u      C  , , -�  !u -�  " .l  " .l  !u -�  !u      C  , , 1�  ! 1�  !� 2�  !� 2�  ! 1�  !      C  , , 3?  ! 3?  !� 3�  !� 3�  ! 3?  !      C  , , '�  % '�  %� (�  %� (�  % '�  %      C  , , *M  % *M  %� *�  %� *�  % *M  %      C  , , ,�  % ,�  %� -E  %� -E  % ,�  %      C  , , 4�  ! 4�  !� 5Q  !� 5Q  ! 4�  !      C  , , �  !u �  "  �  "  �  !u �  !u      C  , , "<  !u "<  " "�  " "�  !u "<  !u      C  , , �  � �    �    �  � �  �      C  , , "<  � "<   "�   "�  � "<  �      C  , , $�  � $�   %4   %4  � $�  �      C  , , &�  � &�   '�   '�  � &�  �      C  , , )&  � )&   )�   )�  � )&  �      C  , , +t  � +t   ,   ,  � +t  �      C  , , �  � �  O  �  O  �  � �  �      C  , , "<  � "<  O "�  O "�  � "<  �      C  , , $�  � $�  O %4  O %4  � $�  �      C  , , &�  � &�  O '�  O '�  � &�  �      C  , , )&  � )&  O )�  O )�  � )&  �      C  , , +t  � +t  O ,  O ,  � +t  �      C  , , -�  � -�  O .l  O .l  � -�  �      C  , , �  = �  �  �  �  �  = �  =      C  , , "<  = "<  � "�  � "�  = "<  =      C  , , 1�  [ 1�   2�   2�  [ 1�  [      C  , , 3?  [ 3?   3�   3�  [ 3?  [      C  , , 4�  [ 4�   5Q   5Q  [ 4�  [      C  , , 1�  # 1�  � 2�  � 2�  # 1�  #      C  , , $�  = $�  � %4  � %4  = $�  =      C  , , &�  = &�  � '�  � '�  = &�  =      C  , , )&  = )&  � )�  � )�  = )&  =      C  , , +t  = +t  � ,  � ,  = +t  =      C  , , -�  = -�  � .l  � .l  = -�  =      C  , , 1�  � 1�  [ 2�  [ 2�  � 1�  �      C  , , 3?  # 3?  � 3�  � 3�  # 3?  #      C  , , 4�  # 4�  � 5Q  � 5Q  # 4�  #      C  , , �  % �  %� q  %� q  % �  %      C  , , !  % !  %� !�  %� !�  % !  %      C  , , 1�  #� 1�  $� 2�  $� 2�  #� 1�  #�      C  , , 3?  #� 3?  $� 3�  $� 3�  #� 3?  #�      C  , , 4�  #� 4�  $� 5Q  $� 5Q  #� 4�  #�      C  , , #c  % #c  %� $  %� $  % #c  %      C  , , %�  % %�  %� &[  %� &[  % %�  %      C  , , -�  � -�   .l   .l  � -�  �      C  , , �    �   �  �   �  �    �         C  , , "<    "<   � "�   � "�    "<         C  , , $�    $�   � %4   � %4    $�         C  , , &�    &�   � '�   � '�    &�         C  , , )&    )&   � )�   � )�    )&         C  , , 3?  � 3?  [ 3�  [ 3�  � 3?  �      C  , , 4�  � 4�  [ 5Q  [ 5Q  � 4�  �      C  , , �  m �    �    �  m �  m      C  , , "<  m "<   "�   "�  m "<  m      C  , , $�  m $�   %4   %4  m $�  m      C  , , &�  m &�   '�   '�  m &�  m      C  , , )&  m )&   )�   )�  m )&  m      C  , , +t  m +t   ,   ,  m +t  m      C  , , -�  m -�   .l   .l  m -�  m      C  , , +t    +t   � ,   � ,    +t         C  , , -�    -�   � .l   � .l    -�         C  , , 1�  � 1�   ? 2�   ? 2�  � 1�  �      C  , , 1�  � 1�  w 2�  w 2�  � 1�  �      C  , , 3?  � 3?  w 3�  w 3�  � 3?  �      C  , , 4�  � 4�  w 5Q  w 5Q  � 4�  �      C  , , 1�  ? 1�  � 2�  � 2�  ? 1�  ?      C  , , �   �  �  �  �  �   �        C  , , "<   "<  � "�  � "�   "<        C  , , $�   $�  � %4  � %4   $�        C  , , &�   &�  � '�  � '�   &�        C  , , )&   )&  � )�  � )�   )&        C  , , +t   +t  � ,  � ,   +t        C  , , -�   -�  � .l  � .l   -�        C  , , 3?  � 3?   ? 3�   ? 3�  � 3?  �      C  , , 4�  � 4�   ? 5Q   ? 5Q  � 4�  �      C  , , �  "� �  #�  �  #�  �  "� �  "�      C  , , "<  "� "<  #� "�  #� "�  "� "<  "�      C  , , $�  "� $�  #� %4  #� %4  "� $�  "�      C  , , &�  "� &�  #� '�  #� '�  "� &�  "�      C  , , )&  "� )&  #� )�  #� )�  "� )&  "�      C  , , +t  "� +t  #� ,  #� ,  "� +t  "�      C  , , -�  "� -�  #� .l  #� .l  "� -�  "�      C  , , 1�  "y 1�  ## 2�  ## 2�  "y 1�  "y      C  , , 3?  "y 3?  ## 3�  ## 3�  "y 3?  "y      C  , , 4�  "y 4�  ## 5Q  ## 5Q  "y 4�  "y      C  , , 3?  ? 3?  � 3�  � 3�  ? 3?  ?      C  , , 4�  ? 4�  � 5Q  � 5Q  ? 4�  ?      C  , , $�  !u $�  " %4  " %4  !u $�  !u      C  , , &�  !u &�  " '�  " '�  !u &�  !u      C  , , 7w  # 7w  � 8!  � 8!  # 7w  #      C  , , 8�  # 8�  � 9�  � 9�  # 8�  #      C  , , :G  # :G  � :�  � :�  # :G  #      C  , , ;�  # ;�  � <Y  � <Y  # ;�  #      C  , , =  # =  � =�  � =�  # =  #      C  , , >  # >  � ?)  � ?)  # >  #      C  , , ?�  # ?�  � @�  � @�  # ?�  #      C  , , D�  � D�  O EU  O EU  � D�  �      C  , , F�  � F�  O G�  O G�  � F�  �      C  , , IG  � IG  O I�  O I�  � IG  �      C  , , K�  � K�  O L?  O L?  � K�  �      C  , , M�  � M�  O N�  O N�  � M�  �      C  , , Jn  % Jn  %� K  %� K  % Jn  %      C  , , L�  % L�  %� Mf  %� Mf  % L�  %      C  , , H   % H   %� H�  %� H�  % H   %      C  , , D�  !u D�  " EU  " EU  !u D�  !u      C  , , F�  !u F�  " G�  " G�  !u F�  !u      C  , , IG  !u IG  " I�  " I�  !u IG  !u      C  , , K�  !u K�  " L?  " L?  !u K�  !u      C  , , M�  !u M�  " N�  " N�  !u M�  !u      C  , , D�    D�   � EU   � EU    D�         C  , , F�    F�   � G�   � G�    F�         C  , , IG    IG   � I�   � I�    IG         C  , , K�    K�   � L?   � L?    K�         C  , , M�    M�   � N�   � N�    M�         C  , , D�  "� D�  #� EU  #� EU  "� D�  "�      C  , , F�  "� F�  #� G�  #� G�  "� F�  "�      C  , , IG  "� IG  #� I�  #� I�  "� IG  "�      C  , , K�  "� K�  #� L?  #� L?  "� K�  "�      C  , , M�  "� M�  #� N�  #� N�  "� M�  "�      C  , , ?�  ! ?�  !� @�  !� @�  ! ?�  !      C  , , =  #� =  $� =�  $� =�  #� =  #�      C  , , >  #� >  $� ?)  $� ?)  #� >  #�      C  , , ?�  #� ?�  $� @�  $� @�  #� ?�  #�      C  , , 7w  � 7w   ? 8!   ? 8!  � 7w  �      C  , , 7w  #� 7w  $� 8!  $� 8!  #� 7w  #�      C  , , 8�  #� 8�  $� 9�  $� 9�  #� 8�  #�      C  , , :G  #� :G  $� :�  $� :�  #� :G  #�      C  , , 8�  � 8�   ? 9�   ? 9�  � 8�  �      C  , , :G  � :G   ? :�   ? :�  � :G  �      C  , , ;�  ! ;�  !� <Y  !� <Y  ! ;�  !      C  , , =  ! =  !� =�  !� =�  ! =  !      C  , , >  ! >  !� ?)  !� ?)  ! >  !      C  , , 8�  ! 8�  !� 9�  !� 9�  ! 8�  !      C  , , :G  ! :G  !� :�  !� :�  ! :G  !      C  , , 7w  ! 7w  !� 8!  !� 8!  ! 7w  !      C  , , 7w  "y 7w  ## 8!  ## 8!  "y 7w  "y      C  , , 8�  "y 8�  ## 9�  ## 9�  "y 8�  "y      C  , , :G  "y :G  ## :�  ## :�  "y :G  "y      C  , , ;�  "y ;�  ## <Y  ## <Y  "y ;�  "y      C  , , =  "y =  ## =�  ## =�  "y =  "y      C  , , >  "y >  ## ?)  ## ?)  "y >  "y      C  , , ?�  "y ?�  ## @�  ## @�  "y ?�  "y      C  , , ;�  � ;�   ? <Y   ? <Y  � ;�  �      C  , , =  � =   ? =�   ? =�  � =  �      C  , , >  � >   ? ?)   ? ?)  � >  �      C  , , ?�  � ?�   ? @�   ? @�  � ?�  �      C  , , ;�  #� ;�  $� <Y  $� <Y  #� ;�  #�      C  , , >  ? >  � ?)  � ?)  ? >  ?      C  , , ?�  ? ?�  � @�  � @�  ? ?�  ?      C  , , >  � >  [ ?)  [ ?)  � >  �      C  , , ?�  � ?�  [ @�  [ @�  � ?�  �      C  , , 8�  � 8�  w 9�  w 9�  � 8�  �      C  , , 7w  [ 7w   8!   8!  [ 7w  [      C  , , 8�  [ 8�   9�   9�  [ 8�  [      C  , , :G  [ :G   :�   :�  [ :G  [      C  , , ;�  [ ;�   <Y   <Y  [ ;�  [      C  , , =  [ =   =�   =�  [ =  [      C  , , >  [ >   ?)   ?)  [ >  [      C  , , ?�  [ ?�   @�   @�  [ ?�  [      C  , , :G  � :G  w :�  w :�  � :G  �      C  , , ;�  � ;�  w <Y  w <Y  � ;�  �      C  , , ;�  ? ;�  � <Y  � <Y  ? ;�  ?      C  , , =  � =  w =�  w =�  � =  �      C  , , >  � >  w ?)  w ?)  � >  �      C  , , ?�  � ?�  w @�  w @�  � ?�  �      C  , , 7w  � 7w  w 8!  w 8!  � 7w  �      C  , , 7w  � 7w  [ 8!  [ 8!  � 7w  �      C  , , 8�  � 8�  [ 9�  [ 9�  � 8�  �      C  , , :G  � :G  [ :�  [ :�  � :G  �      C  , , ;�  � ;�  [ <Y  [ <Y  � ;�  �      C  , , =  � =  [ =�  [ =�  � =  �      C  , , =  ? =  � =�  � =�  ? =  ?      C  , , 7w  ? 7w  � 8!  � 8!  ? 7w  ?      C  , , 8�  ? 8�  � 9�  � 9�  ? 8�  ?      C  , , :G  ? :G  � :�  � :�  ? :G  ?      C  , , K�  � K�   L?   L?  � K�  �      C  , , M�  � M�   N�   N�  � M�  �      C  , , F�   F�  � G�  � G�   F�        C  , , IG   IG  � I�  � I�   IG        C  , , K�   K�  � L?  � L?   K�        C  , , F�  m F�   G�   G�  m F�  m      C  , , IG  m IG   I�   I�  m IG  m      C  , , K�  m K�   L?   L?  m K�  m      C  , , M�  m M�   N�   N�  m M�  m      C  , , D�  � D�   EU   EU  � D�  �      C  , , F�  � F�   G�   G�  � F�  �      C  , , M�   M�  � N�  � N�   M�        C  , , D�  m D�   EU   EU  m D�  m      C  , , D�  = D�  � EU  � EU  = D�  =      C  , , F�  = F�  � G�  � G�  = F�  =      C  , , IG  = IG  � I�  � I�  = IG  =      C  , , K�  = K�  � L?  � L?  = K�  =      C  , , M�  = M�  � N�  � N�  = M�  =      C  , , D�   D�  � EU  � EU   D�        C  , , IG  � IG   I�   I�  � IG  �      C  , ,  ������  �����I  �*���I  �*����  ������      C  , ,  ������  ������  �*����  �*����  ������      C  , ,  �����/  ������  �*����  �*���/  �����/      C  , ,  ����ϕ  �����?  �*���?  �*��ϕ  ����ϕ      C  , ,  ������  ����·  �*��·  �*����  ������      C  , ,  �����%  ������  �*����  �*���%  �����%      C  , ,   1�   2s �  2s �  1�   1�      C  , , h  1� h  2s   2s   1� h  1�      C  , , �  1� �  2s `  2s `  1� �  1�      C  , ,   1�   2s �  2s �  1�   1�      C  , , �  *� �  +k >  +k >  *� �  *�      C  , , �  *� �  +k 	�  +k 	�  *� �  *�      C  , , 0  *� 0  +k �  +k �  *� 0  *�      C  , , ~  *� ~  +k (  +k (  *� ~  *�      C  , , �  *� �  +k v  +k v  *� �  *�      C  , ,   *�   +k �  +k �  *�   *�      C  , , h  *� h  +k   +k   *� h  *�      C  , , �  *� �  +k `  +k `  *� �  *�      C  , ,   *�   +k �  +k �  *�   *�      C  , , R  *� R  +k �  +k �  *� R  *�      C  , , �  ,) �  ,� >  ,� >  ,) �  ,)      C  , , �  ,) �  ,� 	�  ,� 	�  ,) �  ,)      C  , , 0  ,) 0  ,� �  ,� �  ,) 0  ,)      C  , , ~  ,) ~  ,� (  ,� (  ,) ~  ,)      C  , , �  ,) �  ,� v  ,� v  ,) �  ,)      C  , ,   ,)   ,� �  ,� �  ,)   ,)      C  , , h  ,) h  ,�   ,�   ,) h  ,)      C  , , �  ,) �  ,� `  ,� `  ,) �  ,)      C  , ,   ,)   ,� �  ,� �  ,)   ,)      C  , , R  ,) R  ,� �  ,� �  ,) R  ,)      C  , , R  1� R  2s �  2s �  1� R  1�      C  , , �  31 �  3� >  3� >  31 �  31      C  , , �  31 �  3� 	�  3� 	�  31 �  31      C  , , 0  31 0  3� �  3� �  31 0  31      C  , , ~  31 ~  3� (  3� (  31 ~  31      C  , , �  31 �  3� v  3� v  31 �  31      C  , ,   31   3� �  3� �  31   31      C  , , h  31 h  3�   3�   31 h  31      C  , , �  31 �  3� `  3� `  31 �  31      C  , ,   31   3� �  3� �  31   31      C  , , R  31 R  3� �  3� �  31 R  31      C  , , �  .� �  /� >  /� >  .� �  .�      C  , , �  .� �  /� 	�  /� 	�  .� �  .�      C  , , 0  .� 0  /� �  /� �  .� 0  .�      C  , , ~  .� ~  /� (  /� (  .� ~  .�      C  , , �  .� �  /� v  /� v  .� �  .�      C  , ,   .�   /� �  /� �  .�   .�      C  , , h  .� h  /�   /�   .� h  .�      C  , , �  .� �  /� `  /� `  .� �  .�      C  , ,   .�   /� �  /� �  .�   .�      C  , , R  .� R  /� �  /� �  .� R  .�      C  , , �  0a �  1 >  1 >  0a �  0a      C  , , �  0a �  1 	�  1 	�  0a �  0a      C  , , 0  0a 0  1 �  1 �  0a 0  0a      C  , , ~  0a ~  1 (  1 (  0a ~  0a      C  , , �  0a �  1 v  1 v  0a �  0a      C  , ,   0a   1 �  1 �  0a   0a      C  , , h  0a h  1   1   0a h  0a      C  , , �  0a �  1 `  1 `  0a �  0a      C  , ,   0a   1 �  1 �  0a   0a      C  , , R  0a R  1 �  1 �  0a R  0a      C  , , �  1� �  2s >  2s >  1� �  1�      C  , , �  1� �  2s 	�  2s 	�  1� �  1�      C  , , 0  1� 0  2s �  2s �  1� 0  1�      C  , , ~  1� ~  2s (  2s (  1� ~  1�      C  , , �  1� �  2s v  2s v  1� �  1�      C  , , �  -� �  .; >  .; >  -� �  -�      C  , , �  -� �  .; 	�  .; 	�  -� �  -�      C  , , 0  -� 0  .; �  .; �  -� 0  -�      C  , , ~  -� ~  .; (  .; (  -� ~  -�      C  , , �  -� �  .; v  .; v  -� �  -�      C  , , R  )Y R  * �  * �  )Y R  )Y      C  , ,   -�   .; �  .; �  -�   -�      C  , , h  -� h  .;   .;   -� h  -�      C  , , �  -� �  .; `  .; `  -� �  -�      C  , ,   -�   .; �  .; �  -�   -�      C  , , R  -� R  .; �  .; �  -� R  -�      C  , , m  ') m  '�   '�   ') m  ')      C  , , �  ') �  '� e  '� e  ') �  ')      C  , , 
	  ') 
	  '� 
�  '� 
�  ') 
	  ')      C  , , W  ') W  '�   '�   ') W  ')      C  , , �  ') �  '� O  '� O  ') �  ')      C  , , �  ') �  '� �  '� �  ') �  ')      C  , , A  ') A  '� �  '� �  ') A  ')      C  , , �  ') �  '� 9  '� 9  ') �  ')      C  , , �  ') �  '� �  '� �  ') �  ')      C  , , +  ') +  '� �  '� �  ') +  ')      C  , , y  ') y  '� #  '� #  ') y  ')      C  , , �  )Y �  * >  * >  )Y �  )Y      C  , , �  )Y �  * 	�  * 	�  )Y �  )Y      C  , , 0  )Y 0  * �  * �  )Y 0  )Y      C  , , ~  )Y ~  * (  * (  )Y ~  )Y      C  , , �  )Y �  * v  * v  )Y �  )Y      C  , ,   )Y   * �  * �  )Y   )Y      C  , , h  )Y h  *   *   )Y h  )Y      C  , , �  )Y �  * `  * `  )Y �  )Y      C  , ,   )Y   * �  * �  )Y   )Y      C  , ,  �\  1�  �\  2s  �  2s  �  1�  �\  1�      C  , ,  ��  0a  ��  1  �j  1  �j  0a  ��  0a      C  , ,  �  0a  �  1  ��  1  ��  0a  �  0a      C  , ,  �\  0a  �\  1  �  1  �  0a  �\  0a      C  , ,  ��  .�  ��  /�  �j  /�  �j  .�  ��  .�      C  , ,  ��  -�  ��  .;  �j  .;  �j  -�  ��  -�      C  , ,  �  -�  �  .;  ��  .;  ��  -�  �  -�      C  , ,  �\  -�  �\  .;  �  .;  �  -�  �\  -�      C  , ,  ��  -�  ��  .;  T  .;  T  -�  ��  -�      C  , , �  -� �  .; �  .; �  -� �  -�      C  , , F  -� F  .; �  .; �  -� F  -�      C  , ,  �  .�  �  /�  ��  /�  ��  .�  �  .�      C  , ,  �\  .�  �\  /�  �  /�  �  .�  �\  .�      C  , ,  ��  .�  ��  /�  T  /�  T  .�  ��  .�      C  , , �  .� �  /� �  /� �  .� �  .�      C  , , F  .� F  /� �  /� �  .� F  .�      C  , ,  ��  )Y  ��  *  �j  *  �j  )Y  ��  )Y      C  , ,  �  )Y  �  *  ��  *  ��  )Y  �  )Y      C  , ,  ��  ')  ��  '�  �C  '�  �C  ')  ��  ')      C  , ,  ��  ')  ��  '�  ��  '�  ��  ')  ��  ')      C  , ,  �5  ')  �5  '�  ��  '�  ��  ')  �5  ')      C  , ,  ��  ,)  ��  ,�  T  ,�  T  ,)  ��  ,)      C  , , �  ,) �  ,� �  ,� �  ,) �  ,)      C  , ,  ��  31  ��  3�  T  3�  T  31  ��  31      C  , , �  31 �  3� �  3� �  31 �  31      C  , , F  31 F  3� �  3� �  31 F  31      C  , , F  ,) F  ,� �  ,� �  ,) F  ,)      C  , ,  ��  ')  ��  '�  �-  '�  �-  ')  ��  ')      C  , ,  �  ')  �  '� {  '� {  ')  �  ')      C  , ,   ')   '� �  '� �  ')   ')      C  , ,  �  ,)  �  ,�  ��  ,�  ��  ,)  �  ,)      C  , ,  �\  ,)  �\  ,�  �  ,�  �  ,)  �\  ,)      C  , ,  ��  *�  ��  +k  �j  +k  �j  *�  ��  *�      C  , ,  �  *�  �  +k  ��  +k  ��  *�  �  *�      C  , ,  ��  0a  ��  1  T  1  T  0a  ��  0a      C  , , �  0a �  1 �  1 �  0a �  0a      C  , , F  0a F  1 �  1 �  0a F  0a      C  , ,  �\  *�  �\  +k  �  +k  �  *�  �\  *�      C  , ,  ��  *�  ��  +k  T  +k  T  *�  ��  *�      C  , , �  *� �  +k �  +k �  *� �  *�      C  , , F  *� F  +k �  +k �  *� F  *�      C  , ,  �\  )Y  �\  *  �  *  �  )Y  �\  )Y      C  , ,  ��  )Y  ��  *  T  *  T  )Y  ��  )Y      C  , , �  )Y �  * �  * �  )Y �  )Y      C  , , F  )Y F  * �  * �  )Y F  )Y      C  , ,  ��  ,)  ��  ,�  �j  ,�  �j  ,)  ��  ,)      C  , ,  ��  31  ��  3�  �j  3�  �j  31  ��  31      C  , ,  �  31  �  3�  ��  3�  ��  31  �  31      C  , ,  �\  31  �\  3�  �  3�  �  31  �\  31      C  , ,  ��  1�  ��  2s  �j  2s  �j  1�  ��  1�      C  , ,  �  1�  �  2s  ��  2s  ��  1�  �  1�      C  , ,  ��  1�  ��  2s  T  2s  T  1�  ��  1�      C  , , �  1� �  2s �  2s �  1� �  1�      C  , , F  1� F  2s �  2s �  1� F  1�      C  , ,  ��  m  ��    T    T  m  ��  m      C  , , �  m �   �   �  m �  m      C  , , F  m F   �   �  m F  m      C  , ,  �$  �  �$  O  ��  O  ��  �  �$  �      C  , ,  �r  �  �r  O  �  O  �  �  �r  �      C  , ,  ��  �  ��  O  �j  O  �j  �  ��  �      C  , ,  �  �  �  O  ��  O  ��  �  �  �      C  , ,  �\  �  �\  O  �  O  �  �  �\  �      C  , ,  ��  �  ��  O  T  O  T  �  ��  �      C  , , �  � �  O �  O �  � �  �      C  , ,  ��  %  ��  %�  �C  %�  �C  %  ��  %      C  , ,  ��  %  ��  %�  ��  %�  ��  %  ��  %      C  , ,  �5  %  �5  %�  ��  %�  ��  %  �5  %      C  , ,  �$     �$   �  ��   �  ��     �$         C  , ,  �r     �r   �  �   �  �     �r         C  , ,  ��     ��   �  �j   �  �j     ��         C  , ,  �     �   �  ��   �  ��     �         C  , ,  �\     �\   �  �   �  �     �\         C  , ,  ��     ��   �  T   �  T     ��         C  , ,  ��  %  ��  %�  �-  %�  �-  %  ��  %      C  , ,  �  %  �  %� {  %� {  %  �  %      C  , ,   %   %� �  %� �  %   %      C  , , F  � F  O �  O �  � F  �      C  , ,  �$  !u  �$  "  ��  "  ��  !u  �$  !u      C  , ,  �r  !u  �r  "  �  "  �  !u  �r  !u      C  , , �    �   � �   � �    �         C  , , F    F   � �   � �    F         C  , ,  �$    �$  �  ��  �  ��    �$        C  , ,  �r    �r  �  �  �  �    �r        C  , ,  ��    ��  �  �j  �  �j    ��        C  , ,  �    �  �  ��  �  ��    �        C  , ,  �\    �\  �  �  �  �    �\        C  , ,  ��    ��  �  T  �  T    ��        C  , , �   �  � �  � �   �        C  , , F   F  � �  � �   F        C  , ,  ��  !u  ��  "  �j  "  �j  !u  ��  !u      C  , ,  �  !u  �  "  ��  "  ��  !u  �  !u      C  , ,  �\  !u  �\  "  �  "  �  !u  �\  !u      C  , ,  ��  !u  ��  "  T  "  T  !u  ��  !u      C  , ,  �$  �  �$    ��    ��  �  �$  �      C  , ,  �r  �  �r    �    �  �  �r  �      C  , ,  ��  �  ��    �j    �j  �  ��  �      C  , ,  �  �  �    ��    ��  �  �  �      C  , ,  �\  �  �\    �    �  �  �\  �      C  , ,  ��  �  ��    T    T  �  ��  �      C  , , �  � �   �   �  � �  �      C  , , F  � F   �   �  � F  �      C  , , �  !u �  " �  " �  !u �  !u      C  , , F  !u F  " �  " �  !u F  !u      C  , ,  �$  =  �$  �  ��  �  ��  =  �$  =      C  , ,  �r  =  �r  �  �  �  �  =  �r  =      C  , ,  ��  =  ��  �  �j  �  �j  =  ��  =      C  , ,  �  =  �  �  ��  �  ��  =  �  =      C  , ,  �\  =  �\  �  �  �  �  =  �\  =      C  , ,  ��  =  ��  �  T  �  T  =  ��  =      C  , , �  = �  � �  � �  = �  =      C  , , F  = F  � �  � �  = F  =      C  , ,  �$  m  �$    ��    ��  m  �$  m      C  , ,  �r  m  �r    �    �  m  �r  m      C  , ,  ��  m  ��    �j    �j  m  ��  m      C  , ,  �  m  �    ��    ��  m  �  m      C  , ,  �\  m  �\    �    �  m  �\  m      C  , ,  �$  "�  �$  #�  ��  #�  ��  "�  �$  "�      C  , ,  �r  "�  �r  #�  �  #�  �  "�  �r  "�      C  , ,  ��  "�  ��  #�  �j  #�  �j  "�  ��  "�      C  , ,  �  "�  �  #�  ��  #�  ��  "�  �  "�      C  , ,  �\  "�  �\  #�  �  #�  �  "�  �\  "�      C  , ,  ��  "�  ��  #�  T  #�  T  "�  ��  "�      C  , , �  "� �  #� �  #� �  "� �  "�      C  , , F  "� F  #� �  #� �  "� F  "�      C  , , �  % �  %� �  %� �  % �  %      C  , , +  % +  %� �  %� �  % +  %      C  , , y  % y  %� #  %� #  % y  %      C  , ,   m    �   �  m   m      C  , , h  m h        m h  m      C  , , �  m �   `   `  m �  m      C  , ,   m    �   �  m   m      C  , , R  m R   �   �  m R  m      C  , , �  � �  O v  O v  � �  �      C  , ,   �   O �  O �  �   �      C  , , h  � h  O   O   � h  �      C  , , �  � �  O `  O `  � �  �      C  , , �  !u �  " >  " >  !u �  !u      C  , , �   �  � >  � >   �        C  , , �   �  � 	�  � 	�   �        C  , , 0   0  � �  � �   0        C  , , ~   ~  � (  � (   ~        C  , , �   �  � v  � v   �        C  , , �    �   � >   � >    �         C  , , �    �   � 	�   � 	�    �         C  , , 0    0   � �   � �    0         C  , , ~    ~   � (   � (    ~         C  , , �    �   � v   � v    �         C  , ,        � �   � �             C  , , h    h   �    �     h         C  , , �    �   � `   � `    �         C  , ,        � �   � �             C  , , R    R   � �   � �    R         C  , ,      � �  � �           C  , , h   h  �   �    h        C  , , �   �  � `  � `   �        C  , ,      � �  � �           C  , , R   R  � �  � �   R        C  , , �  !u �  " 	�  " 	�  !u �  !u      C  , , 0  !u 0  " �  " �  !u 0  !u      C  , , ~  !u ~  " (  " (  !u ~  !u      C  , , �  !u �  " v  " v  !u �  !u      C  , ,   !u   " �  " �  !u   !u      C  , , h  !u h  "   "   !u h  !u      C  , , �  !u �  " `  " `  !u �  !u      C  , ,   !u   " �  " �  !u   !u      C  , , R  !u R  " �  " �  !u R  !u      C  , ,   �   O �  O �  �   �      C  , , R  � R  O �  O �  � R  �      C  , , �  � �  O >  O >  � �  �      C  , , �  � �  O 	�  O 	�  � �  �      C  , , 0  � 0  O �  O �  � 0  �      C  , , �  = �  � >  � >  = �  =      C  , , �  � �   >   >  � �  �      C  , , �  � �   	�   	�  � �  �      C  , , 0  � 0   �   �  � 0  �      C  , , ~  � ~   (   (  � ~  �      C  , , �  � �   v   v  � �  �      C  , ,   �    �   �  �   �      C  , , h  � h        � h  �      C  , , �  � �   `   `  � �  �      C  , ,   �    �   �  �   �      C  , , R  � R   �   �  � R  �      C  , , �  = �  � 	�  � 	�  = �  =      C  , , 0  = 0  � �  � �  = 0  =      C  , , ~  = ~  � (  � (  = ~  =      C  , , �  = �  � v  � v  = �  =      C  , ,   =   � �  � �  =   =      C  , , h  = h  �   �   = h  =      C  , , �  = �  � `  � `  = �  =      C  , ,   =   � �  � �  =   =      C  , , R  = R  � �  � �  = R  =      C  , , ~  � ~  O (  O (  � ~  �      C  , , �  m �   >   >  m �  m      C  , , �  m �   	�   	�  m �  m      C  , , 0  m 0   �   �  m 0  m      C  , , ~  m ~   (   (  m ~  m      C  , , �  m �   v   v  m �  m      C  , , m  % m  %�   %�   % m  %      C  , , �  % �  %� e  %� e  % �  %      C  , , 
	  % 
	  %� 
�  %� 
�  % 
	  %      C  , , W  % W  %�   %�   % W  %      C  , , �  % �  %� O  %� O  % �  %      C  , , �  % �  %� �  %� �  % �  %      C  , , A  % A  %� �  %� �  % A  %      C  , , �  % �  %� 9  %� 9  % �  %      C  , , �  "� �  #� >  #� >  "� �  "�      C  , , �  "� �  #� 	�  #� 	�  "� �  "�      C  , , 0  "� 0  #� �  #� �  "� 0  "�      C  , , ~  "� ~  #� (  #� (  "� ~  "�      C  , , �  "� �  #� v  #� v  "� �  "�      C  , ,   "�   #� �  #� �  "�   "�      C  , , h  "� h  #�   #�   "� h  "�      C  , , �  "� �  #� `  #� `  "� �  "�      C  , ,   "�   #� �  #� �  "�   "�      C  , , R  "� R  #� �  #� �  "� R  "�      C  , ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      C  , ,  �1  '.  �1  '�  ��  '�  ��  '.  �1  '.      C  , ,  �  '.  �  '�  �)  '�  �)  '.  �  '.      C  , ,  ��  '.  ��  '�  �w  '�  �w  '.  ��  '.      C  , ,  �  '.  �  '�  ��  '�  ��  '.  �  '.      C  , ,  �i  '.  �i  '�  �  '�  �  '.  �i  '.      C  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C  , ,  �3  	�  �3  
�  ��  
�  ��  	�  �3  	�      C  , ,  ā  	�  ā  
�  �+  
�  �+  	�  ā  	�      C  , ,  ��  	�  ��  
�  �y  
�  �y  	�  ��  	�      C  , ,  �  	�  �  
�  ��  
�  ��  	�  �  	�      C  , ,  �k  	�  �k  
�  �  
�  �  	�  �k  	�      C  , ,  ͹  	�  ͹  
�  �c  
�  �c  	�  ͹  	�      C  , ,  �  	�  �  
�  б  
�  б  	�  �  	�      C  , ,  �p  �  �p  �  �  �  �  �  �p  �      C  , ,  ��  �  ��  �  �h  �  �h  �  ��  �      C  , ,  �  �  �  �  ��  �  ��  �  �  �      C  , ,  �Z  �  �Z  �  �  �  �  �  �Z  �      C  , ,  Ũ  �  Ũ  �  �R  �  �R  �  Ũ  �      C  , ,  ��  �  ��  �  Ƞ  �  Ƞ  �  ��  �      C  , ,  �D  �  �D  �  ��  �  ��  �  �D  �      C  , ,  ̒  �  ̒  �  �<  �  �<  �  ̒  �      C  , ,  ��  �  ��  �  ϊ  �  ϊ  �  ��  �      C  , ,  �.  �  �.  �  ��  �  ��  �  �.  �      C  , ,  �p  �  �p  ;  �  ;  �  �  �p  �      C  , ,  ��  �  ��  ;  �h  ;  �h  �  ��  �      C  , ,  �  �  �  ;  ��  ;  ��  �  �  �      C  , ,  �Z  �  �Z  ;  �  ;  �  �  �Z  �      C  , ,  Ũ  �  Ũ  ;  �R  ;  �R  �  Ũ  �      C  , ,  ��  �  ��  ;  Ƞ  ;  Ƞ  �  ��  �      C  , ,  �D  �  �D  ;  ��  ;  ��  �  �D  �      C  , ,  ̒  �  ̒  ;  �<  ;  �<  �  ̒  �      C  , ,  ��  �  ��  ;  ϊ  ;  ϊ  �  ��  �      C  , ,  �.  �  �.  ;  ��  ;  ��  �  �.  �      C  , ,  �p  )  �p  �  �  �  �  )  �p  )      C  , ,  ��  )  ��  �  �h  �  �h  )  ��  )      C  , ,  �  )  �  �  ��  �  ��  )  �  )      C  , ,  �Z  )  �Z  �  �  �  �  )  �Z  )      C  , ,  Ũ  )  Ũ  �  �R  �  �R  )  Ũ  )      C  , ,  ��  )  ��  �  Ƞ  �  Ƞ  )  ��  )      C  , ,  �D  )  �D  �  ��  �  ��  )  �D  )      C  , ,  ̒  )  ̒  �  �<  �  �<  )  ̒  )      C  , ,  ��  )  ��  �  ϊ  �  ϊ  )  ��  )      C  , ,  �.  )  �.  �  ��  �  ��  )  �.  )      C  , ,  �p  �  �p  k  �  k  �  �  �p  �      C  , ,  ��  �  ��  k  �h  k  �h  �  ��  �      C  , ,  �  �  �  k  ��  k  ��  �  �  �      C  , ,  �Z  �  �Z  k  �  k  �  �  �Z  �      C  , ,  Ũ  �  Ũ  k  �R  k  �R  �  Ũ  �      C  , ,  ��  �  ��  k  Ƞ  k  Ƞ  �  ��  �      C  , ,  �D  �  �D  k  ��  k  ��  �  �D  �      C  , ,  ̒  �  ̒  k  �<  k  �<  �  ̒  �      C  , ,  ��  �  ��  k  ϊ  k  ϊ  �  ��  �      C  , ,  �.  �  �.  k  ��  k  ��  �  �.  �      C  , ,  �p  Y  �p    �    �  Y  �p  Y      C  , ,  ��  Y  ��    �h    �h  Y  ��  Y      C  , ,  �  Y  �    ��    ��  Y  �  Y      C  , ,  �Z  Y  �Z    �    �  Y  �Z  Y      C  , ,  Ũ  Y  Ũ    �R    �R  Y  Ũ  Y      C  , ,  ��  Y  ��    Ƞ    Ƞ  Y  ��  Y      C  , ,  �D  Y  �D    ��    ��  Y  �D  Y      C  , ,  ̒  Y  ̒    �<    �<  Y  ̒  Y      C  , ,  ��  Y  ��    ϊ    ϊ  Y  ��  Y      C  , ,  �.  Y  �.    ��    ��  Y  �.  Y      C  , ,  �p  �  �p  �  �  �  �  �  �p  �      C  , ,  ��  �  ��  �  �h  �  �h  �  ��  �      C  , ,  �  �  �  �  ��  �  ��  �  �  �      C  , ,  �Z  �  �Z  �  �  �  �  �  �Z  �      C  , ,  Ũ  �  Ũ  �  �R  �  �R  �  Ũ  �      C  , ,  ��  �  ��  �  Ƞ  �  Ƞ  �  ��  �      C  , ,  �D  �  �D  �  ��  �  ��  �  �D  �      C  , ,  ̒  �  ̒  �  �<  �  �<  �  ̒  �      C  , ,  ��  �  ��  �  ϊ  �  ϊ  �  ��  �      C  , ,  �.  �  �.  �  ��  �  ��  �  �.  �      C  , ,  �p  �  �p  3  �  3  �  �  �p  �      C  , ,  ��  �  ��  3  �h  3  �h  �  ��  �      C  , ,  �  �  �  3  ��  3  ��  �  �  �      C  , ,  �Z  �  �Z  3  �  3  �  �  �Z  �      C  , ,  Ũ  �  Ũ  3  �R  3  �R  �  Ũ  �      C  , ,  ��  �  ��  3  Ƞ  3  Ƞ  �  ��  �      C  , ,  �D  �  �D  3  ��  3  ��  �  �D  �      C  , ,  ̒  �  ̒  3  �<  3  �<  �  ̒  �      C  , ,  ��  �  ��  3  ϊ  3  ϊ  �  ��  �      C  , ,  �.  �  �.  3  ��  3  ��  �  �.  �      C  , ,  �p  !  �p  �  �  �  �  !  �p  !      C  , ,  ��  !  ��  �  �h  �  �h  !  ��  !      C  , ,  �  !  �  �  ��  �  ��  !  �  !      C  , ,  �Z  !  �Z  �  �  �  �  !  �Z  !      C  , ,  Ũ  !  Ũ  �  �R  �  �R  !  Ũ  !      C  , ,  ��  !  ��  �  Ƞ  �  Ƞ  !  ��  !      C  , ,  �D  !  �D  �  ��  �  ��  !  �D  !      C  , ,  ̒  !  ̒  �  �<  �  �<  !  ̒  !      C  , ,  ��  !  ��  �  ϊ  �  ϊ  !  ��  !      C  , ,  �.  !  �.  �  ��  �  ��  !  �.  !      C  , ,  ��  	�  ��  
�  �A  
�  �A  	�  ��  	�      C  , ,  �����  ����w  �����w  ������  �����      C  , ,  �Z����  �Z���w  ����w  �����  �Z����      C  , ,  Ũ����  Ũ���w  �R���w  �R����  Ũ����      C  , ,  ������  �����w  Ƞ���w  Ƞ����  ������      C  , ,  �D����  �D���w  �����w  ������  �D����      C  , ,  ̒����  ̒���w  �<���w  �<����  ̒����      C  , ,  ������  �����w  ϊ���w  ϊ����  ������      C  , ,  �.����  �.���w  �����w  ������  �.����      C  , ,  ��  �  ��    �A    �A  �  ��  �      C  , ,  ��  �  ��    ��    ��  �  ��  �      C  , ,  �3  �  �3    ��    ��  �  �3  �      C  , ,  ā  �  ā    �+    �+  �  ā  �      C  , ,  ��  �  ��    �y    �y  �  ��  �      C  , ,  �  �  �    ��    ��  �  �  �      C  , ,  �k  �  �k    �    �  �  �k  �      C  , ,  ͹  �  ͹    �c    �c  �  ͹  �      C  , ,  �  �  �    б    б  �  �  �      C  , ,  �p  �  �p  O  �  O  �  �  �p  �      C  , ,  ��  �  ��  O  �h  O  �h  �  ��  �      C  , ,  �  �  �  O  ��  O  ��  �  �  �      C  , ,  �Z  �  �Z  O  �  O  �  �  �Z  �      C  , ,  Ũ  �  Ũ  O  �R  O  �R  �  Ũ  �      C  , ,  ��  �  ��  O  Ƞ  O  Ƞ  �  ��  �      C  , ,  �D  �  �D  O  ��  O  ��  �  �D  �      C  , ,  ̒  �  ̒  O  �<  O  �<  �  ̒  �      C  , ,  ��  �  ��  O  ϊ  O  ϊ  �  ��  �      C  , ,  �.  �  �.  O  ��  O  ��  �  �.  �      C  , ,  �p  =  �p  �  �  �  �  =  �p  =      C  , ,  ��  =  ��  �  �h  �  �h  =  ��  =      C  , ,  �  =  �  �  ��  �  ��  =  �  =      C  , ,  �Z  =  �Z  �  �  �  �  =  �Z  =      C  , ,  Ũ  =  Ũ  �  �R  �  �R  =  Ũ  =      C  , ,  ��  =  ��  �  Ƞ  �  Ƞ  =  ��  =      C  , ,  �D  =  �D  �  ��  �  ��  =  �D  =      C  , ,  ̒  =  ̒  �  �<  �  �<  =  ̒  =      C  , ,  ��  =  ��  �  ϊ  �  ϊ  =  ��  =      C  , ,  �.  =  �.  �  ��  �  ��  =  �.  =      C  , ,  �p  �  �p    �    �  �  �p  �      C  , ,  ��  �  ��    �h    �h  �  ��  �      C  , ,  �  �  �    ��    ��  �  �  �      C  , ,  �Z  �  �Z    �    �  �  �Z  �      C  , ,  Ũ  �  Ũ    �R    �R  �  Ũ  �      C  , ,  ��  �  ��    Ƞ    Ƞ  �  ��  �      C  , ,  �D  �  �D    ��    ��  �  �D  �      C  , ,  ̒  �  ̒    �<    �<  �  ̒  �      C  , ,  ��  �  ��    ϊ    ϊ  �  ��  �      C  , ,  �.  �  �.    ��    ��  �  �.  �      C  , ,  �p  m  �p    �    �  m  �p  m      C  , ,  ��  m  ��    �h    �h  m  ��  m      C  , ,  �  m  �    ��    ��  m  �  m      C  , ,  �Z  m  �Z    �    �  m  �Z  m      C  , ,  Ũ  m  Ũ    �R    �R  m  Ũ  m      C  , ,  ��  m  ��    Ƞ    Ƞ  m  ��  m      C  , ,  �D  m  �D    ��    ��  m  �D  m      C  , ,  ̒  m  ̒    �<    �<  m  ̒  m      C  , ,  ��  m  ��    ϊ    ϊ  m  ��  m      C  , ,  �.  m  �.    ��    ��  m  �.  m      C  , ,  �p     �p   �  �   �  �     �p         C  , ,  ��     ��   �  �h   �  �h     ��         C  , ,  �     �   �  ��   �  ��     �         C  , ,  �Z     �Z   �  �   �  �     �Z         C  , ,  Ũ     Ũ   �  �R   �  �R     Ũ         C  , ,  ��     ��   �  Ƞ   �  Ƞ     ��         C  , ,  �D     �D   �  ��   �  ��     �D         C  , ,  ̒     ̒   �  �<   �  �<     ̒         C  , ,  ��     ��   �  ϊ   �  ϊ     ��         C  , ,  �.     �.   �  ��   �  ��     �.         C  , ,  �p����  �p���G  ����G  �����  �p����      C  , ,  ������  �����G  �h���G  �h����  ������      C  , ,  �����  ����G  �����G  ������  �����      C  , ,  �Z����  �Z���G  ����G  �����  �Z����      C  , ,  Ũ����  Ũ���G  �R���G  �R����  Ũ����      C  , ,  ������  �����G  Ƞ���G  Ƞ����  ������      C  , ,  �D����  �D���G  �����G  ������  �D����      C  , ,  ̒����  ̒���G  �<���G  �<����  ̒����      C  , ,  ������  �����G  ϊ���G  ϊ����  ������      C  , ,  �.����  �.���G  �����G  ������  �.����      C  , ,  �p���5  �p����  �����  ����5  �p���5      C  , ,  �����5  ������  �h����  �h���5  �����5      C  , ,  ����5  �����  ������  �����5  ����5      C  , ,  �Z���5  �Z����  �����  ����5  �Z���5      C  , ,  Ũ���5  Ũ����  �R����  �R���5  Ũ���5      C  , ,  �����5  ������  Ƞ����  Ƞ���5  �����5      C  , ,  �D���5  �D����  ������  �����5  �D���5      C  , ,  ̒���5  ̒����  �<����  �<���5  ̒���5      C  , ,  �����5  ������  ϊ����  ϊ���5  �����5      C  , ,  �.���5  �.����  ������  �����5  �.���5      C  , ,  �p����  �p���w  ����w  �����  �p����      C  , ,  ������  �����w  �h���w  �h����  ������      C  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C  , ,  ��  �  ��    ��    ��  �  ��  �      C  , ,  ��  '.  ��  '�  �O  '�  �O  '.  ��  '.      C  , ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      C  , ,  �A  '.  �A  '�  ��  '�  ��  '.  �A  '.      C  , ,  ��  '.  ��  '�  �9  '�  �9  '.  ��  '.      C  , ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      C  , ,  �+  '.  �+  '�  ��  '�  ��  '.  �+  '.      C  , ,  �y  '.  �y  '�  �#  '�  �#  '.  �y  '.      C  , ,  ��  '.  ��  '�  �q  '�  �q  '.  ��  '.      C  , ,  �  '.  �  '�  ��  '�  ��  '.  �  '.      C  , ,  �c  '.  �c  '�  �  '�  �  '.  �c  '.      C  , ,  �%  '.  �%  '�  ��  '�  ��  '.  �%  '.      C  , ,  �s  '.  �s  '�  �  '�  �  '.  �s  '.      C  , ,  ��  '.  ��  '�  �k  '�  �k  '.  ��  '.      C  , ,  �  '.  �  '�  ��  '�  ��  '.  �  '.      C  , ,  �]  '.  �]  '�  �  '�  �  '.  �]  '.      C  , ,  ��  '.  ��  '�  �U  '�  �U  '.  ��  '.      C  , ,  ��  '.  ��  '�  ��  '�  ��  '.  ��  '.      C  , ,  �G  '.  �G  '�  ��  '�  ��  '.  �G  '.      C  , ,  ��  '.  ��  '�  �?  '�  �?  '.  ��  '.      C  , ,  ^�  '.  ^�  '�  __  '�  __  '.  ^�  '.      C  , ,  j;  '.  j;  '�  j�  '�  j�  '.  j;  '.      C  , ,  l�  '.  l�  '�  m3  '�  m3  '.  l�  '.      C  , ,  n�  '.  n�  '�  o�  '�  o�  '.  n�  '.      C  , ,  a  '.  a  '�  a�  '�  a�  '.  a  '.      C  , ,  q%  '.  q%  '�  q�  '�  q�  '.  q%  '.      C  , ,  ss  '.  ss  '�  t  '�  t  '.  ss  '.      C  , ,  u�  '.  u�  '�  vk  '�  vk  '.  u�  '.      C  , ,  x  '.  x  '�  x�  '�  x�  '.  x  '.      C  , ,  z]  '.  z]  '�  {  '�  {  '.  z]  '.      C  , ,  ��  '.  ��  '�  �e  '�  �e  '.  ��  '.      C  , ,  �	  '.  �	  '�  ��  '�  ��  '.  �	  '.      C  , ,  �W  '.  �W  '�  �  '�  �  '.  �W  '.      C  , ,  cQ  '.  cQ  '�  c�  '�  c�  '.  cQ  '.      C  , ,  e�  '.  e�  '�  fI  '�  fI  '.  e�  '.      C  , ,  g�  '.  g�  '�  h�  '�  h�  '.  g�  '.      C  , ,  ��  -�  ��  .@  �>  .@  �>  -�  ��  -�      C  , ,  ��  36  ��  3�  �>  3�  �>  36  ��  36      C  , ,  ��  0f  ��  1  �>  1  �>  0f  ��  0f      C  , ,  ��  1�  ��  2x  �>  2x  �>  1�  ��  1�      C  , ,  ��  *�  ��  +p  �>  +p  �>  *�  ��  *�      C  , ,  ��  )^  ��  *  �>  *  �>  )^  ��  )^      C  , ,  ��  ,.  ��  ,�  �>  ,�  �>  ,.  ��  ,.      C  , ,  ��  .�  ��  /�  �>  /�  �>  .�  ��  .�      C  , ,  Z  '.  Z  '�  Z�  '�  Z�  '.  Z  '.      C  , ,  \g  '.  \g  '�  ]  '�  ]  '.  \g  '.      C  , ,  y�  �  y�  �  zD  �  zD  �  y�  �      C  , ,  {�  �  {�  �  |�  �  |�  �  {�  �      C  , ,  ~6  �  ~6  �  ~�  �  ~�  �  ~6  �      C  , ,  r�  �  r�  3  sZ  3  sZ  �  r�  �      C  , ,  t�  �  t�  3  u�  3  u�  �  t�  �      C  , ,  wL  �  wL  3  w�  3  w�  �  wL  �      C  , ,  y�  �  y�  3  zD  3  zD  �  y�  �      C  , ,  {�  �  {�  3  |�  3  |�  �  {�  �      C  , ,  ~6  �  ~6  3  ~�  3  ~�  �  ~6  �      C  , ,  ��  �  ��  3  �.  3  �.  �  ��  �      C  , ,  ��  �  ��  3  �|  3  �|  �  ��  �      C  , ,  �   �  �   3  ��  3  ��  �  �   �      C  , ,  �n  �  �n  3  �  3  �  �  �n  �      C  , ,  ��  �  ��  3  �f  3  �f  �  ��  �      C  , ,  ��  �  ��  �  �.  �  �.  �  ��  �      C  , ,  ��  �  ��  �  �|  �  �|  �  ��  �      C  , ,  �   �  �   �  ��  �  ��  �  �   �      C  , ,  �n  �  �n  �  �  �  �  �  �n  �      C  , ,  ��  �  ��  �  �f  �  �f  �  ��  �      C  , ,  r�  !  r�  �  sZ  �  sZ  !  r�  !      C  , ,  t�  !  t�  �  u�  �  u�  !  t�  !      C  , ,  wL  !  wL  �  w�  �  w�  !  wL  !      C  , ,  y�  !  y�  �  zD  �  zD  !  y�  !      C  , ,  {�  !  {�  �  |�  �  |�  !  {�  !      C  , ,  ~6  !  ~6  �  ~�  �  ~�  !  ~6  !      C  , ,  ��  !  ��  �  �.  �  �.  !  ��  !      C  , ,  ��  !  ��  �  �|  �  �|  !  ��  !      C  , ,  �   !  �   �  ��  �  ��  !  �   !      C  , ,  �n  !  �n  �  �  �  �  !  �n  !      C  , ,  ��  !  ��  �  �f  �  �f  !  ��  !      C  , ,  s�  	�  s�  
�  t�  
�  t�  	�  s�  	�      C  , ,  v%  	�  v%  
�  v�  
�  v�  	�  v%  	�      C  , ,  xs  	�  xs  
�  y  
�  y  	�  xs  	�      C  , ,  z�  	�  z�  
�  {k  
�  {k  	�  z�  	�      C  , ,  }  	�  }  
�  }�  
�  }�  	�  }  	�      C  , ,  ]  	�  ]  
�  �  
�  �  	�  ]  	�      C  , ,  ��  	�  ��  
�  �U  
�  �U  	�  ��  	�      C  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C  , ,  �G  	�  �G  
�  ��  
�  ��  	�  �G  	�      C  , ,  ��  	�  ��  
�  �?  
�  �?  	�  ��  	�      C  , ,  ��  Y  ��    �.    �.  Y  ��  Y      C  , ,  ��  Y  ��    �|    �|  Y  ��  Y      C  , ,  �   Y  �     ��    ��  Y  �   Y      C  , ,  �n  Y  �n    �    �  Y  �n  Y      C  , ,  ��  Y  ��    �f    �f  Y  ��  Y      C  , ,  t�  Y  t�    u�    u�  Y  t�  Y      C  , ,  wL  Y  wL    w�    w�  Y  wL  Y      C  , ,  y�  Y  y�    zD    zD  Y  y�  Y      C  , ,  {�  Y  {�    |�    |�  Y  {�  Y      C  , ,  ~6  Y  ~6    ~�    ~�  Y  ~6  Y      C  , ,  r�  �  r�  ;  sZ  ;  sZ  �  r�  �      C  , ,  t�  �  t�  ;  u�  ;  u�  �  t�  �      C  , ,  wL  �  wL  ;  w�  ;  w�  �  wL  �      C  , ,  y�  �  y�  ;  zD  ;  zD  �  y�  �      C  , ,  {�  �  {�  ;  |�  ;  |�  �  {�  �      C  , ,  ~6  �  ~6  ;  ~�  ;  ~�  �  ~6  �      C  , ,  ��  �  ��  ;  �.  ;  �.  �  ��  �      C  , ,  ��  �  ��  ;  �|  ;  �|  �  ��  �      C  , ,  �   �  �   ;  ��  ;  ��  �  �   �      C  , ,  �n  �  �n  ;  �  ;  �  �  �n  �      C  , ,  ��  �  ��  ;  �f  ;  �f  �  ��  �      C  , ,  r�  )  r�  �  sZ  �  sZ  )  r�  )      C  , ,  t�  )  t�  �  u�  �  u�  )  t�  )      C  , ,  wL  )  wL  �  w�  �  w�  )  wL  )      C  , ,  y�  )  y�  �  zD  �  zD  )  y�  )      C  , ,  {�  )  {�  �  |�  �  |�  )  {�  )      C  , ,  ~6  )  ~6  �  ~�  �  ~�  )  ~6  )      C  , ,  ��  )  ��  �  �.  �  �.  )  ��  )      C  , ,  ��  )  ��  �  �|  �  �|  )  ��  )      C  , ,  �   )  �   �  ��  �  ��  )  �   )      C  , ,  �n  )  �n  �  �  �  �  )  �n  )      C  , ,  ��  )  ��  �  �f  �  �f  )  ��  )      C  , ,  r�  �  r�  �  sZ  �  sZ  �  r�  �      C  , ,  t�  �  t�  �  u�  �  u�  �  t�  �      C  , ,  wL  �  wL  �  w�  �  w�  �  wL  �      C  , ,  y�  �  y�  �  zD  �  zD  �  y�  �      C  , ,  {�  �  {�  �  |�  �  |�  �  {�  �      C  , ,  ~6  �  ~6  �  ~�  �  ~�  �  ~6  �      C  , ,  ��  �  ��  �  �.  �  �.  �  ��  �      C  , ,  ��  �  ��  �  �|  �  �|  �  ��  �      C  , ,  r�  �  r�  k  sZ  k  sZ  �  r�  �      C  , ,  t�  �  t�  k  u�  k  u�  �  t�  �      C  , ,  wL  �  wL  k  w�  k  w�  �  wL  �      C  , ,  y�  �  y�  k  zD  k  zD  �  y�  �      C  , ,  {�  �  {�  k  |�  k  |�  �  {�  �      C  , ,  ~6  �  ~6  k  ~�  k  ~�  �  ~6  �      C  , ,  ��  �  ��  k  �.  k  �.  �  ��  �      C  , ,  ��  �  ��  k  �|  k  �|  �  ��  �      C  , ,  �   �  �   k  ��  k  ��  �  �   �      C  , ,  �n  �  �n  k  �  k  �  �  �n  �      C  , ,  ��  �  ��  k  �f  k  �f  �  ��  �      C  , ,  �   �  �   �  ��  �  ��  �  �   �      C  , ,  �n  �  �n  �  �  �  �  �  �n  �      C  , ,  ��  �  ��  �  �f  �  �f  �  ��  �      C  , ,  r�  �  r�  �  sZ  �  sZ  �  r�  �      C  , ,  t�  �  t�  �  u�  �  u�  �  t�  �      C  , ,  wL  �  wL  �  w�  �  w�  �  wL  �      C  , ,  r�  Y  r�    sZ    sZ  Y  r�  Y      C  , ,  ix  !  ix  �  j"  �  j"  !  ix  !      C  , ,  b�  �  b�  �  c8  �  c8  �  b�  �      C  , ,  d�  �  d�  �  e�  �  e�  �  d�  �      C  , ,  g*  �  g*  �  g�  �  g�  �  g*  �      C  , ,  ]�  �  ]�  �  ^�  �  ^�  �  ]�  �      C  , ,  `@  �  `@  �  `�  �  `�  �  `@  �      C  , ,  b�  �  b�  �  c8  �  c8  �  b�  �      C  , ,  d�  �  d�  �  e�  �  e�  �  d�  �      C  , ,  g*  �  g*  �  g�  �  g�  �  g*  �      C  , ,  ix  �  ix  �  j"  �  j"  �  ix  �      C  , ,  k�  �  k�  �  lp  �  lp  �  k�  �      C  , ,  ]�  )  ]�  �  ^�  �  ^�  )  ]�  )      C  , ,  `@  )  `@  �  `�  �  `�  )  `@  )      C  , ,  b�  )  b�  �  c8  �  c8  )  b�  )      C  , ,  d�  )  d�  �  e�  �  e�  )  d�  )      C  , ,  g*  )  g*  �  g�  �  g�  )  g*  )      C  , ,  ix  )  ix  �  j"  �  j"  )  ix  )      C  , ,  k�  )  k�  �  lp  �  lp  )  k�  )      C  , ,  n  )  n  �  n�  �  n�  )  n  )      C  , ,  pb  )  pb  �  q  �  q  )  pb  )      C  , ,  k�  !  k�  �  lp  �  lp  !  k�  !      C  , ,  n  !  n  �  n�  �  n�  !  n  !      C  , ,  pb  !  pb  �  q  �  q  !  pb  !      C  , ,  n  �  n  3  n�  3  n�  �  n  �      C  , ,  pb  �  pb  3  q  3  q  �  pb  �      C  , ,  ]�  �  ]�  3  ^�  3  ^�  �  ]�  �      C  , ,  `@  �  `@  3  `�  3  `�  �  `@  �      C  , ,  b�  �  b�  3  c8  3  c8  �  b�  �      C  , ,  d�  �  d�  3  e�  3  e�  �  d�  �      C  , ,  g*  �  g*  3  g�  3  g�  �  g*  �      C  , ,  ix  �  ix  3  j"  3  j"  �  ix  �      C  , ,  n  �  n  �  n�  �  n�  �  n  �      C  , ,  pb  �  pb  �  q  �  q  �  pb  �      C  , ,  k�  �  k�  3  lp  3  lp  �  k�  �      C  , ,  ]�  !  ]�  �  ^�  �  ^�  !  ]�  !      C  , ,  `@  !  `@  �  `�  �  `�  !  `@  !      C  , ,  _  	�  _  
�  _�  
�  _�  	�  _  	�      C  , ,  ag  	�  ag  
�  b  
�  b  	�  ag  	�      C  , ,  ]�  �  ]�  �  ^�  �  ^�  �  ]�  �      C  , ,  `@  �  `@  �  `�  �  `�  �  `@  �      C  , ,  ]�  �  ]�  ;  ^�  ;  ^�  �  ]�  �      C  , ,  ]�  �  ]�  k  ^�  k  ^�  �  ]�  �      C  , ,  `@  �  `@  k  `�  k  `�  �  `@  �      C  , ,  b�  �  b�  k  c8  k  c8  �  b�  �      C  , ,  d�  �  d�  k  e�  k  e�  �  d�  �      C  , ,  g*  �  g*  k  g�  k  g�  �  g*  �      C  , ,  ix  �  ix  k  j"  k  j"  �  ix  �      C  , ,  k�  �  k�  k  lp  k  lp  �  k�  �      C  , ,  n  �  n  k  n�  k  n�  �  n  �      C  , ,  pb  �  pb  k  q  k  q  �  pb  �      C  , ,  `@  �  `@  ;  `�  ;  `�  �  `@  �      C  , ,  b�  �  b�  ;  c8  ;  c8  �  b�  �      C  , ,  d�  �  d�  ;  e�  ;  e�  �  d�  �      C  , ,  g*  �  g*  ;  g�  ;  g�  �  g*  �      C  , ,  ix  �  ix  ;  j"  ;  j"  �  ix  �      C  , ,  k�  �  k�  ;  lp  ;  lp  �  k�  �      C  , ,  n  �  n  ;  n�  ;  n�  �  n  �      C  , ,  pb  �  pb  ;  q  ;  q  �  pb  �      C  , ,  c�  	�  c�  
�  d_  
�  d_  	�  c�  	�      C  , ,  f  	�  f  
�  f�  
�  f�  	�  f  	�      C  , ,  hQ  	�  hQ  
�  h�  
�  h�  	�  hQ  	�      C  , ,  j�  	�  j�  
�  kI  
�  kI  	�  j�  	�      C  , ,  l�  	�  l�  
�  m�  
�  m�  	�  l�  	�      C  , ,  o;  	�  o;  
�  o�  
�  o�  	�  o;  	�      C  , ,  ix  �  ix  �  j"  �  j"  �  ix  �      C  , ,  k�  �  k�  �  lp  �  lp  �  k�  �      C  , ,  n  �  n  �  n�  �  n�  �  n  �      C  , ,  pb  �  pb  �  q  �  q  �  pb  �      C  , ,  q�  	�  q�  
�  r3  
�  r3  	�  q�  	�      C  , ,  b�  !  b�  �  c8  �  c8  !  b�  !      C  , ,  d�  !  d�  �  e�  �  e�  !  d�  !      C  , ,  ]�  Y  ]�    ^�    ^�  Y  ]�  Y      C  , ,  `@  Y  `@    `�    `�  Y  `@  Y      C  , ,  b�  Y  b�    c8    c8  Y  b�  Y      C  , ,  d�  Y  d�    e�    e�  Y  d�  Y      C  , ,  g*  Y  g*    g�    g�  Y  g*  Y      C  , ,  ix  Y  ix    j"    j"  Y  ix  Y      C  , ,  k�  Y  k�    lp    lp  Y  k�  Y      C  , ,  n  Y  n    n�    n�  Y  n  Y      C  , ,  pb  Y  pb    q    q  Y  pb  Y      C  , ,  g*  !  g*  �  g�  �  g�  !  g*  !      C  , ,  n  =  n  �  n�  �  n�  =  n  =      C  , ,  pb  =  pb  �  q  �  q  =  pb  =      C  , ,  `@  �  `@  O  `�  O  `�  �  `@  �      C  , ,  b�  �  b�  O  c8  O  c8  �  b�  �      C  , ,  ]����5  ]�����  ^�����  ^����5  ]����5      C  , ,  `@���5  `@����  `�����  `����5  `@���5      C  , ,  b����5  b�����  c8����  c8���5  b����5      C  , ,  d����5  d�����  e�����  e����5  d����5      C  , ,  g*���5  g*����  g�����  g����5  g*���5      C  , ,  ix���5  ix����  j"����  j"���5  ix���5      C  , ,  k����5  k�����  lp����  lp���5  k����5      C  , ,  n���5  n����  n�����  n����5  n���5      C  , ,  pb���5  pb����  q����  q���5  pb���5      C  , ,  d�  �  d�  O  e�  O  e�  �  d�  �      C  , ,  g*  �  g*  O  g�  O  g�  �  g*  �      C  , ,  ix  �  ix  O  j"  O  j"  �  ix  �      C  , ,  k�  �  k�  O  lp  O  lp  �  k�  �      C  , ,  n  �  n  O  n�  O  n�  �  n  �      C  , ,  pb  �  pb  O  q  O  q  �  pb  �      C  , ,  ]�  �  ]�    ^�    ^�  �  ]�  �      C  , ,  `@  �  `@    `�    `�  �  `@  �      C  , ,  b�  �  b�    c8    c8  �  b�  �      C  , ,  ]�����  ]����w  ^����w  ^�����  ]�����      C  , ,  `@����  `@���w  `����w  `�����  `@����      C  , ,  b�����  b����w  c8���w  c8����  b�����      C  , ,  d�����  d����w  e����w  e�����  d�����      C  , ,  g*����  g*���w  g����w  g�����  g*����      C  , ,  ix����  ix���w  j"���w  j"����  ix����      C  , ,  k�����  k����w  lp���w  lp����  k�����      C  , ,  n����  n���w  n����w  n�����  n����      C  , ,  pb����  pb���w  q���w  q����  pb����      C  , ,  d�  �  d�    e�    e�  �  d�  �      C  , ,  g*  �  g*    g�    g�  �  g*  �      C  , ,  ix  �  ix    j"    j"  �  ix  �      C  , ,  k�  �  k�    lp    lp  �  k�  �      C  , ,  n  �  n    n�    n�  �  n  �      C  , ,  pb  �  pb    q    q  �  pb  �      C  , ,  ]�  m  ]�    ^�    ^�  m  ]�  m      C  , ,  `@  m  `@    `�    `�  m  `@  m      C  , ,  b�  m  b�    c8    c8  m  b�  m      C  , ,  d�  m  d�    e�    e�  m  d�  m      C  , ,  g*  m  g*    g�    g�  m  g*  m      C  , ,  ix  m  ix    j"    j"  m  ix  m      C  , ,  k�  m  k�    lp    lp  m  k�  m      C  , ,  n  m  n    n�    n�  m  n  m      C  , ,  pb  m  pb    q    q  m  pb  m      C  , ,  ag  �  ag    b    b  �  ag  �      C  , ,  ]�     ]�   �  ^�   �  ^�     ]�         C  , ,  `@     `@   �  `�   �  `�     `@         C  , ,  b�     b�   �  c8   �  c8     b�         C  , ,  d�     d�   �  e�   �  e�     d�         C  , ,  g*     g*   �  g�   �  g�     g*         C  , ,  ix     ix   �  j"   �  j"     ix         C  , ,  k�     k�   �  lp   �  lp     k�         C  , ,  n     n   �  n�   �  n�     n         C  , ,  pb     pb   �  q   �  q     pb         C  , ,  c�  �  c�    d_    d_  �  c�  �      C  , ,  f  �  f    f�    f�  �  f  �      C  , ,  hQ  �  hQ    h�    h�  �  hQ  �      C  , ,  j�  �  j�    kI    kI  �  j�  �      C  , ,  l�  �  l�    m�    m�  �  l�  �      C  , ,  o;  �  o;    o�    o�  �  o;  �      C  , ,  q�  �  q�    r3    r3  �  q�  �      C  , ,  _  �  _    _�    _�  �  _  �      C  , ,  ]�  �  ]�  O  ^�  O  ^�  �  ]�  �      C  , ,  ]�  =  ]�  �  ^�  �  ^�  =  ]�  =      C  , ,  ]�����  ]����G  ^����G  ^�����  ]�����      C  , ,  `@����  `@���G  `����G  `�����  `@����      C  , ,  b�����  b����G  c8���G  c8����  b�����      C  , ,  d�����  d����G  e����G  e�����  d�����      C  , ,  g*����  g*���G  g����G  g�����  g*����      C  , ,  ix����  ix���G  j"���G  j"����  ix����      C  , ,  k�����  k����G  lp���G  lp����  k�����      C  , ,  n����  n���G  n����G  n�����  n����      C  , ,  pb����  pb���G  q���G  q����  pb����      C  , ,  `@  =  `@  �  `�  �  `�  =  `@  =      C  , ,  b�  =  b�  �  c8  �  c8  =  b�  =      C  , ,  d�  =  d�  �  e�  �  e�  =  d�  =      C  , ,  g*  =  g*  �  g�  �  g�  =  g*  =      C  , ,  ix  =  ix  �  j"  �  j"  =  ix  =      C  , ,  k�  =  k�  �  lp  �  lp  =  k�  =      C  , ,  wL  =  wL  �  w�  �  w�  =  wL  =      C  , ,  y�  =  y�  �  zD  �  zD  =  y�  =      C  , ,  {�  =  {�  �  |�  �  |�  =  {�  =      C  , ,  r�  m  r�    sZ    sZ  m  r�  m      C  , ,  t�  m  t�    u�    u�  m  t�  m      C  , ,  wL  m  wL    w�    w�  m  wL  m      C  , ,  y�  m  y�    zD    zD  m  y�  m      C  , ,  {�  m  {�    |�    |�  m  {�  m      C  , ,  r����5  r�����  sZ����  sZ���5  r����5      C  , ,  t����5  t�����  u�����  u����5  t����5      C  , ,  wL���5  wL����  w�����  w����5  wL���5      C  , ,  y����5  y�����  zD����  zD���5  y����5      C  , ,  {����5  {�����  |�����  |����5  {����5      C  , ,  ~6���5  ~6����  ~�����  ~����5  ~6���5      C  , ,  �����5  ������  �.����  �.���5  �����5      C  , ,  �����5  ������  �|����  �|���5  �����5      C  , ,  � ���5  � ����  ������  �����5  � ���5      C  , ,  �n���5  �n����  �����  ����5  �n���5      C  , ,  �����5  ������  �f����  �f���5  �����5      C  , ,  ~6  m  ~6    ~�    ~�  m  ~6  m      C  , ,  ��  m  ��    �.    �.  m  ��  m      C  , ,  ��  m  ��    �|    �|  m  ��  m      C  , ,  �   m  �     ��    ��  m  �   m      C  , ,  �n  m  �n    �    �  m  �n  m      C  , ,  ��  m  ��    �f    �f  m  ��  m      C  , ,  ~6  =  ~6  �  ~�  �  ~�  =  ~6  =      C  , ,  ��  =  ��  �  �.  �  �.  =  ��  =      C  , ,  ��  =  ��  �  �|  �  �|  =  ��  =      C  , ,  �   =  �   �  ��  �  ��  =  �   =      C  , ,  �n  =  �n  �  �  �  �  =  �n  =      C  , ,  ��  =  ��  �  �f  �  �f  =  ��  =      C  , ,  �n  �  �n  O  �  O  �  �  �n  �      C  , ,  ��  �  ��  O  �f  O  �f  �  ��  �      C  , ,  ��  �  ��    �?    �?  �  ��  �      C  , ,  s�  �  s�    t�    t�  �  s�  �      C  , ,  r�     r�   �  sZ   �  sZ     r�         C  , ,  t�     t�   �  u�   �  u�     t�         C  , ,  r�����  r����w  sZ���w  sZ����  r�����      C  , ,  t�����  t����w  u����w  u�����  t�����      C  , ,  wL����  wL���w  w����w  w�����  wL����      C  , ,  y�����  y����w  zD���w  zD����  y�����      C  , ,  {�����  {����w  |����w  |�����  {�����      C  , ,  ~6����  ~6���w  ~����w  ~�����  ~6����      C  , ,  ������  �����w  �.���w  �.����  ������      C  , ,  ������  �����w  �|���w  �|����  ������      C  , ,  � ����  � ���w  �����w  ������  � ����      C  , ,  �n����  �n���w  ����w  �����  �n����      C  , ,  ������  �����w  �f���w  �f����  ������      C  , ,  wL     wL   �  w�   �  w�     wL         C  , ,  y�     y�   �  zD   �  zD     y�         C  , ,  {�     {�   �  |�   �  |�     {�         C  , ,  ~6     ~6   �  ~�   �  ~�     ~6         C  , ,  ��     ��   �  �.   �  �.     ��         C  , ,  ��     ��   �  �|   �  �|     ��         C  , ,  �      �    �  ��   �  ��     �          C  , ,  �n     �n   �  �   �  �     �n         C  , ,  ��     ��   �  �f   �  �f     ��         C  , ,  v%  �  v%    v�    v�  �  v%  �      C  , ,  xs  �  xs    y    y  �  xs  �      C  , ,  z�  �  z�    {k    {k  �  z�  �      C  , ,  }  �  }    }�    }�  �  }  �      C  , ,  ]  �  ]    �    �  �  ]  �      C  , ,  ��  �  ��    �U    �U  �  ��  �      C  , ,  ��  �  ��    ��    ��  �  ��  �      C  , ,  �G  �  �G    ��    ��  �  �G  �      C  , ,  r�  �  r�  O  sZ  O  sZ  �  r�  �      C  , ,  t�  �  t�  O  u�  O  u�  �  t�  �      C  , ,  wL  �  wL  O  w�  O  w�  �  wL  �      C  , ,  y�  �  y�  O  zD  O  zD  �  y�  �      C  , ,  {�  �  {�  O  |�  O  |�  �  {�  �      C  , ,  r�  �  r�    sZ    sZ  �  r�  �      C  , ,  t�  �  t�    u�    u�  �  t�  �      C  , ,  wL  �  wL    w�    w�  �  wL  �      C  , ,  y�  �  y�    zD    zD  �  y�  �      C  , ,  {�  �  {�    |�    |�  �  {�  �      C  , ,  ~6  �  ~6    ~�    ~�  �  ~6  �      C  , ,  r�����  r����G  sZ���G  sZ����  r�����      C  , ,  t�����  t����G  u����G  u�����  t�����      C  , ,  wL����  wL���G  w����G  w�����  wL����      C  , ,  y�����  y����G  zD���G  zD����  y�����      C  , ,  {�����  {����G  |����G  |�����  {�����      C  , ,  ~6����  ~6���G  ~����G  ~�����  ~6����      C  , ,  ������  �����G  �.���G  �.����  ������      C  , ,  ������  �����G  �|���G  �|����  ������      C  , ,  � ����  � ���G  �����G  ������  � ����      C  , ,  �n����  �n���G  ����G  �����  �n����      C  , ,  ������  �����G  �f���G  �f����  ������      C  , ,  ��  �  ��    �.    �.  �  ��  �      C  , ,  ��  �  ��    �|    �|  �  ��  �      C  , ,  �   �  �     ��    ��  �  �   �      C  , ,  �n  �  �n    �    �  �  �n  �      C  , ,  ��  �  ��    �f    �f  �  ��  �      C  , ,  ~6  �  ~6  O  ~�  O  ~�  �  ~6  �      C  , ,  ��  �  ��  O  �.  O  �.  �  ��  �      C  , ,  ��  �  ��  O  �|  O  �|  �  ��  �      C  , ,  �   �  �   O  ��  O  ��  �  �   �      C  , ,  r�  =  r�  �  sZ  �  sZ  =  r�  =      C  , ,  t�  =  t�  �  u�  �  u�  =  t�  =      C  , ,  �  �  �    ��    ��  �  �  �      C  , ,  �  �  �  ;  ��  ;  ��  �  �  �      C  , ,  �  m  �    ��    ��  m  �  m      C  , ,  �  �  �  3  ��  3  ��  �  �  �      C  , ,  �  �  �  �  ��  �  ��  �  �  �      C  , ,  �     �   �  ��   �  ��     �         C  , ,  �����  ����G  �����G  ������  �����      C  , ,  �  Y  �    ��    ��  Y  �  Y      C  , ,  �  �  �  O  ��  O  ��  �  �  �      C  , ,  ����5  �����  ������  �����5  ����5      C  , ,  �  !  �  �  ��  �  ��  !  �  !      C  , ,  �����  ����w  �����w  ������  �����      C  , ,  �  )  �  �  ��  �  ��  )  �  )      C  , ,  �  �  �  �  ��  �  ��  �  �  �      C  , ,  �  =  �  �  ��  �  ��  =  �  =      C  , ,  �  �  �  k  ��  k  ��  �  �  �      C  , ,  �8  �  �8  �  ��  �  ��  �  �8  �      C  , ,  ��  �  ��  �  �0  �  �0  �  ��  �      C  , ,  ��  �  ��  �  �~  �  �~  �  ��  �      C  , ,  �"  �  �"  �  ��  �  ��  �  �"  �      C  , ,  �=  	�  �=  
�  ��  
�  ��  	�  �=  	�      C  , ,  ��  �  ��  ;  �\  ;  �\  �  ��  �      C  , ,  �   �  �   ;  ��  ;  ��  �  �   �      C  , ,  �N  �  �N  ;  ��  ;  ��  �  �N  �      C  , ,  ��  �  ��  ;  �F  ;  �F  �  ��  �      C  , ,  ��  �  ��  ;  ��  ;  ��  �  ��  �      C  , ,  �8  �  �8  ;  ��  ;  ��  �  �8  �      C  , ,  ��  �  ��  ;  �0  ;  �0  �  ��  �      C  , ,  ��  �  ��  ;  �~  ;  �~  �  ��  �      C  , ,  �"  �  �"  ;  ��  ;  ��  �  �"  �      C  , ,  �d  �  �d  ;  �  ;  �  �  �d  �      C  , ,  �d  �  �d  3  �  3  �  �  �d  �      C  , ,  ��  �  ��  3  �\  3  �\  �  ��  �      C  , ,  �   �  �   3  ��  3  ��  �  �   �      C  , ,  �N  �  �N  3  ��  3  ��  �  �N  �      C  , ,  ��  �  ��  3  �F  3  �F  �  ��  �      C  , ,  ��  �  ��  3  ��  3  ��  �  ��  �      C  , ,  �8  �  �8  3  ��  3  ��  �  �8  �      C  , ,  ��  �  ��  3  �0  3  �0  �  ��  �      C  , ,  ��  �  ��  3  �~  3  �~  �  ��  �      C  , ,  �"  �  �"  3  ��  3  ��  �  �"  �      C  , ,  ��  	�  ��  
�  �5  
�  �5  	�  ��  	�      C  , ,  �d  �  �d  �  �  �  �  �  �d  �      C  , ,  ��  �  ��  �  �\  �  �\  �  ��  �      C  , ,  �   �  �   �  ��  �  ��  �  �   �      C  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C  , ,  �N  �  �N  �  ��  �  ��  �  �N  �      C  , ,  ��  �  ��  �  �F  �  �F  �  ��  �      C  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      C  , ,  �8  �  �8  �  ��  �  ��  �  �8  �      C  , ,  ��  �  ��  �  �0  �  �0  �  ��  �      C  , ,  ��  �  ��  �  �~  �  �~  �  ��  �      C  , ,  �'  	�  �'  
�  ��  
�  ��  	�  �'  	�      C  , ,  �"  �  �"  �  ��  �  ��  �  �"  �      C  , ,  �u  	�  �u  
�  �  
�  �  	�  �u  	�      C  , ,  �d  Y  �d    �    �  Y  �d  Y      C  , ,  ��  Y  ��    �\    �\  Y  ��  Y      C  , ,  �   Y  �     ��    ��  Y  �   Y      C  , ,  �N  Y  �N    ��    ��  Y  �N  Y      C  , ,  ��  Y  ��    �F    �F  Y  ��  Y      C  , ,  ��  Y  ��    ��    ��  Y  ��  Y      C  , ,  �8  Y  �8    ��    ��  Y  �8  Y      C  , ,  ��  Y  ��    �0    �0  Y  ��  Y      C  , ,  ��  Y  ��    �~    �~  Y  ��  Y      C  , ,  �"  Y  �"    ��    ��  Y  �"  Y      C  , ,  ��  	�  ��  
�  �m  
�  �m  	�  ��  	�      C  , ,  �  	�  �  
�  ��  
�  ��  	�  �  	�      C  , ,  �_  	�  �_  
�  �	  
�  �	  	�  �_  	�      C  , ,  �d  !  �d  �  �  �  �  !  �d  !      C  , ,  ��  !  ��  �  �\  �  �\  !  ��  !      C  , ,  �   !  �   �  ��  �  ��  !  �   !      C  , ,  �N  !  �N  �  ��  �  ��  !  �N  !      C  , ,  ��  !  ��  �  �F  �  �F  !  ��  !      C  , ,  ��  !  ��  �  ��  �  ��  !  ��  !      C  , ,  �8  !  �8  �  ��  �  ��  !  �8  !      C  , ,  ��  !  ��  �  �0  �  �0  !  ��  !      C  , ,  ��  !  ��  �  �~  �  �~  !  ��  !      C  , ,  �"  !  �"  �  ��  �  ��  !  �"  !      C  , ,  ��  	�  ��  
�  �W  
�  �W  	�  ��  	�      C  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C  , ,  �d  )  �d  �  �  �  �  )  �d  )      C  , ,  ��  )  ��  �  �\  �  �\  )  ��  )      C  , ,  �   )  �   �  ��  �  ��  )  �   )      C  , ,  �N  )  �N  �  ��  �  ��  )  �N  )      C  , ,  ��  )  ��  �  �F  �  �F  )  ��  )      C  , ,  ��  )  ��  �  ��  �  ��  )  ��  )      C  , ,  �8  )  �8  �  ��  �  ��  )  �8  )      C  , ,  ��  )  ��  �  �0  �  �0  )  ��  )      C  , ,  ��  )  ��  �  �~  �  �~  )  ��  )      C  , ,  �"  )  �"  �  ��  �  ��  )  �"  )      C  , ,  �I  	�  �I  
�  ��  
�  ��  	�  �I  	�      C  , ,  �d  �  �d  �  �  �  �  �  �d  �      C  , ,  ��  �  ��  �  �\  �  �\  �  ��  �      C  , ,  �   �  �   �  ��  �  ��  �  �   �      C  , ,  �N  �  �N  �  ��  �  ��  �  �N  �      C  , ,  ��  �  ��  �  �F  �  �F  �  ��  �      C  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      C  , ,  �d  �  �d  k  �  k  �  �  �d  �      C  , ,  ��  �  ��  k  �\  k  �\  �  ��  �      C  , ,  �   �  �   k  ��  k  ��  �  �   �      C  , ,  �N  �  �N  k  ��  k  ��  �  �N  �      C  , ,  ��  �  ��  k  �F  k  �F  �  ��  �      C  , ,  ��  �  ��  k  ��  k  ��  �  ��  �      C  , ,  �8  �  �8  k  ��  k  ��  �  �8  �      C  , ,  ��  �  ��  k  �0  k  �0  �  ��  �      C  , ,  ��  �  ��  k  �~  k  �~  �  ��  �      C  , ,  �"  �  �"  k  ��  k  ��  �  �"  �      C  , ,  ��  !  ��  �  ��  �  ��  !  ��  !      C  , ,  �,  !  �,  �  ��  �  ��  !  �,  !      C  , ,  �z  !  �z  �  �$  �  �$  !  �z  !      C  , ,  ��  !  ��  �  �r  �  �r  !  ��  !      C  , ,  ��  �  ��  3  ��  3  ��  �  ��  �      C  , ,  ��  	�  ��  
�  �w  
�  �w  	�  ��  	�      C  , ,  �  	�  �  
�  ��  
�  ��  	�  �  	�      C  , ,  �i  	�  �i  
�  �  
�  �  	�  �i  	�      C  , ,  ��  	�  ��  
�  �a  
�  �a  	�  ��  	�      C  , ,  �
  �  �
  �  ��  �  ��  �  �
  �      C  , ,  �X  �  �X  �  �  �  �  �  �X  �      C  , ,  ��  �  ��  �  �P  �  �P  �  ��  �      C  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      C  , ,  �B  �  �B  �  ��  �  ��  �  �B  �      C  , ,  �  	�  �  
�  ��  
�  ��  	�  �  	�      C  , ,  ��  �  ��  �  �:  �  �:  �  ��  �      C  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      C  , ,  �,  �  �,  �  ��  �  ��  �  �,  �      C  , ,  �S  	�  �S  
�  ��  
�  ��  	�  �S  	�      C  , ,  �X  )  �X  �  �  �  �  )  �X  )      C  , ,  ��  )  ��  �  �P  �  �P  )  ��  )      C  , ,  ��  )  ��  �  ��  �  ��  )  ��  )      C  , ,  �B  )  �B  �  ��  �  ��  )  �B  )      C  , ,  ��  )  ��  �  �:  �  �:  )  ��  )      C  , ,  ��  )  ��  �  ��  �  ��  )  ��  )      C  , ,  �,  )  �,  �  ��  �  ��  )  �,  )      C  , ,  �z  )  �z  �  �$  �  �$  )  �z  )      C  , ,  ��  )  ��  �  �r  �  �r  )  ��  )      C  , ,  ��  	�  ��  
�  �K  
�  �K  	�  ��  	�      C  , ,  ��  	�  ��  
�  ��  
�  ��  	�  ��  	�      C  , ,  �1  	�  �1  
�  ��  
�  ��  	�  �1  	�      C  , ,  �  	�  �  
�  �)  
�  �)  	�  �  	�      C  , ,  �,  �  �,  3  ��  3  ��  �  �,  �      C  , ,  �z  �  �z  3  �$  3  �$  �  �z  �      C  , ,  ��  Y  ��    �r    �r  Y  ��  Y      C  , ,  ��  �  ��  3  �r  3  �r  �  ��  �      C  , ,  ��  �  ��  ;  �P  ;  �P  �  ��  �      C  , ,  ��  �  ��  ;  ��  ;  ��  �  ��  �      C  , ,  �B  �  �B  ;  ��  ;  ��  �  �B  �      C  , ,  �z  �  �z  �  �$  �  �$  �  �z  �      C  , ,  ��  �  ��  �  �r  �  �r  �  ��  �      C  , ,  ��  �  ��  ;  �:  ;  �:  �  ��  �      C  , ,  ��  �  ��  ;  ��  ;  ��  �  ��  �      C  , ,  �,  �  �,  ;  ��  ;  ��  �  �,  �      C  , ,  �z  �  �z  ;  �$  ;  �$  �  �z  �      C  , ,  ��  �  ��  ;  �r  ;  �r  �  ��  �      C  , ,  �X  Y  �X    �    �  Y  �X  Y      C  , ,  ��  Y  ��    �P    �P  Y  ��  Y      C  , ,  ��  Y  ��    ��    ��  Y  ��  Y      C  , ,  ��  �  ��  3  ��  3  ��  �  ��  �      C  , ,  �
  �  �
  k  ��  k  ��  �  �
  �      C  , ,  �X  �  �X  k  �  k  �  �  �X  �      C  , ,  ��  �  ��  k  �P  k  �P  �  ��  �      C  , ,  ��  �  ��  k  ��  k  ��  �  ��  �      C  , ,  �B  �  �B  k  ��  k  ��  �  �B  �      C  , ,  ��  �  ��  k  �:  k  �:  �  ��  �      C  , ,  ��  �  ��  k  ��  k  ��  �  ��  �      C  , ,  �,  �  �,  k  ��  k  ��  �  �,  �      C  , ,  �z  �  �z  k  �$  k  �$  �  �z  �      C  , ,  ��  �  ��  k  �r  k  �r  �  ��  �      C  , ,  �B  �  �B  3  ��  3  ��  �  �B  �      C  , ,  �
  Y  �
    ��    ��  Y  �
  Y      C  , ,  �
  !  �
  �  ��  �  ��  !  �
  !      C  , ,  �X  !  �X  �  �  �  �  !  �X  !      C  , ,  ��  !  ��  �  �P  �  �P  !  ��  !      C  , ,  ��  !  ��  �  ��  �  ��  !  ��  !      C  , ,  ��  �  ��  3  �:  3  �:  �  ��  �      C  , ,  ��  �  ��  �  �r  �  �r  �  ��  �      C  , ,  �
  )  �
  �  ��  �  ��  )  �
  )      C  , ,  �B  !  �B  �  ��  �  ��  !  �B  !      C  , ,  ��  !  ��  �  �:  �  �:  !  ��  !      C  , ,  �B  Y  �B    ��    ��  Y  �B  Y      C  , ,  ��  Y  ��    �:    �:  Y  ��  Y      C  , ,  ��  Y  ��    ��    ��  Y  ��  Y      C  , ,  �,  Y  �,    ��    ��  Y  �,  Y      C  , ,  �z  Y  �z    �$    �$  Y  �z  Y      C  , ,  �
  �  �
  �  ��  �  ��  �  �
  �      C  , ,  �X  �  �X  �  �  �  �  �  �X  �      C  , ,  ��  �  ��  �  �P  �  �P  �  ��  �      C  , ,  �
  �  �
  ;  ��  ;  ��  �  �
  �      C  , ,  �X  �  �X  ;  �  ;  �  �  �X  �      C  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      C  , ,  �B  �  �B  �  ��  �  ��  �  �B  �      C  , ,  ��  �  ��  �  �:  �  �:  �  ��  �      C  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      C  , ,  �,  �  �,  �  ��  �  ��  �  �,  �      C  , ,  �z  �  �z  �  �$  �  �$  �  �z  �      C  , ,  �
  �  �
  3  ��  3  ��  �  �
  �      C  , ,  �X  �  �X  3  �  3  �  �  �X  �      C  , ,  ��  �  ��  3  �P  3  �P  �  ��  �      C  , ,  ������  �����w  �P���w  �P����  ������      C  , ,  ������  �����w  �����w  ������  ������      C  , ,  �B����  �B���w  �����w  ������  �B����      C  , ,  ������  �����w  �:���w  �:����  ������      C  , ,  ������  �����w  �����w  ������  ������      C  , ,  �,����  �,���w  �����w  ������  �,����      C  , ,  �z����  �z���w  �$���w  �$����  �z����      C  , ,  ������  �����w  �r���w  �r����  ������      C  , ,  ������  �����G  �P���G  �P����  ������      C  , ,  ������  �����G  �����G  ������  ������      C  , ,  �B����  �B���G  �����G  ������  �B����      C  , ,  ������  �����G  �:���G  �:����  ������      C  , ,  ������  �����G  �����G  ������  ������      C  , ,  �,����  �,���G  �����G  ������  �,����      C  , ,  �z����  �z���G  �$���G  �$����  �z����      C  , ,  ������  �����G  �r���G  �r����  ������      C  , ,  ��  �  ��    �P    �P  �  ��  �      C  , ,  ��  �  ��    ��    ��  �  ��  �      C  , ,  �B  �  �B    ��    ��  �  �B  �      C  , ,  ��  �  ��    �:    �:  �  ��  �      C  , ,  ��  �  ��    ��    ��  �  ��  �      C  , ,  �,  �  �,    ��    ��  �  �,  �      C  , ,  �z  �  �z    �$    �$  �  �z  �      C  , ,  ��  �  ��    �r    �r  �  ��  �      C  , ,  �1  �  �1    ��    ��  �  �1  �      C  , ,  �  �  �    �)    �)  �  �  �      C  , ,  �
     �
   �  ��   �  ��     �
         C  , ,  �X     �X   �  �   �  �     �X         C  , ,  ��     ��   �  �P   �  �P     ��         C  , ,  ��     ��   �  ��   �  ��     ��         C  , ,  �B     �B   �  ��   �  ��     �B         C  , ,  ��     ��   �  �:   �  �:     ��         C  , ,  ��     ��   �  ��   �  ��     ��         C  , ,  �,     �,   �  ��   �  ��     �,         C  , ,  �z     �z   �  �$   �  �$     �z         C  , ,  �
  �  �
  O  ��  O  ��  �  �
  �      C  , ,  �X  �  �X  O  �  O  �  �  �X  �      C  , ,  ��  �  ��  O  �P  O  �P  �  ��  �      C  , ,  ��  �  ��  O  ��  O  ��  �  ��  �      C  , ,  �
  =  �
  �  ��  �  ��  =  �
  =      C  , ,  �X  =  �X  �  �  �  �  =  �X  =      C  , ,  ��  =  ��  �  �P  �  �P  =  ��  =      C  , ,  ��  =  ��  �  ��  �  ��  =  ��  =      C  , ,  �B  =  �B  �  ��  �  ��  =  �B  =      C  , ,  ��  =  ��  �  �:  �  �:  =  ��  =      C  , ,  ��  =  ��  �  ��  �  ��  =  ��  =      C  , ,  �,  =  �,  �  ��  �  ��  =  �,  =      C  , ,  �z  =  �z  �  �$  �  �$  =  �z  =      C  , ,  ��  =  ��  �  �r  �  �r  =  ��  =      C  , ,  �B  �  �B  O  ��  O  ��  �  �B  �      C  , ,  ��  �  ��  O  �:  O  �:  �  ��  �      C  , ,  ��  �  ��  O  ��  O  ��  �  ��  �      C  , ,  �,  �  �,  O  ��  O  ��  �  �,  �      C  , ,  �z  �  �z  O  �$  O  �$  �  �z  �      C  , ,  ��  �  ��  O  �r  O  �r  �  ��  �      C  , ,  ��     ��   �  �r   �  �r     ��         C  , ,  �
���5  �
����  ������  �����5  �
���5      C  , ,  �X���5  �X����  �����  ����5  �X���5      C  , ,  �����5  ������  �P����  �P���5  �����5      C  , ,  �����5  ������  ������  �����5  �����5      C  , ,  �B���5  �B����  ������  �����5  �B���5      C  , ,  �����5  ������  �:����  �:���5  �����5      C  , ,  �����5  ������  ������  �����5  �����5      C  , ,  �,���5  �,����  ������  �����5  �,���5      C  , ,  �z���5  �z����  �$����  �$���5  �z���5      C  , ,  �����5  ������  �r����  �r���5  �����5      C  , ,  �
  �  �
    ��    ��  �  �
  �      C  , ,  ��  �  ��    �w    �w  �  ��  �      C  , ,  �  �  �    ��    ��  �  �  �      C  , ,  �i  �  �i    �    �  �  �i  �      C  , ,  ��  �  ��    �a    �a  �  ��  �      C  , ,  �  �  �    ��    ��  �  �  �      C  , ,  �S  �  �S    ��    ��  �  �S  �      C  , ,  ��  �  ��    �K    �K  �  ��  �      C  , ,  ��  �  ��    ��    ��  �  ��  �      C  , ,  �
  m  �
    ��    ��  m  �
  m      C  , ,  �X  m  �X    �    �  m  �X  m      C  , ,  ��  m  ��    �P    �P  m  ��  m      C  , ,  ��  m  ��    ��    ��  m  ��  m      C  , ,  �B  m  �B    ��    ��  m  �B  m      C  , ,  ��  m  ��    �:    �:  m  ��  m      C  , ,  ��  m  ��    ��    ��  m  ��  m      C  , ,  �,  m  �,    ��    ��  m  �,  m      C  , ,  �z  m  �z    �$    �$  m  �z  m      C  , ,  ��  m  ��    �r    �r  m  ��  m      C  , ,  �X  �  �X    �    �  �  �X  �      C  , ,  �
����  �
���G  �����G  ������  �
����      C  , ,  �X����  �X���G  ����G  �����  �X����      C  , ,  �
����  �
���w  �����w  ������  �
����      C  , ,  �X����  �X���w  ����w  �����  �X����      C  , ,  ��  m  ��    �\    �\  m  ��  m      C  , ,  �   m  �     ��    ��  m  �   m      C  , ,  �N  m  �N    ��    ��  m  �N  m      C  , ,  ��  m  ��    �F    �F  m  ��  m      C  , ,  ��  m  ��    ��    ��  m  ��  m      C  , ,  �8  m  �8    ��    ��  m  �8  m      C  , ,  ��  m  ��    �0    �0  m  ��  m      C  , ,  ��  m  ��    �~    �~  m  ��  m      C  , ,  �d  �  �d  O  �  O  �  �  �d  �      C  , ,  �"  m  �"    ��    ��  m  �"  m      C  , ,  ��  �  ��    �\    �\  �  ��  �      C  , ,  �d     �d   �  �   �  �     �d         C  , ,  ��     ��   �  �\   �  �\     ��         C  , ,  �      �    �  ��   �  ��     �          C  , ,  �N     �N   �  ��   �  ��     �N         C  , ,  ��     ��   �  �F   �  �F     ��         C  , ,  ��     ��   �  ��   �  ��     ��         C  , ,  �8     �8   �  ��   �  ��     �8         C  , ,  ��     ��   �  �0   �  �0     ��         C  , ,  ��     ��   �  �~   �  �~     ��         C  , ,  �d���5  �d����  �����  ����5  �d���5      C  , ,  �����5  ������  �\����  �\���5  �����5      C  , ,  � ���5  � ����  ������  �����5  � ���5      C  , ,  �N���5  �N����  ������  �����5  �N���5      C  , ,  �����5  ������  �F����  �F���5  �����5      C  , ,  �����5  ������  ������  �����5  �����5      C  , ,  �8���5  �8����  ������  �����5  �8���5      C  , ,  �����5  ������  �0����  �0���5  �����5      C  , ,  �����5  ������  �~����  �~���5  �����5      C  , ,  �"���5  �"����  ������  �����5  �"���5      C  , ,  ��  �  ��  O  �\  O  �\  �  ��  �      C  , ,  �   �  �   O  ��  O  ��  �  �   �      C  , ,  �N  �  �N  O  ��  O  ��  �  �N  �      C  , ,  ��  �  ��  O  �F  O  �F  �  ��  �      C  , ,  ��  �  ��  O  ��  O  ��  �  ��  �      C  , ,  �8  �  �8  O  ��  O  ��  �  �8  �      C  , ,  ��  �  ��  O  �0  O  �0  �  ��  �      C  , ,  ��  �  ��  O  �~  O  �~  �  ��  �      C  , ,  �"  �  �"  O  ��  O  ��  �  �"  �      C  , ,  �"     �"   �  ��   �  ��     �"         C  , ,  �d����  �d���G  ����G  �����  �d����      C  , ,  �d  =  �d  �  �  �  �  =  �d  =      C  , ,  ��  =  ��  �  �\  �  �\  =  ��  =      C  , ,  �   =  �   �  ��  �  ��  =  �   =      C  , ,  �N  =  �N  �  ��  �  ��  =  �N  =      C  , ,  ��  =  ��  �  �F  �  �F  =  ��  =      C  , ,  ��  =  ��  �  ��  �  ��  =  ��  =      C  , ,  �8  =  �8  �  ��  �  ��  =  �8  =      C  , ,  ��  =  ��  �  �0  �  �0  =  ��  =      C  , ,  ��  =  ��  �  �~  �  �~  =  ��  =      C  , ,  ������  �����G  �\���G  �\����  ������      C  , ,  � ����  � ���G  �����G  ������  � ����      C  , ,  �N����  �N���G  �����G  ������  �N����      C  , ,  ������  �����G  �F���G  �F����  ������      C  , ,  ������  �����G  �����G  ������  ������      C  , ,  �8����  �8���G  �����G  ������  �8����      C  , ,  ������  �����G  �0���G  �0����  ������      C  , ,  ������  �����G  �~���G  �~����  ������      C  , ,  �"����  �"���G  �����G  ������  �"����      C  , ,  �   �  �     ��    ��  �  �   �      C  , ,  �N  �  �N    ��    ��  �  �N  �      C  , ,  ��  �  ��    �F    �F  �  ��  �      C  , ,  ��  �  ��    ��    ��  �  ��  �      C  , ,  �8  �  �8    ��    ��  �  �8  �      C  , ,  ��  �  ��    �0    �0  �  ��  �      C  , ,  ��  �  ��    �~    �~  �  ��  �      C  , ,  �"  �  �"    ��    ��  �  �"  �      C  , ,  �=  �  �=    ��    ��  �  �=  �      C  , ,  ��  �  ��    �5    �5  �  ��  �      C  , ,  ��  �  ��    ��    ��  �  ��  �      C  , ,  �'  �  �'    ��    ��  �  �'  �      C  , ,  �"  =  �"  �  ��  �  ��  =  �"  =      C  , ,  �u  �  �u    �    �  �  �u  �      C  , ,  ��  �  ��    �m    �m  �  ��  �      C  , ,  �  �  �    ��    ��  �  �  �      C  , ,  �_  �  �_    �	    �	  �  �_  �      C  , ,  ��  �  ��    �W    �W  �  ��  �      C  , ,  ��  �  ��    ��    ��  �  ��  �      C  , ,  �I  �  �I    ��    ��  �  �I  �      C  , ,  �d  �  �d    �    �  �  �d  �      C  , ,  �d  m  �d    �    �  m  �d  m      C  , ,  �d����  �d���w  ����w  �����  �d����      C  , ,  ������  �����w  �\���w  �\����  ������      C  , ,  � ����  � ���w  �����w  ������  � ����      C  , ,  �N����  �N���w  �����w  ������  �N����      C  , ,  ������  �����w  �F���w  �F����  ������      C  , ,  ������  �����w  �����w  ������  ������      C  , ,  �8����  �8���w  �����w  ������  �8����      C  , ,  ������  �����w  �0���w  �0����  ������      C  , ,  ������  �����w  �~���w  �~����  ������      C  , ,  �"����  �"���w  �����w  ������  �"����      C  , ,  ������  �����  �����  ������  ������      C  , ,  ������  �����u  �����u  ������  ������      C  , ,  �����  ����  �����  ������  �����      C  , ,  ����  ����1  �����1  �����  ����      C  , ,  ����  �����  ������  �����  ����      C  , ,  ����  ����a  �����a  �����  ����      C  , ,  ����O  �����  ������  �����O  ����O      C  , ,  �����  ����  �����  ������  �����      C  , ,  ����  ����)  �����)  �����  ����      C  , ,  ����  �����  ������  �����  ����      C  , ,  ���ݛ  ����E  �����E  ����ݛ  ���ݛ      C  , ,  �@����  �@����  ������  ������  �@����      C  , ,  ������  ������  �R����  �R����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �x����  �x����  �"����  �"����  �x����      C  , ,  ������  ������  ������  ������  ������      C  , ,  �H����  �H����  ������  ������  �H����      C  , ,  ������  ������  �Z����  �Z����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �����/  ������  �B����  �B���/  �����/      C  , ,  � ���/  � ����  ������  �����/  � ���/      C  , ,  �h���/  �h����  �����  ����/  �h���/      C  , ,  �����/  ������  �z����  �z���/  �����/      C  , ,  �8���/  �8����  ������  �����/  �8���/      C  , ,  �����/  ������  �J����  �J���/  �����/      C  , ,  ����/  �����  ������  �����/  ����/      C  , ,  �p���/  �p����  �����  ����/  �p���/      C  , ,  �����/  ������  ������  �����/  �����/      C  , ,  �@���/  �@����  ������  �����/  �@���/      C  , ,  �����/  ������  �R����  �R���/  �����/      C  , ,  ����/  �����  ������  �����/  ����/      C  , ,  �x���/  �x����  �"����  �"���/  �x���/      C  , ,  �����/  ������  ������  �����/  �����/      C  , ,  �H���/  �H����  ������  �����/  �H���/      C  , ,  �����/  ������  �Z����  �Z���/  �����/      C  , ,  ����/  �����  ������  �����/  ����/      C  , ,  ������  ������  �B����  �B����  ������      C  , ,  �d����  �d���  ����  �����  �d����      C  , ,  ������  �����  �\���  �\����  ������      C  , ,  � ����  � ���  �����  ������  � ����      C  , ,  �N����  �N���  �����  ������  �N����      C  , ,  ������  �����  �F���  �F����  ������      C  , ,  ������  �����  �����  ������  ������      C  , ,  �8����  �8���  �����  ������  �8����      C  , ,  ������  �����  �0���  �0����  ������      C  , ,  ������  �����  �~���  �~����  ������      C  , ,  �"����  �"���  �����  ������  �"����      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  �d���  �d���1  ����1  ����  �d���      C  , ,  �����  �����1  �\���1  �\���  �����      C  , ,  � ���  � ���1  �����1  �����  � ���      C  , ,  �N���  �N���1  �����1  �����  �N���      C  , ,  �����  �����1  �F���1  �F���  �����      C  , ,  �����  �����1  �����1  �����  �����      C  , ,  �8���  �8���1  �����1  �����  �8���      C  , ,  �����  �����1  �0���1  �0���  �����      C  , ,  �����  �����1  �~���1  �~���  �����      C  , ,  �"���  �"���1  �����1  �����  �"���      C  , ,  �h����  �h����  �����  �����  �h����      C  , ,  ������  ������  �z����  �z����  ������      C  , ,  �8����  �8����  ������  ������  �8����      C  , ,  ������  ������  �J����  �J����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �p����  �p����  �����  �����  �p����      C  , ,  ������  ������  ������  ������  ������      C  , ,  ������  �����I  �B���I  �B����  ������      C  , ,  � ����  � ���I  �����I  ������  � ����      C  , ,  �h����  �h���I  ����I  �����  �h����      C  , ,  ������  �����I  �z���I  �z����  ������      C  , ,  �8����  �8���I  �����I  ������  �8����      C  , ,  ������  �����I  �J���I  �J����  ������      C  , ,  �����  ����I  �����I  ������  �����      C  , ,  �p����  �p���I  ����I  �����  �p����      C  , ,  ������  �����I  �����I  ������  ������      C  , ,  �@����  �@���I  �����I  ������  �@����      C  , ,  ������  �����I  �R���I  �R����  ������      C  , ,  �����  ����I  �����I  ������  �����      C  , ,  �x����  �x���I  �"���I  �"����  �x����      C  , ,  ������  �����I  �����I  ������  ������      C  , ,  �H����  �H���I  �����I  ������  �H����      C  , ,  ������  �����I  �Z���I  �Z����  ������      C  , ,  �����  ����I  �����I  ������  �����      C  , ,  � ���/  � ����  ������  �����/  � ���/      C  , ,  �����/  ������  �2����  �2���/  �����/      C  , ,  �����/  ������  ������  �����/  �����/      C  , ,  �X���/  �X����  �����  ����/  �X���/      C  , ,  �����/  ������  �j����  �j���/  �����/      C  , ,  �(���/  �(����  ������  �����/  �(���/      C  , ,  �����/  ������  �:����  �:���/  �����/      C  , ,  �
���  �
���1  �����1  �����  �
���      C  , ,  �X���  �X���1  ����1  ����  �X���      C  , ,  �����  �����1  �P���1  �P���  �����      C  , ,  �����  �����1  �����1  �����  �����      C  , ,  �B���  �B���1  �����1  �����  �B���      C  , ,  �����  �����1  �:���1  �:���  �����      C  , ,  �����  �����1  �����1  �����  �����      C  , ,  �,���  �,���1  �����1  �����  �,���      C  , ,  �z���  �z���1  �$���1  �$���  �z���      C  , ,  �����  �����1  �r���1  �r���  �����      C  , ,  �����/  ������  ������  �����/  �����/      C  , ,  �`���/  �`����  �
����  �
���/  �`���/      C  , ,  �����/  ������  �r����  �r���/  �����/      C  , ,  �0���/  �0����  ������  �����/  �0���/      C  , ,  �P����  �P����  ������  ������  �P����      C  , ,  ������  ������  �b����  �b����  ������      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  ������  ������  �2����  �2����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �X����  �X����  �����  �����  �X����      C  , ,  ������  ������  �j����  �j����  ������      C  , ,  �(����  �(����  ������  ������  �(����      C  , ,  ������  ������  �:����  �:����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �`����  �`����  �
����  �
����  �`����      C  , ,  ������  ������  �r����  �r����  ������      C  , ,  �0����  �0����  ������  ������  �0����      C  , ,  ������  ������  �Z����  �Z����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  ������  ������  �*����  �*����  ������      C  , ,  ������  �����I  �Z���I  �Z����  ������      C  , ,  �����  ����I  �����I  ������  �����      C  , ,  ������  �����I  �*���I  �*����  ������      C  , ,  ������  �����I  �����I  ������  ������      C  , ,  �P����  �P���I  �����I  ������  �P����      C  , ,  ������  �����I  �b���I  �b����  ������      C  , ,  � ����  � ���I  �����I  ������  � ����      C  , ,  ������  �����I  �2���I  �2����  ������      C  , ,  ������  �����I  �����I  ������  ������      C  , ,  �X����  �X���I  ����I  �����  �X����      C  , ,  ������  �����I  �j���I  �j����  ������      C  , ,  �(����  �(���I  �����I  ������  �(����      C  , ,  ������  �����I  �:���I  �:����  ������      C  , ,  ������  �����I  �����I  ������  ������      C  , ,  �`����  �`���I  �
���I  �
����  �`����      C  , ,  ������  �����I  �r���I  �r����  ������      C  , ,  �0����  �0���I  �����I  ������  �0����      C  , ,  ������  ������  ������  ������  ������      C  , ,  �����/  ������  �Z����  �Z���/  �����/      C  , ,  ����/  �����  ������  �����/  ����/      C  , ,  �
����  �
���  �����  ������  �
����      C  , ,  �X����  �X���  ����  �����  �X����      C  , ,  ������  �����  �P���  �P����  ������      C  , ,  ������  �����  �����  ������  ������      C  , ,  �B����  �B���  �����  ������  �B����      C  , ,  ������  �����  �:���  �:����  ������      C  , ,  ������  �����  �����  ������  ������      C  , ,  �,����  �,���  �����  ������  �,����      C  , ,  �z����  �z���  �$���  �$����  �z����      C  , ,  ������  �����  �r���  �r����  ������      C  , ,  �����/  ������  �*����  �*���/  �����/      C  , ,  �����/  ������  ������  �����/  �����/      C  , ,  �P���/  �P����  ������  �����/  �P���/      C  , ,  �����/  ������  �b����  �b���/  �����/      C  , ,  �����  ������  ������  �����  �����      C  , ,  �
���  �
���)  �����)  �����  �
���      C  , ,  �X���  �X���)  ����)  ����  �X���      C  , ,  �����  �����)  �P���)  �P���  �����      C  , ,  �����  �����)  �����)  �����  �����      C  , ,  �B���  �B���)  �����)  �����  �B���      C  , ,  �����  �����)  �:���)  �:���  �����      C  , ,  �����  �����)  �����)  �����  �����      C  , ,  �,���  �,���)  �����)  �����  �,���      C  , ,  �z���  �z���)  �$���)  �$���  �z���      C  , ,  �����  �����)  �r���)  �r���  �����      C  , ,  �B���  �B����  ������  �����  �B���      C  , ,  �
���  �
����  ������  �����  �
���      C  , ,  �X���  �X����  �����  ����  �X���      C  , ,  �����  ������  �P����  �P���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �B���  �B����  ������  �����  �B���      C  , ,  �����  ������  �:����  �:���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �,���  �,����  ������  �����  �,���      C  , ,  �z���  �z����  �$����  �$���  �z���      C  , ,  �����  ������  �r����  �r���  �����      C  , ,  �����  ������  �:����  �:���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �1����  �1���  �����  ������  �1����      C  , ,  �����  ����  �)���  �)����  �����      C  , ,  ������  �����  �w���  �w����  ������      C  , ,  �����  ����  �����  ������  �����      C  , ,  �i����  �i���  ����  �����  �i����      C  , ,  ������  �����  �a���  �a����  ������      C  , ,  �����  ����  �����  ������  �����      C  , ,  �S����  �S���  �����  ������  �S����      C  , ,  ������  �����  �K���  �K����  ������      C  , ,  ������  �����  �����  ������  ������      C  , ,  �,���  �,����  ������  �����  �,���      C  , ,  �1����  �1���u  �����u  ������  �1����      C  , ,  �����  ����u  �)���u  �)����  �����      C  , ,  ������  �����u  �w���u  �w����  ������      C  , ,  �����  ����u  �����u  ������  �����      C  , ,  �i����  �i���u  ����u  �����  �i����      C  , ,  ������  �����u  �a���u  �a����  ������      C  , ,  �����  ����u  �����u  ������  �����      C  , ,  �S����  �S���u  �����u  ������  �S����      C  , ,  ������  �����u  �K���u  �K����  ������      C  , ,  ������  �����u  �����u  ������  ������      C  , ,  �
��ݛ  �
���E  �����E  ����ݛ  �
��ݛ      C  , ,  �X��ݛ  �X���E  ����E  ���ݛ  �X��ݛ      C  , ,  ����ݛ  �����E  �P���E  �P��ݛ  ����ݛ      C  , ,  ����ݛ  �����E  �����E  ����ݛ  ����ݛ      C  , ,  �B��ݛ  �B���E  �����E  ����ݛ  �B��ݛ      C  , ,  ����ݛ  �����E  �:���E  �:��ݛ  ����ݛ      C  , ,  ����ݛ  �����E  �����E  ����ݛ  ����ݛ      C  , ,  �,��ݛ  �,���E  �����E  ����ݛ  �,��ݛ      C  , ,  �z��ݛ  �z���E  �$���E  �$��ݛ  �z��ݛ      C  , ,  ����ݛ  �����E  �r���E  �r��ݛ  ����ݛ      C  , ,  �z���  �z����  �$����  �$���  �z���      C  , ,  �����  ������  �r����  �r���  �����      C  , ,  �
���  �
����  ������  �����  �
���      C  , ,  �
���  �
���a  �����a  �����  �
���      C  , ,  �X���  �X���a  ����a  ����  �X���      C  , ,  �����  �����a  �P���a  �P���  �����      C  , ,  �����  �����a  �����a  �����  �����      C  , ,  �B���  �B���a  �����a  �����  �B���      C  , ,  �����  �����a  �:���a  �:���  �����      C  , ,  �����  �����a  �����a  �����  �����      C  , ,  �,���  �,���a  �����a  �����  �,���      C  , ,  �z���  �z���a  �$���a  �$���  �z���      C  , ,  �����  �����a  �r���a  �r���  �����      C  , ,  �X���  �X����  �����  ����  �X���      C  , ,  �
���O  �
����  ������  �����O  �
���O      C  , ,  �X���O  �X����  �����  ����O  �X���O      C  , ,  �����O  ������  �P����  �P���O  �����O      C  , ,  �����O  ������  ������  �����O  �����O      C  , ,  �B���O  �B����  ������  �����O  �B���O      C  , ,  �����O  ������  �:����  �:���O  �����O      C  , ,  �����O  ������  ������  �����O  �����O      C  , ,  �,���O  �,����  ������  �����O  �,���O      C  , ,  �z���O  �z����  �$����  �$���O  �z���O      C  , ,  �����O  ������  �r����  �r���O  �����O      C  , ,  �����  ������  �P����  �P���  �����      C  , ,  �
����  �
���  �����  ������  �
����      C  , ,  �X����  �X���  ����  �����  �X����      C  , ,  ������  �����  �P���  �P����  ������      C  , ,  ������  �����  �����  ������  ������      C  , ,  �B����  �B���  �����  ������  �B����      C  , ,  ������  �����  �:���  �:����  ������      C  , ,  ������  �����  �����  ������  ������      C  , ,  �,����  �,���  �����  ������  �,����      C  , ,  �z����  �z���  �$���  �$����  �z����      C  , ,  ������  �����  �r���  �r����  ������      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �d����  �d���  ����  �����  �d����      C  , ,  ������  �����  �\���  �\����  ������      C  , ,  � ����  � ���  �����  ������  � ����      C  , ,  �=����  �=���  �����  ������  �=����      C  , ,  ������  �����  �5���  �5����  ������      C  , ,  ������  �����  �����  ������  ������      C  , ,  �'����  �'���  �����  ������  �'����      C  , ,  �u����  �u���  ����  �����  �u����      C  , ,  ������  �����  �m���  �m����  ������      C  , ,  �����  ����  �����  ������  �����      C  , ,  �_����  �_���  �	���  �	����  �_����      C  , ,  ������  �����  �W���  �W����  ������      C  , ,  ������  �����  �����  ������  ������      C  , ,  �I����  �I���  �����  ������  �I����      C  , ,  �N����  �N���  �����  ������  �N����      C  , ,  ������  �����  �F���  �F����  ������      C  , ,  ������  �����  �����  ������  ������      C  , ,  �8����  �8���  �����  ������  �8����      C  , ,  ������  �����  �0���  �0����  ������      C  , ,  ������  �����  �~���  �~����  ������      C  , ,  �"����  �"���  �����  ������  �"����      C  , ,  �N���  �N����  ������  �����  �N���      C  , ,  �����  ������  �F����  �F���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �8���  �8����  ������  �����  �8���      C  , ,  �=����  �=���u  �����u  ������  �=����      C  , ,  ������  �����u  �5���u  �5����  ������      C  , ,  ������  �����u  �����u  ������  ������      C  , ,  �'����  �'���u  �����u  ������  �'����      C  , ,  �u����  �u���u  ����u  �����  �u����      C  , ,  ������  �����u  �m���u  �m����  ������      C  , ,  �����  ����u  �����u  ������  �����      C  , ,  �_����  �_���u  �	���u  �	����  �_����      C  , ,  ������  �����u  �W���u  �W����  ������      C  , ,  ������  �����u  �����u  ������  ������      C  , ,  �I����  �I���u  �����u  ������  �I����      C  , ,  �����  ������  �0����  �0���  �����      C  , ,  �����  ������  �~����  �~���  �����      C  , ,  �"���  �"����  ������  �����  �"���      C  , ,  �d���  �d����  �����  ����  �d���      C  , ,  �d���  �d���a  ����a  ����  �d���      C  , ,  �d���O  �d����  �����  ����O  �d���O      C  , ,  �����O  ������  �\����  �\���O  �����O      C  , ,  �d���  �d���)  ����)  ����  �d���      C  , ,  �����  �����)  �\���)  �\���  �����      C  , ,  � ���  � ���)  �����)  �����  � ���      C  , ,  �N���  �N���)  �����)  �����  �N���      C  , ,  �d��ݛ  �d���E  ����E  ���ݛ  �d��ݛ      C  , ,  ����ݛ  �����E  �\���E  �\��ݛ  ����ݛ      C  , ,  � ��ݛ  � ���E  �����E  ����ݛ  � ��ݛ      C  , ,  �N��ݛ  �N���E  �����E  ����ݛ  �N��ݛ      C  , ,  ����ݛ  �����E  �F���E  �F��ݛ  ����ݛ      C  , ,  ����ݛ  �����E  �����E  ����ݛ  ����ݛ      C  , ,  �8��ݛ  �8���E  �����E  ����ݛ  �8��ݛ      C  , ,  ����ݛ  �����E  �0���E  �0��ݛ  ����ݛ      C  , ,  ����ݛ  �����E  �~���E  �~��ݛ  ����ݛ      C  , ,  �"��ݛ  �"���E  �����E  ����ݛ  �"��ݛ      C  , ,  �����  �����)  �F���)  �F���  �����      C  , ,  �����  �����)  �����)  �����  �����      C  , ,  �8���  �8���)  �����)  �����  �8���      C  , ,  �����  �����)  �0���)  �0���  �����      C  , ,  �����  �����)  �~���)  �~���  �����      C  , ,  �"���  �"���)  �����)  �����  �"���      C  , ,  � ���O  � ����  ������  �����O  � ���O      C  , ,  �N���O  �N����  ������  �����O  �N���O      C  , ,  �����O  ������  �F����  �F���O  �����O      C  , ,  �����O  ������  ������  �����O  �����O      C  , ,  �8���O  �8����  ������  �����O  �8���O      C  , ,  �����O  ������  �0����  �0���O  �����O      C  , ,  �����O  ������  �~����  �~���O  �����O      C  , ,  �"���O  �"����  ������  �����O  �"���O      C  , ,  �����  �����a  �\���a  �\���  �����      C  , ,  � ���  � ���a  �����a  �����  � ���      C  , ,  �N���  �N���a  �����a  �����  �N���      C  , ,  �d���  �d����  �����  ����  �d���      C  , ,  �����  ������  �\����  �\���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �N���  �N����  ������  �����  �N���      C  , ,  �����  ������  �F����  �F���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �8���  �8����  ������  �����  �8���      C  , ,  �����  ������  �0����  �0���  �����      C  , ,  �����  ������  �~����  �~���  �����      C  , ,  �"���  �"����  ������  �����  �"���      C  , ,  �����  �����a  �F���a  �F���  �����      C  , ,  �����  �����a  �����a  �����  �����      C  , ,  �8���  �8���a  �����a  �����  �8���      C  , ,  �����  �����a  �0���a  �0���  �����      C  , ,  �����  �����a  �~���a  �~���  �����      C  , ,  �"���  �"���a  �����a  �����  �"���      C  , ,  �����  ������  �\����  �\���  �����      C  , ,  r`����  r`����  s
����  s
����  r`����      C  , ,  r`���/  r`����  s
����  s
���/  r`���/      C  , ,  r`����  r`���I  s
���I  s
����  r`����      C  , ,  y����  y����1  zD���1  zD���  y����      C  , ,  {����  {����1  |����1  |����  {����      C  , ,  ~6���  ~6���1  ~����1  ~����  ~6���      C  , ,  �����  �����1  �.���1  �.���  �����      C  , ,  �����  �����1  �|���1  �|���  �����      C  , ,  � ���  � ���1  �����1  �����  � ���      C  , ,  �n���  �n���1  ����1  ����  �n���      C  , ,  �����  �����1  �f���1  �f���  �����      C  , ,  ������  ������  �R����  �R����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �x����  �x����  �"����  �"����  �x����      C  , ,  ������  ������  ������  ������  ������      C  , ,  �H����  �H����  ������  ������  �H����      C  , ,  r����  r����1  sZ���1  sZ���  r����      C  , ,  s�����  s�����  tr����  tr����  s�����      C  , ,  u0����  u0����  u�����  u�����  u0����      C  , ,  v�����  v�����  wB����  wB����  v�����      C  , ,  x ����  x ����  x�����  x�����  x ����      C  , ,  yh����  yh����  z����  z����  yh����      C  , ,  z�����  z�����  {z����  {z����  z�����      C  , ,  |8����  |8����  |�����  |�����  |8����      C  , ,  }�����  }�����  ~J����  ~J����  }�����      C  , ,  ����  ����  �����  �����  ����      C  , ,  �p����  �p����  �����  �����  �p����      C  , ,  ������  ������  ������  ������  ������      C  , ,  r�����  r����  sZ���  sZ����  r�����      C  , ,  t�����  t����  u����  u�����  t�����      C  , ,  wL����  wL���  w����  w�����  wL����      C  , ,  y�����  y����  zD���  zD����  y�����      C  , ,  {�����  {����  |����  |�����  {�����      C  , ,  ~6����  ~6���  ~����  ~�����  ~6����      C  , ,  ������  �����  �.���  �.����  ������      C  , ,  ������  �����  �|���  �|����  ������      C  , ,  � ����  � ���  �����  ������  � ����      C  , ,  �n����  �n���  ����  �����  �n����      C  , ,  ������  �����  �f���  �f����  ������      C  , ,  t����  t����1  u����1  u����  t����      C  , ,  s����/  s�����  tr����  tr���/  s����/      C  , ,  u0���/  u0����  u�����  u����/  u0���/      C  , ,  v����/  v�����  wB����  wB���/  v����/      C  , ,  x ���/  x ����  x�����  x����/  x ���/      C  , ,  yh���/  yh����  z����  z���/  yh���/      C  , ,  z����/  z�����  {z����  {z���/  z����/      C  , ,  wL���  wL���1  w����1  w����  wL���      C  , ,  s�����  s����I  tr���I  tr����  s�����      C  , ,  u0����  u0���I  u����I  u�����  u0����      C  , ,  v�����  v����I  wB���I  wB����  v�����      C  , ,  x ����  x ���I  x����I  x�����  x ����      C  , ,  yh����  yh���I  z���I  z����  yh����      C  , ,  z�����  z����I  {z���I  {z����  z�����      C  , ,  |8����  |8���I  |����I  |�����  |8����      C  , ,  }�����  }����I  ~J���I  ~J����  }�����      C  , ,  ����  ���I  ����I  �����  ����      C  , ,  �p����  �p���I  ����I  �����  �p����      C  , ,  ������  �����I  �����I  ������  ������      C  , ,  �@����  �@���I  �����I  ������  �@����      C  , ,  ������  �����I  �R���I  �R����  ������      C  , ,  �����  ����I  �����I  ������  �����      C  , ,  �x����  �x���I  �"���I  �"����  �x����      C  , ,  ������  �����I  �����I  ������  ������      C  , ,  �H����  �H���I  �����I  ������  �H����      C  , ,  |8���/  |8����  |�����  |����/  |8���/      C  , ,  }����/  }�����  ~J����  ~J���/  }����/      C  , ,  ���/  ����  �����  ����/  ���/      C  , ,  �p���/  �p����  �����  ����/  �p���/      C  , ,  �����/  ������  ������  �����/  �����/      C  , ,  �@���/  �@����  ������  �����/  �@���/      C  , ,  �����/  ������  �R����  �R���/  �����/      C  , ,  ����/  �����  ������  �����/  ����/      C  , ,  �x���/  �x����  �"����  �"���/  �x���/      C  , ,  �����/  ������  ������  �����/  �����/      C  , ,  �H���/  �H����  ������  �����/  �H���/      C  , ,  �@����  �@����  ������  ������  �@����      C  , ,  dP����  dP���I  d����I  d�����  dP����      C  , ,  e�����  e����I  fb���I  fb����  e�����      C  , ,  g ����  g ���I  g����I  g�����  g ����      C  , ,  h�����  h����I  i2���I  i2����  h�����      C  , ,  i�����  i����I  j����I  j�����  i�����      C  , ,  kX����  kX���I  l���I  l����  kX����      C  , ,  l�����  l����I  mj���I  mj����  l�����      C  , ,  n(����  n(���I  n����I  n�����  n(����      C  , ,  o�����  o����I  p:���I  p:����  o�����      C  , ,  p�����  p����I  q����I  q�����  p�����      C  , ,  `@����  `@���  `����  `�����  `@����      C  , ,  b�����  b����  c8���  c8����  b�����      C  , ,  d�����  d����  e����  e�����  d�����      C  , ,  g*����  g*���  g����  g�����  g*����      C  , ,  ix����  ix���  j"���  j"����  ix����      C  , ,  k�����  k����  lp���  lp����  k�����      C  , ,  n����  n���  n����  n�����  n����      C  , ,  pb����  pb���  q���  q����  pb����      C  , ,  o�����  o�����  p:����  p:����  o�����      C  , ,  p�����  p�����  q�����  q�����  p�����      C  , ,  ^�����  ^����I  _Z���I  _Z����  ^�����      C  , ,  ]H���/  ]H����  ]�����  ]����/  ]H���/      C  , ,  ^����/  ^�����  _Z����  _Z���/  ^����/      C  , ,  `���/  `����  `�����  `����/  `���/      C  , ,  a����/  a�����  b*����  b*���/  a����/      C  , ,  b����/  b�����  c�����  c����/  b����/      C  , ,  dP���/  dP����  d�����  d����/  dP���/      C  , ,  e����/  e�����  fb����  fb���/  e����/      C  , ,  g ���/  g ����  g�����  g����/  g ���/      C  , ,  o����/  o�����  p:����  p:���/  o����/      C  , ,  p����/  p�����  q�����  q����/  p����/      C  , ,  h����/  h�����  i2����  i2���/  h����/      C  , ,  i����/  i�����  j�����  j����/  i����/      C  , ,  kX���/  kX����  l����  l���/  kX���/      C  , ,  l����/  l�����  mj����  mj���/  l����/      C  , ,  n(���/  n(����  n�����  n����/  n(���/      C  , ,  `����  `���I  `����I  `�����  `����      C  , ,  ]�����  ]����  ^����  ^�����  ]�����      C  , ,  a�����  a����I  b*���I  b*����  a�����      C  , ,  b�����  b����I  c����I  c�����  b�����      C  , ,  ]����  ]����1  ^����1  ^����  ]����      C  , ,  `@���  `@���1  `����1  `����  `@���      C  , ,  b����  b����1  c8���1  c8���  b����      C  , ,  d����  d����1  e����1  e����  d����      C  , ,  g*���  g*���1  g����1  g����  g*���      C  , ,  ix���  ix���1  j"���1  j"���  ix���      C  , ,  k����  k����1  lp���1  lp���  k����      C  , ,  n���  n���1  n����1  n����  n���      C  , ,  pb���  pb���1  q���1  q���  pb���      C  , ,  ]H����  ]H���I  ]����I  ]�����  ]H����      C  , ,  ]H����  ]H����  ]�����  ]�����  ]H����      C  , ,  ^�����  ^�����  _Z����  _Z����  ^�����      C  , ,  `����  `����  `�����  `�����  `����      C  , ,  a�����  a�����  b*����  b*����  a�����      C  , ,  b�����  b�����  c�����  c�����  b�����      C  , ,  dP����  dP����  d�����  d�����  dP����      C  , ,  e�����  e�����  fb����  fb����  e�����      C  , ,  g ����  g ����  g�����  g�����  g ����      C  , ,  h�����  h�����  i2����  i2����  h�����      C  , ,  i�����  i�����  j�����  j�����  i�����      C  , ,  kX����  kX����  l����  l����  kX����      C  , ,  l�����  l�����  mj����  mj����  l�����      C  , ,  n(����  n(����  n�����  n�����  n(����      C  , ,  ]����O  ]�����  ^�����  ^����O  ]����O      C  , ,  `@���O  `@����  `�����  `����O  `@���O      C  , ,  b����O  b�����  c8����  c8���O  b����O      C  , ,  d����O  d�����  e�����  e����O  d����O      C  , ,  g*���O  g*����  g�����  g����O  g*���O      C  , ,  ix���O  ix����  j"����  j"���O  ix���O      C  , ,  k����O  k�����  lp����  lp���O  k����O      C  , ,  n���O  n����  n�����  n����O  n���O      C  , ,  pb���O  pb����  q����  q���O  pb���O      C  , ,  c�����  c����  d_���  d_����  c�����      C  , ,  f����  f���  f����  f�����  f����      C  , ,  hQ����  hQ���  h����  h�����  hQ����      C  , ,  j�����  j����  kI���  kI����  j�����      C  , ,  l�����  l����  m����  m�����  l�����      C  , ,  o;����  o;���  o����  o�����  o;����      C  , ,  q�����  q����  r3���  r3����  q�����      C  , ,  ]����  ]�����  ^�����  ^����  ]����      C  , ,  `@���  `@����  `�����  `����  `@���      C  , ,  b����  b�����  c8����  c8���  b����      C  , ,  d����  d�����  e�����  e����  d����      C  , ,  g*���  g*����  g�����  g����  g*���      C  , ,  ix���  ix����  j"����  j"���  ix���      C  , ,  k����  k�����  lp����  lp���  k����      C  , ,  n���  n����  n�����  n����  n���      C  , ,  pb���  pb����  q����  q���  pb���      C  , ,  ]����  ]�����  ^�����  ^����  ]����      C  , ,  ]����  ]����a  ^����a  ^����  ]����      C  , ,  `@���  `@���a  `����a  `����  `@���      C  , ,  b����  b����a  c8���a  c8���  b����      C  , ,  d����  d����a  e����a  e����  d����      C  , ,  g*���  g*���a  g����a  g����  g*���      C  , ,  ix���  ix���a  j"���a  j"���  ix���      C  , ,  k����  k����a  lp���a  lp���  k����      C  , ,  n���  n���a  n����a  n����  n���      C  , ,  pb���  pb���a  q���a  q���  pb���      C  , ,  _����  _���u  _����u  _�����  _����      C  , ,  ag����  ag���u  b���u  b����  ag����      C  , ,  c�����  c����u  d_���u  d_����  c�����      C  , ,  f����  f���u  f����u  f�����  f����      C  , ,  hQ����  hQ���u  h����u  h�����  hQ����      C  , ,  j�����  j����u  kI���u  kI����  j�����      C  , ,  l�����  l����u  m����u  m�����  l�����      C  , ,  o;����  o;���u  o����u  o�����  o;����      C  , ,  q�����  q����u  r3���u  r3����  q�����      C  , ,  `@���  `@����  `�����  `����  `@���      C  , ,  b����  b�����  c8����  c8���  b����      C  , ,  d����  d�����  e�����  e����  d����      C  , ,  g*���  g*����  g�����  g����  g*���      C  , ,  ix���  ix����  j"����  j"���  ix���      C  , ,  k����  k�����  lp����  lp���  k����      C  , ,  n���  n����  n�����  n����  n���      C  , ,  pb���  pb����  q����  q���  pb���      C  , ,  pb����  pb���  q���  q����  pb����      C  , ,  n����  n���  n����  n�����  n����      C  , ,  ]����  ]����)  ^����)  ^����  ]����      C  , ,  `@���  `@���)  `����)  `����  `@���      C  , ,  b����  b����)  c8���)  c8���  b����      C  , ,  d����  d����)  e����)  e����  d����      C  , ,  ]���ݛ  ]����E  ^����E  ^���ݛ  ]���ݛ      C  , ,  `@��ݛ  `@���E  `����E  `���ݛ  `@��ݛ      C  , ,  ]�����  ]����  ^����  ^�����  ]�����      C  , ,  `@����  `@���  `����  `�����  `@����      C  , ,  b�����  b����  c8���  c8����  b�����      C  , ,  d�����  d����  e����  e�����  d�����      C  , ,  g*����  g*���  g����  g�����  g*����      C  , ,  ix����  ix���  j"���  j"����  ix����      C  , ,  k�����  k����  lp���  lp����  k�����      C  , ,  b���ݛ  b����E  c8���E  c8��ݛ  b���ݛ      C  , ,  d���ݛ  d����E  e����E  e���ݛ  d���ݛ      C  , ,  g*��ݛ  g*���E  g����E  g���ݛ  g*��ݛ      C  , ,  ix��ݛ  ix���E  j"���E  j"��ݛ  ix��ݛ      C  , ,  k���ݛ  k����E  lp���E  lp��ݛ  k���ݛ      C  , ,  n��ݛ  n���E  n����E  n���ݛ  n��ݛ      C  , ,  pb��ݛ  pb���E  q���E  q��ݛ  pb��ݛ      C  , ,  g*���  g*���)  g����)  g����  g*���      C  , ,  ix���  ix���)  j"���)  j"���  ix���      C  , ,  k����  k����)  lp���)  lp���  k����      C  , ,  n���  n���)  n����)  n����  n���      C  , ,  pb���  pb���)  q���)  q���  pb���      C  , ,  _����  _���  _����  _�����  _����      C  , ,  ag����  ag���  b���  b����  ag����      C  , ,  ������  �����  �?���  �?����  ������      C  , ,  t�����  t����  u����  u�����  t�����      C  , ,  wL����  wL���  w����  w�����  wL����      C  , ,  y�����  y����  zD���  zD����  y�����      C  , ,  r����  r�����  sZ����  sZ���  r����      C  , ,  t����  t�����  u�����  u����  t����      C  , ,  wL���  wL����  w�����  w����  wL���      C  , ,  y����  y�����  zD����  zD���  y����      C  , ,  {����  {�����  |�����  |����  {����      C  , ,  ~6���  ~6����  ~�����  ~����  ~6���      C  , ,  �����  ������  �.����  �.���  �����      C  , ,  �����  ������  �|����  �|���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �n���  �n����  �����  ����  �n���      C  , ,  r����O  r�����  sZ����  sZ���O  r����O      C  , ,  t����O  t�����  u�����  u����O  t����O      C  , ,  wL���O  wL����  w�����  w����O  wL���O      C  , ,  y����O  y�����  zD����  zD���O  y����O      C  , ,  {����O  {�����  |�����  |����O  {����O      C  , ,  �����  ������  �f����  �f���  �����      C  , ,  t����  t�����  u�����  u����  t����      C  , ,  wL���  wL����  w�����  w����  wL���      C  , ,  y����  y�����  zD����  zD���  y����      C  , ,  {����  {�����  |�����  |����  {����      C  , ,  ~6���  ~6����  ~�����  ~����  ~6���      C  , ,  r����  r����a  sZ���a  sZ���  r����      C  , ,  t����  t����a  u����a  u����  t����      C  , ,  wL���  wL���a  w����a  w����  wL���      C  , ,  �����  ������  �.����  �.���  �����      C  , ,  �����  ������  �|����  �|���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �n���  �n����  �����  ����  �n���      C  , ,  �����  ������  �f����  �f���  �����      C  , ,  {�����  {����  |����  |�����  {�����      C  , ,  ~6����  ~6���  ~����  ~�����  ~6����      C  , ,  ������  �����  �.���  �.����  ������      C  , ,  ������  �����  �|���  �|����  ������      C  , ,  s�����  s����u  t����u  t�����  s�����      C  , ,  v%����  v%���u  v����u  v�����  v%����      C  , ,  xs����  xs���u  y���u  y����  xs����      C  , ,  z�����  z����u  {k���u  {k����  z�����      C  , ,  }����  }���u  }����u  }�����  }����      C  , ,  ]����  ]���u  ����u  �����  ]����      C  , ,  ������  �����u  �U���u  �U����  ������      C  , ,  ������  �����u  �����u  ������  ������      C  , ,  �G����  �G���u  �����u  ������  �G����      C  , ,  ������  �����u  �?���u  �?����  ������      C  , ,  y����  y����a  zD���a  zD���  y����      C  , ,  {����  {����a  |����a  |����  {����      C  , ,  ~6���O  ~6����  ~�����  ~����O  ~6���O      C  , ,  �����O  ������  �.����  �.���O  �����O      C  , ,  �����O  ������  �|����  �|���O  �����O      C  , ,  � ���O  � ����  ������  �����O  � ���O      C  , ,  �n���O  �n����  �����  ����O  �n���O      C  , ,  �����O  ������  �f����  �f���O  �����O      C  , ,  ~6���  ~6���a  ~����a  ~����  ~6���      C  , ,  �����  �����a  �.���a  �.���  �����      C  , ,  �����  �����a  �|���a  �|���  �����      C  , ,  � ���  � ���a  �����a  �����  � ���      C  , ,  �n���  �n���a  ����a  ����  �n���      C  , ,  �����  �����a  �f���a  �f���  �����      C  , ,  r����  r����)  sZ���)  sZ���  r����      C  , ,  t����  t����)  u����)  u����  t����      C  , ,  wL���  wL���)  w����)  w����  wL���      C  , ,  y����  y����)  zD���)  zD���  y����      C  , ,  {����  {����)  |����)  |����  {����      C  , ,  ~6���  ~6���)  ~����)  ~����  ~6���      C  , ,  �����  �����)  �.���)  �.���  �����      C  , ,  �����  �����)  �|���)  �|���  �����      C  , ,  � ���  � ���)  �����)  �����  � ���      C  , ,  r����  r�����  sZ����  sZ���  r����      C  , ,  �n���  �n���)  ����)  ����  �n���      C  , ,  �����  �����)  �f���)  �f���  �����      C  , ,  � ����  � ���  �����  ������  � ����      C  , ,  �n����  �n���  ����  �����  �n����      C  , ,  ������  �����  �f���  �f����  ������      C  , ,  r�����  r����  sZ���  sZ����  r�����      C  , ,  s�����  s����  t����  t�����  s�����      C  , ,  v%����  v%���  v����  v�����  v%����      C  , ,  xs����  xs���  y���  y����  xs����      C  , ,  z�����  z����  {k���  {k����  z�����      C  , ,  }����  }���  }����  }�����  }����      C  , ,  ]����  ]���  ����  �����  ]����      C  , ,  ������  �����  �U���  �U����  ������      C  , ,  r���ݛ  r����E  sZ���E  sZ��ݛ  r���ݛ      C  , ,  t���ݛ  t����E  u����E  u���ݛ  t���ݛ      C  , ,  wL��ݛ  wL���E  w����E  w���ݛ  wL��ݛ      C  , ,  y���ݛ  y����E  zD���E  zD��ݛ  y���ݛ      C  , ,  {���ݛ  {����E  |����E  |���ݛ  {���ݛ      C  , ,  ~6��ݛ  ~6���E  ~����E  ~���ݛ  ~6��ݛ      C  , ,  ����ݛ  �����E  �.���E  �.��ݛ  ����ݛ      C  , ,  ����ݛ  �����E  �|���E  �|��ݛ  ����ݛ      C  , ,  � ��ݛ  � ���E  �����E  ����ݛ  � ��ݛ      C  , ,  �n��ݛ  �n���E  ����E  ���ݛ  �n��ݛ      C  , ,  ����ݛ  �����E  �f���E  �f��ݛ  ����ݛ      C  , ,  ������  �����  �����  ������  ������      C  , ,  �G����  �G���  �����  ������  �G����      C  , ,  r`��ϕ  r`���?  s
���?  s
��ϕ  r`��ϕ      C  , ,  r`����  r`��·  s
��·  s
����  r`����      C  , ,  r`���%  r`����  s
����  s
���%  r`���%      C  , ,  t���֓  t����=  u����=  u���֓  t���֓      C  , ,  wL��֓  wL���=  w����=  w���֓  wL��֓      C  , ,  y���֓  y����=  zD���=  zD��֓  y���֓      C  , ,  {���֓  {����=  |����=  |���֓  {���֓      C  , ,  ~6��֓  ~6���=  ~����=  ~���֓  ~6��֓      C  , ,  ����֓  �����=  �.���=  �.��֓  ����֓      C  , ,  ����֓  �����=  �|���=  �|��֓  ����֓      C  , ,  � ��֓  � ���=  �����=  ����֓  � ��֓      C  , ,  �n��֓  �n���=  ����=  ���֓  �n��֓      C  , ,  ����֓  �����=  �f���=  �f��֓  ����֓      C  , ,  r����+  r�����  sZ����  sZ���+  r����+      C  , ,  t����+  t�����  u�����  u����+  t����+      C  , ,  wL���+  wL����  w�����  w����+  wL���+      C  , ,  y����+  y�����  zD����  zD���+  y����+      C  , ,  {����+  {�����  |�����  |����+  {����+      C  , ,  ~6���+  ~6����  ~�����  ~����+  ~6���+      C  , ,  �����+  ������  �.����  �.���+  �����+      C  , ,  �����+  ������  �|����  �|���+  �����+      C  , ,  � ���+  � ����  ������  �����+  � ���+      C  , ,  �n���+  �n����  �����  ����+  �n���+      C  , ,  �����+  ������  �f����  �f���+  �����+      C  , ,  r�����  r����m  sZ���m  sZ����  r�����      C  , ,  t�����  t����m  u����m  u�����  t�����      C  , ,  wL����  wL���m  w����m  w�����  wL����      C  , ,  y�����  y����m  zD���m  zD����  y�����      C  , ,  {�����  {����m  |����m  |�����  {�����      C  , ,  ~6����  ~6���m  ~����m  ~�����  ~6����      C  , ,  ������  �����m  �.���m  �.����  ������      C  , ,  ������  �����m  �|���m  �|����  ������      C  , ,  � ����  � ���m  �����m  ������  � ����      C  , ,  �n����  �n���m  ����m  �����  �n����      C  , ,  ������  �����m  �f���m  �f����  ������      C  , ,  �n����  �n��إ  ���إ  �����  �n����      C  , ,  s���ϕ  s����?  tr���?  tr��ϕ  s���ϕ      C  , ,  u0��ϕ  u0���?  u����?  u���ϕ  u0��ϕ      C  , ,  v���ϕ  v����?  wB���?  wB��ϕ  v���ϕ      C  , ,  x ��ϕ  x ���?  x����?  x���ϕ  x ��ϕ      C  , ,  yh��ϕ  yh���?  z���?  z��ϕ  yh��ϕ      C  , ,  z���ϕ  z����?  {z���?  {z��ϕ  z���ϕ      C  , ,  |8��ϕ  |8���?  |����?  |���ϕ  |8��ϕ      C  , ,  }���ϕ  }����?  ~J���?  ~J��ϕ  }���ϕ      C  , ,  ��ϕ  ���?  ����?  ���ϕ  ��ϕ      C  , ,  �p��ϕ  �p���?  ����?  ���ϕ  �p��ϕ      C  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      C  , ,  �@��ϕ  �@���?  �����?  ����ϕ  �@��ϕ      C  , ,  ����ϕ  �����?  �R���?  �R��ϕ  ����ϕ      C  , ,  ���ϕ  ����?  �����?  ����ϕ  ���ϕ      C  , ,  �x��ϕ  �x���?  �"���?  �"��ϕ  �x��ϕ      C  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      C  , ,  �H��ϕ  �H���?  �����?  ����ϕ  �H��ϕ      C  , ,  ������  ����إ  �f��إ  �f����  ������      C  , ,  r���֓  r����=  sZ���=  sZ��֓  r���֓      C  , ,  r����3  r�����  sZ����  sZ���3  r����3      C  , ,  t����3  t�����  u�����  u����3  t����3      C  , ,  wL���3  wL����  w�����  w����3  wL���3      C  , ,  y����3  y�����  zD����  zD���3  y����3      C  , ,  {����3  {�����  |�����  |����3  {����3      C  , ,  ~6���3  ~6����  ~�����  ~����3  ~6���3      C  , ,  �����3  ������  �.����  �.���3  �����3      C  , ,  �����3  ������  �|����  �|���3  �����3      C  , ,  � ���3  � ����  ������  �����3  � ���3      C  , ,  �n���3  �n����  �����  ����3  �n���3      C  , ,  �����3  ������  �f����  �f���3  �����3      C  , ,  r�����  r����u  sZ���u  sZ����  r�����      C  , ,  t�����  t����u  u����u  u�����  t�����      C  , ,  wL����  wL���u  w����u  w�����  wL����      C  , ,  y�����  y����u  zD���u  zD����  y�����      C  , ,  {�����  {����u  |����u  |�����  {�����      C  , ,  ~6����  ~6���u  ~����u  ~�����  ~6����      C  , ,  ������  �����u  �.���u  �.����  ������      C  , ,  ������  �����u  �|���u  �|����  ������      C  , ,  � ����  � ���u  �����u  ������  � ����      C  , ,  �n����  �n���u  ����u  �����  �n����      C  , ,  ������  �����u  �f���u  �f����  ������      C  , ,  r����c  r����  sZ���  sZ���c  r����c      C  , ,  t����c  t����  u����  u����c  t����c      C  , ,  wL���c  wL���  w����  w����c  wL���c      C  , ,  y����c  y����  zD���  zD���c  y����c      C  , ,  {����c  {����  |����  |����c  {����c      C  , ,  ~6���c  ~6���  ~����  ~����c  ~6���c      C  , ,  �����c  �����  �.���  �.���c  �����c      C  , ,  �����c  �����  �|���  �|���c  �����c      C  , ,  � ���c  � ���  �����  �����c  � ���c      C  , ,  �n���c  �n���  ����  ����c  �n���c      C  , ,  �����c  �����  �f���  �f���c  �����c      C  , ,  r�����  r���إ  sZ��إ  sZ����  r�����      C  , ,  t�����  t���إ  u���إ  u�����  t�����      C  , ,  wL����  wL��إ  w���إ  w�����  wL����      C  , ,  y�����  y���إ  zD��إ  zD����  y�����      C  , ,  {�����  {���إ  |���إ  |�����  {�����      C  , ,  ~6����  ~6��إ  ~���إ  ~�����  ~6����      C  , ,  ������  ����إ  �.��إ  �.����  ������      C  , ,  ������  ����إ  �|��إ  �|����  ������      C  , ,  � ����  � ��إ  ����إ  ������  � ����      C  , ,  `@���3  `@����  `�����  `����3  `@���3      C  , ,  ix���+  ix����  j"����  j"���+  ix���+      C  , ,  b����3  b�����  c8����  c8���3  b����3      C  , ,  d����3  d�����  e�����  e����3  d����3      C  , ,  g*���3  g*����  g�����  g����3  g*���3      C  , ,  ix���3  ix����  j"����  j"���3  ix���3      C  , ,  k����3  k�����  lp����  lp���3  k����3      C  , ,  n���3  n����  n�����  n����3  n���3      C  , ,  pb���3  pb����  q����  q���3  pb���3      C  , ,  k����+  k�����  lp����  lp���+  k����+      C  , ,  n���+  n����  n�����  n����+  n���+      C  , ,  pb���+  pb����  q����  q���+  pb���+      C  , ,  b���֓  b����=  c8���=  c8��֓  b���֓      C  , ,  d���֓  d����=  e����=  e���֓  d���֓      C  , ,  g*��֓  g*���=  g����=  g���֓  g*��֓      C  , ,  ix��֓  ix���=  j"���=  j"��֓  ix��֓      C  , ,  ]H��ϕ  ]H���?  ]����?  ]���ϕ  ]H��ϕ      C  , ,  ^���ϕ  ^����?  _Z���?  _Z��ϕ  ^���ϕ      C  , ,  `��ϕ  `���?  `����?  `���ϕ  `��ϕ      C  , ,  a���ϕ  a����?  b*���?  b*��ϕ  a���ϕ      C  , ,  ]�����  ]����u  ^����u  ^�����  ]�����      C  , ,  `@����  `@���u  `����u  `�����  `@����      C  , ,  b�����  b����u  c8���u  c8����  b�����      C  , ,  d�����  d����u  e����u  e�����  d�����      C  , ,  g*����  g*���u  g����u  g�����  g*����      C  , ,  ix����  ix���u  j"���u  j"����  ix����      C  , ,  k�����  k����u  lp���u  lp����  k�����      C  , ,  n����  n���u  n����u  n�����  n����      C  , ,  pb����  pb���u  q���u  q����  pb����      C  , ,  b���ϕ  b����?  c����?  c���ϕ  b���ϕ      C  , ,  dP��ϕ  dP���?  d����?  d���ϕ  dP��ϕ      C  , ,  e���ϕ  e����?  fb���?  fb��ϕ  e���ϕ      C  , ,  g ��ϕ  g ���?  g����?  g���ϕ  g ��ϕ      C  , ,  h���ϕ  h����?  i2���?  i2��ϕ  h���ϕ      C  , ,  i���ϕ  i����?  j����?  j���ϕ  i���ϕ      C  , ,  kX��ϕ  kX���?  l���?  l��ϕ  kX��ϕ      C  , ,  l���ϕ  l����?  mj���?  mj��ϕ  l���ϕ      C  , ,  n(��ϕ  n(���?  n����?  n���ϕ  n(��ϕ      C  , ,  o���ϕ  o����?  p:���?  p:��ϕ  o���ϕ      C  , ,  p���ϕ  p����?  q����?  q���ϕ  p���ϕ      C  , ,  ]����c  ]����  ^����  ^����c  ]����c      C  , ,  `@���c  `@���  `����  `����c  `@���c      C  , ,  b����c  b����  c8���  c8���c  b����c      C  , ,  d����c  d����  e����  e����c  d����c      C  , ,  g*���c  g*���  g����  g����c  g*���c      C  , ,  ix���c  ix���  j"���  j"���c  ix���c      C  , ,  k����c  k����  lp���  lp���c  k����c      C  , ,  n���c  n���  n����  n����c  n���c      C  , ,  pb���c  pb���  q���  q���c  pb���c      C  , ,  k���֓  k����=  lp���=  lp��֓  k���֓      C  , ,  n��֓  n���=  n����=  n���֓  n��֓      C  , ,  pb��֓  pb���=  q���=  q��֓  pb��֓      C  , ,  ]���֓  ]����=  ^����=  ^���֓  ]���֓      C  , ,  `@��֓  `@���=  `����=  `���֓  `@��֓      C  , ,  ]����+  ]�����  ^�����  ^����+  ]����+      C  , ,  `@���+  `@����  `�����  `����+  `@���+      C  , ,  ]�����  ]����m  ^����m  ^�����  ]�����      C  , ,  `@����  `@���m  `����m  `�����  `@����      C  , ,  b�����  b����m  c8���m  c8����  b�����      C  , ,  d�����  d����m  e����m  e�����  d�����      C  , ,  ]�����  ]���إ  ^���إ  ^�����  ]�����      C  , ,  `@����  `@��إ  `���إ  `�����  `@����      C  , ,  b�����  b���إ  c8��إ  c8����  b�����      C  , ,  d�����  d���إ  e���إ  e�����  d�����      C  , ,  g*����  g*��إ  g���إ  g�����  g*����      C  , ,  ix����  ix��إ  j"��إ  j"����  ix����      C  , ,  k�����  k���إ  lp��إ  lp����  k�����      C  , ,  n����  n��إ  n���إ  n�����  n����      C  , ,  pb����  pb��إ  q��إ  q����  pb����      C  , ,  g*����  g*���m  g����m  g�����  g*����      C  , ,  ix����  ix���m  j"���m  j"����  ix����      C  , ,  k�����  k����m  lp���m  lp����  k�����      C  , ,  n����  n���m  n����m  n�����  n����      C  , ,  pb����  pb���m  q���m  q����  pb����      C  , ,  b����+  b�����  c8����  c8���+  b����+      C  , ,  d����+  d�����  e�����  e����+  d����+      C  , ,  ]����3  ]�����  ^�����  ^����3  ]����3      C  , ,  g*���+  g*����  g�����  g����+  g*���+      C  , ,  o�����  o���·  p:��·  p:����  o�����      C  , ,  p�����  p���·  q���·  q�����  p�����      C  , ,  ]H����  ]H��·  ]���·  ]�����  ]H����      C  , ,  ^�����  ^���·  _Z��·  _Z����  ^�����      C  , ,  ]H���%  ]H����  ]�����  ]����%  ]H���%      C  , ,  ^����%  ^�����  _Z����  _Z���%  ^����%      C  , ,  `���%  `����  `�����  `����%  `���%      C  , ,  a����%  a�����  b*����  b*���%  a����%      C  , ,  b����%  b�����  c�����  c����%  b����%      C  , ,  dP���%  dP����  d�����  d����%  dP���%      C  , ,  e����%  e�����  fb����  fb���%  e����%      C  , ,  g ���%  g ����  g�����  g����%  g ���%      C  , ,  h����%  h�����  i2����  i2���%  h����%      C  , ,  i����%  i�����  j�����  j����%  i����%      C  , ,  kX���%  kX����  l����  l���%  kX���%      C  , ,  l����%  l�����  mj����  mj���%  l����%      C  , ,  n(���%  n(����  n�����  n����%  n(���%      C  , ,  o����%  o�����  p:����  p:���%  o����%      C  , ,  p����%  p�����  q�����  q����%  p����%      C  , ,  `����  `��·  `���·  `�����  `����      C  , ,  a�����  a���·  b*��·  b*����  a�����      C  , ,  ]�����  ]���Ə  ^���Ə  ^�����  ]�����      C  , ,  `@����  `@��Ə  `���Ə  `�����  `@����      C  , ,  b�����  b���Ə  c8��Ə  c8����  b�����      C  , ,  d�����  d���Ə  e���Ə  e�����  d�����      C  , ,  g*����  g*��Ə  g���Ə  g�����  g*����      C  , ,  ix����  ix��Ə  j"��Ə  j"����  ix����      C  , ,  k�����  k���Ə  lp��Ə  lp����  k�����      C  , ,  n����  n��Ə  n���Ə  n�����  n����      C  , ,  pb����  pb��Ə  q��Ə  q����  pb����      C  , ,  ]����}  ]����'  ^����'  ^����}  ]����}      C  , ,  `@���}  `@���'  `����'  `����}  `@���}      C  , ,  b����}  b����'  c8���'  c8���}  b����}      C  , ,  d����}  d����'  e����'  e����}  d����}      C  , ,  g*���}  g*���'  g����'  g����}  g*���}      C  , ,  ix���}  ix���'  j"���'  j"���}  ix���}      C  , ,  k����}  k����'  lp���'  lp���}  k����}      C  , ,  n���}  n���'  n����'  n����}  n���}      C  , ,  pb���}  pb���'  q���'  q���}  pb���}      C  , ,  ]����  ]���ÿ  ^���ÿ  ^����  ]����      C  , ,  `@���  `@��ÿ  `���ÿ  `����  `@���      C  , ,  b����  b���ÿ  c8��ÿ  c8���  b����      C  , ,  d����  d���ÿ  e���ÿ  e����  d����      C  , ,  g*���  g*��ÿ  g���ÿ  g����  g*���      C  , ,  ix���  ix��ÿ  j"��ÿ  j"���  ix���      C  , ,  k����  k���ÿ  lp��ÿ  lp���  k����      C  , ,  n���  n��ÿ  n���ÿ  n����  n���      C  , ,  pb���  pb��ÿ  q��ÿ  q���  pb���      C  , ,  ]�����  ]����W  ^����W  ^�����  ]�����      C  , ,  `@����  `@���W  `����W  `�����  `@����      C  , ,  b�����  b����W  c8���W  c8����  b�����      C  , ,  d�����  d����W  e����W  e�����  d�����      C  , ,  g*����  g*���W  g����W  g�����  g*����      C  , ,  ix����  ix���W  j"���W  j"����  ix����      C  , ,  k�����  k����W  lp���W  lp����  k�����      C  , ,  n����  n���W  n����W  n�����  n����      C  , ,  pb����  pb���W  q���W  q����  pb����      C  , ,  b�����  b���·  c���·  c�����  b�����      C  , ,  dP����  dP��·  d���·  d�����  dP����      C  , ,  e�����  e���·  fb��·  fb����  e�����      C  , ,  g ����  g ��·  g���·  g�����  g ����      C  , ,  h�����  h���·  i2��·  i2����  h�����      C  , ,  i�����  i���·  j���·  j�����  i�����      C  , ,  kX����  kX��·  l��·  l����  kX����      C  , ,  l�����  l���·  mj��·  mj����  l�����      C  , ,  n(����  n(��·  n���·  n�����  n(����      C  , ,  � ����  � ���W  �����W  ������  � ����      C  , ,  �n����  �n���W  ����W  �����  �n����      C  , ,  ������  �����W  �f���W  �f����  ������      C  , ,  x ����  x ��·  x���·  x�����  x ����      C  , ,  yh����  yh��·  z��·  z����  yh����      C  , ,  z�����  z���·  {z��·  {z����  z�����      C  , ,  |8����  |8��·  |���·  |�����  |8����      C  , ,  }�����  }���·  ~J��·  ~J����  }�����      C  , ,  ����  ��·  ���·  �����  ����      C  , ,  �p����  �p��·  ���·  �����  �p����      C  , ,  r�����  r���Ə  sZ��Ə  sZ����  r�����      C  , ,  t�����  t���Ə  u���Ə  u�����  t�����      C  , ,  wL����  wL��Ə  w���Ə  w�����  wL����      C  , ,  y�����  y���Ə  zD��Ə  zD����  y�����      C  , ,  {�����  {���Ə  |���Ə  |�����  {�����      C  , ,  ~6����  ~6��Ə  ~���Ə  ~�����  ~6����      C  , ,  ������  ����Ə  �.��Ə  �.����  ������      C  , ,  ������  ����Ə  �|��Ə  �|����  ������      C  , ,  � ����  � ��Ə  ����Ə  ������  � ����      C  , ,  �n����  �n��Ə  ���Ə  �����  �n����      C  , ,  ������  ����Ə  �f��Ə  �f����  ������      C  , ,  ������  ����·  ����·  ������  ������      C  , ,  �@����  �@��·  ����·  ������  �@����      C  , ,  ������  ����·  �R��·  �R����  ������      C  , ,  �����  ���·  ����·  ������  �����      C  , ,  �x����  �x��·  �"��·  �"����  �x����      C  , ,  ������  ����·  ����·  ������  ������      C  , ,  �H����  �H��·  ����·  ������  �H����      C  , ,  s����%  s�����  tr����  tr���%  s����%      C  , ,  u0���%  u0����  u�����  u����%  u0���%      C  , ,  r����}  r����'  sZ���'  sZ���}  r����}      C  , ,  t����}  t����'  u����'  u����}  t����}      C  , ,  wL���}  wL���'  w����'  w����}  wL���}      C  , ,  y����}  y����'  zD���'  zD���}  y����}      C  , ,  {����}  {����'  |����'  |����}  {����}      C  , ,  ~6���}  ~6���'  ~����'  ~����}  ~6���}      C  , ,  �����}  �����'  �.���'  �.���}  �����}      C  , ,  �����}  �����'  �|���'  �|���}  �����}      C  , ,  � ���}  � ���'  �����'  �����}  � ���}      C  , ,  �n���}  �n���'  ����'  ����}  �n���}      C  , ,  �����}  �����'  �f���'  �f���}  �����}      C  , ,  v����%  v�����  wB����  wB���%  v����%      C  , ,  x ���%  x ����  x�����  x����%  x ���%      C  , ,  yh���%  yh����  z����  z���%  yh���%      C  , ,  z����%  z�����  {z����  {z���%  z����%      C  , ,  |8���%  |8����  |�����  |����%  |8���%      C  , ,  }����%  }�����  ~J����  ~J���%  }����%      C  , ,  ���%  ����  �����  ����%  ���%      C  , ,  �p���%  �p����  �����  ����%  �p���%      C  , ,  �����%  ������  ������  �����%  �����%      C  , ,  r����  r���ÿ  sZ��ÿ  sZ���  r����      C  , ,  t����  t���ÿ  u���ÿ  u����  t����      C  , ,  wL���  wL��ÿ  w���ÿ  w����  wL���      C  , ,  y����  y���ÿ  zD��ÿ  zD���  y����      C  , ,  {����  {���ÿ  |���ÿ  |����  {����      C  , ,  ~6���  ~6��ÿ  ~���ÿ  ~����  ~6���      C  , ,  �����  ����ÿ  �.��ÿ  �.���  �����      C  , ,  �����  ����ÿ  �|��ÿ  �|���  �����      C  , ,  � ���  � ��ÿ  ����ÿ  �����  � ���      C  , ,  �n���  �n��ÿ  ���ÿ  ����  �n���      C  , ,  �����  ����ÿ  �f��ÿ  �f���  �����      C  , ,  �@���%  �@����  ������  �����%  �@���%      C  , ,  �����%  ������  �R����  �R���%  �����%      C  , ,  ����%  �����  ������  �����%  ����%      C  , ,  �x���%  �x����  �"����  �"���%  �x���%      C  , ,  �����%  ������  ������  �����%  �����%      C  , ,  �H���%  �H����  ������  �����%  �H���%      C  , ,  s�����  s���·  tr��·  tr����  s�����      C  , ,  u0����  u0��·  u���·  u�����  u0����      C  , ,  v�����  v���·  wB��·  wB����  v�����      C  , ,  r�����  r����W  sZ���W  sZ����  r�����      C  , ,  t�����  t����W  u����W  u�����  t�����      C  , ,  wL����  wL���W  w����W  w�����  wL����      C  , ,  y�����  y����W  zD���W  zD����  y�����      C  , ,  {�����  {����W  |����W  |�����  {�����      C  , ,  ~6����  ~6���W  ~����W  ~�����  ~6����      C  , ,  ������  �����W  �.���W  �.����  ������      C  , ,  ������  �����W  �|���W  �|����  ������      C  , ,  ����c  ����  �����  �����c  ����c      C  , ,  ����+  �����  ������  �����+  ����+      C  , ,  �����  ����u  �����u  ������  �����      C  , ,  �����  ���Ə  ����Ə  ������  �����      C  , ,  �����  ����m  �����m  ������  �����      C  , ,  ����}  ����'  �����'  �����}  ����}      C  , ,  �����  ���إ  ����إ  ������  �����      C  , ,  ����  ���ÿ  ����ÿ  �����  ����      C  , ,  �����  ����W  �����W  ������  �����      C  , ,  ����3  �����  ������  �����3  ����3      C  , ,  ���֓  ����=  �����=  ����֓  ���֓      C  , ,  � ���+  � ����  ������  �����+  � ���+      C  , ,  �N���+  �N����  ������  �����+  �N���+      C  , ,  �����+  ������  �F����  �F���+  �����+      C  , ,  �����+  ������  ������  �����+  �����+      C  , ,  �8���+  �8����  ������  �����+  �8���+      C  , ,  �����+  ������  �0����  �0���+  �����+      C  , ,  �����+  ������  �~����  �~���+  �����+      C  , ,  �"���+  �"����  ������  �����+  �"���+      C  , ,  �����c  �����  �0���  �0���c  �����c      C  , ,  �����c  �����  �~���  �~���c  �����c      C  , ,  �"���c  �"���  �����  �����c  �"���c      C  , ,  �����3  ������  �~����  �~���3  �����3      C  , ,  �����c  �����  �\���  �\���c  �����c      C  , ,  �d����  �d���u  ����u  �����  �d����      C  , ,  � ���c  � ���  �����  �����c  � ���c      C  , ,  ������  �����u  �\���u  �\����  ������      C  , ,  � ����  � ���u  �����u  ������  � ����      C  , ,  �N����  �N���u  �����u  ������  �N����      C  , ,  ������  �����u  �F���u  �F����  ������      C  , ,  �N���c  �N���  �����  �����c  �N���c      C  , ,  �d����  �d���m  ����m  �����  �d����      C  , ,  ������  �����m  �\���m  �\����  ������      C  , ,  � ����  � ���m  �����m  ������  � ����      C  , ,  �N����  �N���m  �����m  ������  �N����      C  , ,  ������  �����m  �F���m  �F����  ������      C  , ,  �����c  �����  �F���  �F���c  �����c      C  , ,  ������  �����m  �����m  ������  ������      C  , ,  �8����  �8���m  �����m  ������  �8����      C  , ,  ������  �����m  �0���m  �0����  ������      C  , ,  ������  �����m  �~���m  �~����  ������      C  , ,  �"����  �"���m  �����m  ������  �"����      C  , ,  ������  �����u  �����u  ������  ������      C  , ,  �8����  �8���u  �����u  ������  �8����      C  , ,  ������  �����u  �0���u  �0����  ������      C  , ,  �����c  �����  �����  �����c  �����c      C  , ,  �d����  �d��إ  ���إ  �����  �d����      C  , ,  �8���c  �8���  �����  �����c  �8���c      C  , ,  ������  ����إ  �\��إ  �\����  ������      C  , ,  � ����  � ��إ  ����إ  ������  � ����      C  , ,  �N����  �N��إ  ����إ  ������  �N����      C  , ,  ������  ����إ  �F��إ  �F����  ������      C  , ,  ������  ����إ  ����إ  ������  ������      C  , ,  �8����  �8��إ  ����إ  ������  �8����      C  , ,  ������  ����إ  �0��إ  �0����  ������      C  , ,  ������  ����إ  �~��إ  �~����  ������      C  , ,  �"����  �"��إ  ����إ  ������  �"����      C  , ,  ������  �����u  �~���u  �~����  ������      C  , ,  �"����  �"���u  �����u  ������  �"����      C  , ,  �"���3  �"����  ������  �����3  �"���3      C  , ,  �d���c  �d���  ����  ����c  �d���c      C  , ,  ����ϕ  �����?  �B���?  �B��ϕ  ����ϕ      C  , ,  � ��ϕ  � ���?  �����?  ����ϕ  � ��ϕ      C  , ,  �h��ϕ  �h���?  ����?  ���ϕ  �h��ϕ      C  , ,  ����ϕ  �����?  �z���?  �z��ϕ  ����ϕ      C  , ,  �8��ϕ  �8���?  �����?  ����ϕ  �8��ϕ      C  , ,  ����ϕ  �����?  �J���?  �J��ϕ  ����ϕ      C  , ,  ���ϕ  ����?  �����?  ����ϕ  ���ϕ      C  , ,  �p��ϕ  �p���?  ����?  ���ϕ  �p��ϕ      C  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      C  , ,  �@��ϕ  �@���?  �����?  ����ϕ  �@��ϕ      C  , ,  ����ϕ  �����?  �R���?  �R��ϕ  ����ϕ      C  , ,  ���ϕ  ����?  �����?  ����ϕ  ���ϕ      C  , ,  �x��ϕ  �x���?  �"���?  �"��ϕ  �x��ϕ      C  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      C  , ,  �H��ϕ  �H���?  �����?  ����ϕ  �H��ϕ      C  , ,  ����ϕ  �����?  �Z���?  �Z��ϕ  ����ϕ      C  , ,  ���ϕ  ����?  �����?  ����ϕ  ���ϕ      C  , ,  �d���+  �d����  �����  ����+  �d���+      C  , ,  �d���3  �d����  �����  ����3  �d���3      C  , ,  �����3  ������  �\����  �\���3  �����3      C  , ,  � ���3  � ����  ������  �����3  � ���3      C  , ,  �N���3  �N����  ������  �����3  �N���3      C  , ,  �����3  ������  �F����  �F���3  �����3      C  , ,  �����3  ������  ������  �����3  �����3      C  , ,  �����+  ������  �\����  �\���+  �����+      C  , ,  �d��֓  �d���=  ����=  ���֓  �d��֓      C  , ,  ����֓  �����=  �\���=  �\��֓  ����֓      C  , ,  � ��֓  � ���=  �����=  ����֓  � ��֓      C  , ,  �N��֓  �N���=  �����=  ����֓  �N��֓      C  , ,  ����֓  �����=  �F���=  �F��֓  ����֓      C  , ,  ����֓  �����=  �����=  ����֓  ����֓      C  , ,  �8��֓  �8���=  �����=  ����֓  �8��֓      C  , ,  ����֓  �����=  �0���=  �0��֓  ����֓      C  , ,  ����֓  �����=  �~���=  �~��֓  ����֓      C  , ,  �"��֓  �"���=  �����=  ����֓  �"��֓      C  , ,  �8���3  �8����  ������  �����3  �8���3      C  , ,  �����3  ������  �0����  �0���3  �����3      C  , ,  ������  �����u  �:���u  �:����  ������      C  , ,  ������  �����u  �����u  ������  ������      C  , ,  �,����  �,���u  �����u  ������  �,����      C  , ,  �z����  �z���u  �$���u  �$����  �z����      C  , ,  ������  �����u  �r���u  �r����  ������      C  , ,  �����+  ������  �:����  �:���+  �����+      C  , ,  �����+  ������  ������  �����+  �����+      C  , ,  �,���+  �,����  ������  �����+  �,���+      C  , ,  �z���+  �z����  �$����  �$���+  �z���+      C  , ,  �����+  ������  �r����  �r���+  �����+      C  , ,  �z���c  �z���  �$���  �$���c  �z���c      C  , ,  �����c  �����  �r���  �r���c  �����c      C  , ,  �
���3  �
����  ������  �����3  �
���3      C  , ,  �X���3  �X����  �����  ����3  �X���3      C  , ,  �����3  ������  �P����  �P���3  �����3      C  , ,  �����3  ������  ������  �����3  �����3      C  , ,  �B���3  �B����  ������  �����3  �B���3      C  , ,  �����3  ������  �:����  �:���3  �����3      C  , ,  ����ϕ  �����?  �Z���?  �Z��ϕ  ����ϕ      C  , ,  ���ϕ  ����?  �����?  ����ϕ  ���ϕ      C  , ,  �
����  �
���m  �����m  ������  �
����      C  , ,  ����ϕ  �����?  �*���?  �*��ϕ  ����ϕ      C  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      C  , ,  �P��ϕ  �P���?  �����?  ����ϕ  �P��ϕ      C  , ,  ����ϕ  �����?  �b���?  �b��ϕ  ����ϕ      C  , ,  � ��ϕ  � ���?  �����?  ����ϕ  � ��ϕ      C  , ,  ����ϕ  �����?  �2���?  �2��ϕ  ����ϕ      C  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      C  , ,  �X��ϕ  �X���?  ����?  ���ϕ  �X��ϕ      C  , ,  ����ϕ  �����?  �j���?  �j��ϕ  ����ϕ      C  , ,  �(��ϕ  �(���?  �����?  ����ϕ  �(��ϕ      C  , ,  ����ϕ  �����?  �:���?  �:��ϕ  ����ϕ      C  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      C  , ,  �`��ϕ  �`���?  �
���?  �
��ϕ  �`��ϕ      C  , ,  ����ϕ  �����?  �r���?  �r��ϕ  ����ϕ      C  , ,  �0��ϕ  �0���?  �����?  ����ϕ  �0��ϕ      C  , ,  �X����  �X���m  ����m  �����  �X����      C  , ,  ������  �����m  �P���m  �P����  ������      C  , ,  ������  �����m  �����m  ������  ������      C  , ,  �B����  �B���m  �����m  ������  �B����      C  , ,  ������  �����m  �:���m  �:����  ������      C  , ,  ������  �����m  �����m  ������  ������      C  , ,  �,����  �,���m  �����m  ������  �,����      C  , ,  �z����  �z���m  �$���m  �$����  �z����      C  , ,  ������  �����m  �r���m  �r����  ������      C  , ,  �
���c  �
���  �����  �����c  �
���c      C  , ,  �X���c  �X���  ����  ����c  �X���c      C  , ,  �����c  �����  �P���  �P���c  �����c      C  , ,  �����c  �����  �����  �����c  �����c      C  , ,  �B���c  �B���  �����  �����c  �B���c      C  , ,  �����c  �����  �:���  �:���c  �����c      C  , ,  �����c  �����  �����  �����c  �����c      C  , ,  �,���c  �,���  �����  �����c  �,���c      C  , ,  �����3  ������  ������  �����3  �����3      C  , ,  �,���3  �,����  ������  �����3  �,���3      C  , ,  �z���3  �z����  �$����  �$���3  �z���3      C  , ,  �����3  ������  �r����  �r���3  �����3      C  , ,  �
���+  �
����  ������  �����+  �
���+      C  , ,  �X���+  �X����  �����  ����+  �X���+      C  , ,  �����+  ������  �P����  �P���+  �����+      C  , ,  �����+  ������  ������  �����+  �����+      C  , ,  �B���+  �B����  ������  �����+  �B���+      C  , ,  �
����  �
���u  �����u  ������  �
����      C  , ,  �X����  �X���u  ����u  �����  �X����      C  , ,  �
��֓  �
���=  �����=  ����֓  �
��֓      C  , ,  �X��֓  �X���=  ����=  ���֓  �X��֓      C  , ,  ����֓  �����=  �P���=  �P��֓  ����֓      C  , ,  ����֓  �����=  �����=  ����֓  ����֓      C  , ,  �B��֓  �B���=  �����=  ����֓  �B��֓      C  , ,  ����֓  �����=  �:���=  �:��֓  ����֓      C  , ,  ����֓  �����=  �����=  ����֓  ����֓      C  , ,  �,��֓  �,���=  �����=  ����֓  �,��֓      C  , ,  �z��֓  �z���=  �$���=  �$��֓  �z��֓      C  , ,  ����֓  �����=  �r���=  �r��֓  ����֓      C  , ,  �
����  �
��إ  ����إ  ������  �
����      C  , ,  �X����  �X��إ  ���إ  �����  �X����      C  , ,  ������  ����إ  �P��إ  �P����  ������      C  , ,  ������  ����إ  ����إ  ������  ������      C  , ,  �B����  �B��إ  ����إ  ������  �B����      C  , ,  ������  ����إ  �:��إ  �:����  ������      C  , ,  ������  ����إ  ����إ  ������  ������      C  , ,  �,����  �,��إ  ����إ  ������  �,����      C  , ,  �z����  �z��إ  �$��إ  �$����  �z����      C  , ,  ������  ����إ  �r��إ  �r����  ������      C  , ,  ������  �����u  �P���u  �P����  ������      C  , ,  ������  �����u  �����u  ������  ������      C  , ,  �B����  �B���u  �����u  ������  �B����      C  , ,  �����}  �����'  �r���'  �r���}  �����}      C  , ,  �X���%  �X����  �����  ����%  �X���%      C  , ,  �����%  ������  �j����  �j���%  �����%      C  , ,  �(���%  �(����  ������  �����%  �(���%      C  , ,  �����%  ������  �:����  �:���%  �����%      C  , ,  �
����  �
��Ə  ����Ə  ������  �
����      C  , ,  �X����  �X��Ə  ���Ə  �����  �X����      C  , ,  ������  ����Ə  �P��Ə  �P����  ������      C  , ,  ������  ����Ə  ����Ə  ������  ������      C  , ,  �B����  �B��Ə  ����Ə  ������  �B����      C  , ,  ������  ����Ə  �:��Ə  �:����  ������      C  , ,  ������  ����Ə  ����Ə  ������  ������      C  , ,  �,����  �,��Ə  ����Ə  ������  �,����      C  , ,  �z����  �z��Ə  �$��Ə  �$����  �z����      C  , ,  ������  ����Ə  �r��Ə  �r����  ������      C  , ,  �����%  ������  ������  �����%  �����%      C  , ,  �`���%  �`����  �
����  �
���%  �`���%      C  , ,  �����%  ������  �r����  �r���%  �����%      C  , ,  �0���%  �0����  ������  �����%  �0���%      C  , ,  �(����  �(��·  ����·  ������  �(����      C  , ,  ������  ����·  �:��·  �:����  ������      C  , ,  ������  ����·  ����·  ������  ������      C  , ,  �
���  �
��ÿ  ����ÿ  �����  �
���      C  , ,  �X���  �X��ÿ  ���ÿ  ����  �X���      C  , ,  �����  ����ÿ  �P��ÿ  �P���  �����      C  , ,  �����  ����ÿ  ����ÿ  �����  �����      C  , ,  �B���  �B��ÿ  ����ÿ  �����  �B���      C  , ,  �����  ����ÿ  �:��ÿ  �:���  �����      C  , ,  �����  ����ÿ  ����ÿ  �����  �����      C  , ,  �,���  �,��ÿ  ����ÿ  �����  �,���      C  , ,  �z���  �z��ÿ  �$��ÿ  �$���  �z���      C  , ,  �����  ����ÿ  �r��ÿ  �r���  �����      C  , ,  �`����  �`��·  �
��·  �
����  �`����      C  , ,  ������  ����·  �r��·  �r����  ������      C  , ,  �0����  �0��·  ����·  ������  �0����      C  , ,  �X����  �X��·  ���·  �����  �X����      C  , ,  ������  ����·  �j��·  �j����  ������      C  , ,  �����%  ������  �Z����  �Z���%  �����%      C  , ,  ����%  �����  ������  �����%  ����%      C  , ,  �����%  ������  �*����  �*���%  �����%      C  , ,  �����%  ������  ������  �����%  �����%      C  , ,  �P���%  �P����  ������  �����%  �P���%      C  , ,  �����%  ������  �b����  �b���%  �����%      C  , ,  � ���%  � ����  ������  �����%  � ���%      C  , ,  �����%  ������  �2����  �2���%  �����%      C  , ,  �����%  ������  ������  �����%  �����%      C  , ,  �
���}  �
���'  �����'  �����}  �
���}      C  , ,  �X���}  �X���'  ����'  ����}  �X���}      C  , ,  �����}  �����'  �P���'  �P���}  �����}      C  , ,  �����}  �����'  �����'  �����}  �����}      C  , ,  �B���}  �B���'  �����'  �����}  �B���}      C  , ,  �����}  �����'  �:���'  �:���}  �����}      C  , ,  �����}  �����'  �����'  �����}  �����}      C  , ,  �
����  �
���W  �����W  ������  �
����      C  , ,  �X����  �X���W  ����W  �����  �X����      C  , ,  ������  �����W  �P���W  �P����  ������      C  , ,  ������  �����W  �����W  ������  ������      C  , ,  �B����  �B���W  �����W  ������  �B����      C  , ,  ������  �����W  �:���W  �:����  ������      C  , ,  ������  �����W  �����W  ������  ������      C  , ,  �,����  �,���W  �����W  ������  �,����      C  , ,  �z����  �z���W  �$���W  �$����  �z����      C  , ,  ������  �����W  �r���W  �r����  ������      C  , ,  �,���}  �,���'  �����'  �����}  �,���}      C  , ,  �z���}  �z���'  �$���'  �$���}  �z���}      C  , ,  ������  ����·  �Z��·  �Z����  ������      C  , ,  �����  ���·  ����·  ������  �����      C  , ,  ������  ����·  �*��·  �*����  ������      C  , ,  ������  ����·  ����·  ������  ������      C  , ,  �P����  �P��·  ����·  ������  �P����      C  , ,  ������  ����·  �b��·  �b����  ������      C  , ,  � ����  � ��·  ����·  ������  � ����      C  , ,  ������  ����·  �2��·  �2����  ������      C  , ,  ������  ����·  ����·  ������  ������      C  , ,  �8����  �8��Ə  ����Ə  ������  �8����      C  , ,  ������  ����Ə  �0��Ə  �0����  ������      C  , ,  ������  ����Ə  �~��Ə  �~����  ������      C  , ,  �"����  �"��Ə  ����Ə  ������  �"����      C  , ,  �����%  ������  �Z����  �Z���%  �����%      C  , ,  ����%  �����  ������  �����%  ����%      C  , ,  ������  ����·  �B��·  �B����  ������      C  , ,  � ����  � ��·  ����·  ������  � ����      C  , ,  �h����  �h��·  ���·  �����  �h����      C  , ,  ������  ����·  �z��·  �z����  ������      C  , ,  �8����  �8��·  ����·  ������  �8����      C  , ,  ������  ����·  �J��·  �J����  ������      C  , ,  �����  ���·  ����·  ������  �����      C  , ,  �p����  �p��·  ���·  �����  �p����      C  , ,  ������  ����·  ����·  ������  ������      C  , ,  �@����  �@��·  ����·  ������  �@����      C  , ,  ������  ����·  �R��·  �R����  ������      C  , ,  �����  ���·  ����·  ������  �����      C  , ,  �x����  �x��·  �"��·  �"����  �x����      C  , ,  ������  ����·  ����·  ������  ������      C  , ,  �H����  �H��·  ����·  ������  �H����      C  , ,  ������  ����·  �Z��·  �Z����  ������      C  , ,  �d���  �d��ÿ  ���ÿ  ����  �d���      C  , ,  �����  ����ÿ  �\��ÿ  �\���  �����      C  , ,  � ���  � ��ÿ  ����ÿ  �����  � ���      C  , ,  �N���  �N��ÿ  ����ÿ  �����  �N���      C  , ,  �����  ����ÿ  �F��ÿ  �F���  �����      C  , ,  �����  ����ÿ  ����ÿ  �����  �����      C  , ,  �8���  �8��ÿ  ����ÿ  �����  �8���      C  , ,  �����  ����ÿ  �0��ÿ  �0���  �����      C  , ,  �����  ����ÿ  �~��ÿ  �~���  �����      C  , ,  �"���  �"��ÿ  ����ÿ  �����  �"���      C  , ,  �����  ���·  ����·  ������  �����      C  , ,  �����%  ������  �B����  �B���%  �����%      C  , ,  � ���%  � ����  ������  �����%  � ���%      C  , ,  �h���%  �h����  �����  ����%  �h���%      C  , ,  �����%  ������  �z����  �z���%  �����%      C  , ,  �8���%  �8����  ������  �����%  �8���%      C  , ,  �����%  ������  �J����  �J���%  �����%      C  , ,  ����%  �����  ������  �����%  ����%      C  , ,  �p���%  �p����  �����  ����%  �p���%      C  , ,  �����%  ������  ������  �����%  �����%      C  , ,  �@���%  �@����  ������  �����%  �@���%      C  , ,  �����%  ������  �R����  �R���%  �����%      C  , ,  ����%  �����  ������  �����%  ����%      C  , ,  �d���}  �d���'  ����'  ����}  �d���}      C  , ,  �����}  �����'  �\���'  �\���}  �����}      C  , ,  � ���}  � ���'  �����'  �����}  � ���}      C  , ,  �N���}  �N���'  �����'  �����}  �N���}      C  , ,  �����}  �����'  �F���'  �F���}  �����}      C  , ,  �����}  �����'  �����'  �����}  �����}      C  , ,  �8���}  �8���'  �����'  �����}  �8���}      C  , ,  �����}  �����'  �0���'  �0���}  �����}      C  , ,  �����}  �����'  �~���'  �~���}  �����}      C  , ,  �"���}  �"���'  �����'  �����}  �"���}      C  , ,  �x���%  �x����  �"����  �"���%  �x���%      C  , ,  �����%  ������  ������  �����%  �����%      C  , ,  �H���%  �H����  ������  �����%  �H���%      C  , ,  �d����  �d��Ə  ���Ə  �����  �d����      C  , ,  ������  ����Ə  �\��Ə  �\����  ������      C  , ,  � ����  � ��Ə  ����Ə  ������  � ����      C  , ,  �N����  �N��Ə  ����Ə  ������  �N����      C  , ,  ������  ����Ə  �F��Ə  �F����  ������      C  , ,  �d����  �d���W  ����W  �����  �d����      C  , ,  ������  �����W  �\���W  �\����  ������      C  , ,  � ����  � ���W  �����W  ������  � ����      C  , ,  �N����  �N���W  �����W  ������  �N����      C  , ,  ������  �����W  �F���W  �F����  ������      C  , ,  ������  �����W  �����W  ������  ������      C  , ,  �8����  �8���W  �����W  ������  �8����      C  , ,  ������  �����W  �0���W  �0����  ������      C  , ,  ������  �����W  �~���W  �~����  ������      C  , ,  �"����  �"���W  �����W  ������  �"����      C  , ,  ������  ����Ə  ����Ə  ������  ������      C  , ,  ������  ������  Ě����  Ě����  ������      C  , ,  �X����  �X����  �����  �����  �X����      C  , ,  ������  ������  �j����  �j����  ������      C  , ,  �(����  �(����  ������  ������  �(����      C  , ,  ɐ����  ɐ����  �:����  �:����  ɐ����      C  , ,  ������  ������  ˢ����  ˢ����  ������      C  , ,  �`����  �`����  �
����  �
����  �`����      C  , ,  ������  ������  �r����  �r����  ������      C  , ,  �0����  �0����  ������  ������  �0����      C  , ,  И����  И����  �B����  �B����  И����      C  , ,  � ����  � ����  Ҫ����  Ҫ����  � ����      C  , ,  ����  ���I  �2���I  �2����  ����      C  , ,  ������  �����I  Ě���I  Ě����  ������      C  , ,  �X����  �X���I  ����I  �����  �X����      C  , ,  ������  �����I  �j���I  �j����  ������      C  , ,  �����/  ������  ������  �����/  �����/      C  , ,  �P���/  �P����  ������  �����/  �P���/      C  , ,  �p���  �p���1  ����1  ����  �p���      C  , ,  �����  �����1  �h���1  �h���  �����      C  , ,  ����  ����1  �����1  �����  ����      C  , ,  �Z���  �Z���1  ����1  ����  �Z���      C  , ,  Ũ���  Ũ���1  �R���1  �R���  Ũ���      C  , ,  �����  �����1  Ƞ���1  Ƞ���  �����      C  , ,  �D���  �D���1  �����1  �����  �D���      C  , ,  ̒���  ̒���1  �<���1  �<���  ̒���      C  , ,  �����  �����1  ϊ���1  ϊ���  �����      C  , ,  �.���  �.���1  �����1  �����  �.���      C  , ,  �����/  ������  �b����  �b���/  �����/      C  , ,  � ���/  � ����  ������  �����/  � ���/      C  , ,  ���/  ����  �2����  �2���/  ���/      C  , ,  �����/  ������  Ě����  Ě���/  �����/      C  , ,  �X���/  �X����  �����  ����/  �X���/      C  , ,  �����/  ������  �j����  �j���/  �����/      C  , ,  �(���/  �(����  ������  �����/  �(���/      C  , ,  �p����  �p���  ����  �����  �p����      C  , ,  ������  �����  �h���  �h����  ������      C  , ,  �����  ����  �����  ������  �����      C  , ,  �Z����  �Z���  ����  �����  �Z����      C  , ,  Ũ����  Ũ���  �R���  �R����  Ũ����      C  , ,  ������  �����  Ƞ���  Ƞ����  ������      C  , ,  �D����  �D���  �����  ������  �D����      C  , ,  ̒����  ̒���  �<���  �<����  ̒����      C  , ,  ������  �����  ϊ���  ϊ����  ������      C  , ,  �.����  �.���  �����  ������  �.����      C  , ,  ɐ���/  ɐ����  �:����  �:���/  ɐ���/      C  , ,  �����/  ������  ˢ����  ˢ���/  �����/      C  , ,  �`���/  �`����  �
����  �
���/  �`���/      C  , ,  �����/  ������  �r����  �r���/  �����/      C  , ,  �0���/  �0����  ������  �����/  �0���/      C  , ,  И���/  И����  �B����  �B���/  И���/      C  , ,  � ���/  � ����  Ҫ����  Ҫ���/  � ���/      C  , ,  �(����  �(���I  �����I  ������  �(����      C  , ,  ɐ����  ɐ���I  �:���I  �:����  ɐ����      C  , ,  ������  �����I  ˢ���I  ˢ����  ������      C  , ,  �`����  �`���I  �
���I  �
����  �`����      C  , ,  ������  �����I  �r���I  �r����  ������      C  , ,  �0����  �0���I  �����I  ������  �0����      C  , ,  И����  И���I  �B���I  �B����  И����      C  , ,  � ����  � ���I  Ҫ���I  Ҫ����  � ����      C  , ,  ������  �����I  �����I  ������  ������      C  , ,  �P����  �P���I  �����I  ������  �P����      C  , ,  ������  �����I  �b���I  �b����  ������      C  , ,  � ����  � ���I  �����I  ������  � ����      C  , ,  ������  ������  ������  ������  ������      C  , ,  �P����  �P����  ������  ������  �P����      C  , ,  ������  ������  �b����  �b����  ������      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  ����  ����  �2����  �2����  ����      C  , ,  Ũ��ݛ  Ũ���E  �R���E  �R��ݛ  Ũ��ݛ      C  , ,  ����ݛ  �����E  Ƞ���E  Ƞ��ݛ  ����ݛ      C  , ,  �D��ݛ  �D���E  �����E  ����ݛ  �D��ݛ      C  , ,  ̒��ݛ  ̒���E  �<���E  �<��ݛ  ̒��ݛ      C  , ,  ����ݛ  �����E  ϊ���E  ϊ��ݛ  ����ݛ      C  , ,  �.��ݛ  �.���E  �����E  ����ݛ  �.��ݛ      C  , ,  �����  ������  Ƞ����  Ƞ���  �����      C  , ,  �D���  �D����  ������  �����  �D���      C  , ,  ̒���  ̒����  �<����  �<���  ̒���      C  , ,  �����  ������  ϊ����  ϊ���  �����      C  , ,  �.���  �.����  ������  �����  �.���      C  , ,  �����O  ������  Ƞ����  Ƞ���O  �����O      C  , ,  �D���O  �D����  ������  �����O  �D���O      C  , ,  ̒���O  ̒����  �<����  �<���O  ̒���O      C  , ,  �����O  ������  ϊ����  ϊ���O  �����O      C  , ,  �.���O  �.����  ������  �����O  �.���O      C  , ,  �����  �����)  Ƞ���)  Ƞ���  �����      C  , ,  �D���  �D���)  �����)  �����  �D���      C  , ,  ̒���  ̒���)  �<���)  �<���  ̒���      C  , ,  �����  �����)  ϊ���)  ϊ���  �����      C  , ,  �.���  �.���)  �����)  �����  �.���      C  , ,  �����  ������  ϊ����  ϊ���  �����      C  , ,  �.���  �.����  ������  �����  �.���      C  , ,  �p���  �p���a  ����a  ����  �p���      C  , ,  �����  �����a  �h���a  �h���  �����      C  , ,  ����  ����a  �����a  �����  ����      C  , ,  �Z���  �Z���a  ����a  ����  �Z���      C  , ,  �p����  �p���  ����  �����  �p����      C  , ,  ������  �����  �h���  �h����  ������      C  , ,  �����  ����  �����  ������  �����      C  , ,  �Z����  �Z���  ����  �����  �Z����      C  , ,  Ũ����  Ũ���  �R���  �R����  Ũ����      C  , ,  ������  �����  Ƞ���  Ƞ����  ������      C  , ,  �D����  �D���  �����  ������  �D����      C  , ,  ̒����  ̒���  �<���  �<����  ̒����      C  , ,  ������  �����  ϊ���  ϊ����  ������      C  , ,  �.����  �.���  �����  ������  �.����      C  , ,  Ũ���  Ũ���a  �R���a  �R���  Ũ���      C  , ,  �����  �����a  Ƞ���a  Ƞ���  �����      C  , ,  �D���  �D���a  �����a  �����  �D���      C  , ,  ̒���  ̒���a  �<���a  �<���  ̒���      C  , ,  �����  �����a  ϊ���a  ϊ���  �����      C  , ,  �.���  �.���a  �����a  �����  �.���      C  , ,  �����  �����)  �h���)  �h���  �����      C  , ,  ����  ����)  �����)  �����  ����      C  , ,  �Z���  �Z���)  ����)  ����  �Z���      C  , ,  ������  �����u  �A���u  �A����  ������      C  , ,  ������  �����u  �����u  ������  ������      C  , ,  �3����  �3���u  �����u  ������  �3����      C  , ,  ā����  ā���u  �+���u  �+����  ā����      C  , ,  ������  �����u  �y���u  �y����  ������      C  , ,  �����  ����u  �����u  ������  �����      C  , ,  ������  �����  �A���  �A����  ������      C  , ,  ������  �����  �����  ������  ������      C  , ,  �3����  �3���  �����  ������  �3����      C  , ,  ā����  ā���  �+���  �+����  ā����      C  , ,  ������  �����  �y���  �y����  ������      C  , ,  �����  ����  �����  ������  �����      C  , ,  �k����  �k���  ����  �����  �k����      C  , ,  ͹����  ͹���  �c���  �c����  ͹����      C  , ,  �����  ����  б���  б����  �����      C  , ,  �k����  �k���u  ����u  �����  �k����      C  , ,  ͹����  ͹���u  �c���u  �c����  ͹����      C  , ,  �����  ����u  б���u  б����  �����      C  , ,  Ũ���  Ũ���)  �R���)  �R���  Ũ���      C  , ,  �p���O  �p����  �����  ����O  �p���O      C  , ,  �����O  ������  �h����  �h���O  �����O      C  , ,  ����O  �����  ������  �����O  ����O      C  , ,  �Z���O  �Z����  �����  ����O  �Z���O      C  , ,  Ũ���O  Ũ����  �R����  �R���O  Ũ���O      C  , ,  �p���  �p����  �����  ����  �p���      C  , ,  �����  ������  �h����  �h���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �Z���  �Z����  �����  ����  �Z���      C  , ,  Ũ���  Ũ����  �R����  �R���  Ũ���      C  , ,  �p��ݛ  �p���E  ����E  ���ݛ  �p��ݛ      C  , ,  ����ݛ  �����E  �h���E  �h��ݛ  ����ݛ      C  , ,  ���ݛ  ����E  �����E  ����ݛ  ���ݛ      C  , ,  �Z��ݛ  �Z���E  ����E  ���ݛ  �Z��ݛ      C  , ,  �p���  �p����  �����  ����  �p���      C  , ,  �����  ������  �h����  �h���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �Z���  �Z����  �����  ����  �Z���      C  , ,  Ũ���  Ũ����  �R����  �R���  Ũ���      C  , ,  �����  ������  Ƞ����  Ƞ���  �����      C  , ,  �D���  �D����  ������  �����  �D���      C  , ,  ̒���  ̒����  �<����  �<���  ̒���      C  , ,  �p���  �p���)  ����)  ����  �p���      C  , ,  �`��ϕ  �`���?  �
���?  �
��ϕ  �`��ϕ      C  , ,  ����ϕ  �����?  �r���?  �r��ϕ  ����ϕ      C  , ,  �0��ϕ  �0���?  �����?  ����ϕ  �0��ϕ      C  , ,  И��ϕ  И���?  �B���?  �B��ϕ  И��ϕ      C  , ,  � ��ϕ  � ���?  Ҫ���?  Ҫ��ϕ  � ��ϕ      C  , ,  ������  ����إ  Ƞ��إ  Ƞ����  ������      C  , ,  �D����  �D��إ  ����إ  ������  �D����      C  , ,  ̒����  ̒��إ  �<��إ  �<����  ̒����      C  , ,  ������  ����إ  ϊ��إ  ϊ����  ������      C  , ,  �.����  �.��إ  ����إ  ������  �.����      C  , ,  ̒���c  ̒���  �<���  �<���c  ̒���c      C  , ,  �����c  �����  ϊ���  ϊ���c  �����c      C  , ,  �.���c  �.���  �����  �����c  �.���c      C  , ,  �p����  �p���m  ����m  �����  �p����      C  , ,  ������  �����m  �h���m  �h����  ������      C  , ,  �����  ����m  �����m  ������  �����      C  , ,  �Z����  �Z���m  ����m  �����  �Z����      C  , ,  Ũ����  Ũ���m  �R���m  �R����  Ũ����      C  , ,  ������  �����m  Ƞ���m  Ƞ����  ������      C  , ,  �D����  �D���m  �����m  ������  �D����      C  , ,  ̒����  ̒���m  �<���m  �<����  ̒����      C  , ,  ������  �����m  ϊ���m  ϊ����  ������      C  , ,  �.����  �.���m  �����m  ������  �.����      C  , ,  �.����  �.���u  �����u  ������  �.����      C  , ,  ������  �����u  ϊ���u  ϊ����  ������      C  , ,  �p���3  �p����  �����  ����3  �p���3      C  , ,  �����3  ������  �h����  �h���3  �����3      C  , ,  ����3  �����  ������  �����3  ����3      C  , ,  �Z���3  �Z����  �����  ����3  �Z���3      C  , ,  Ũ���3  Ũ����  �R����  �R���3  Ũ���3      C  , ,  �����3  ������  Ƞ����  Ƞ���3  �����3      C  , ,  �D���3  �D����  ������  �����3  �D���3      C  , ,  ̒���3  ̒����  �<����  �<���3  ̒���3      C  , ,  �p��֓  �p���=  ����=  ���֓  �p��֓      C  , ,  ����֓  �����=  �h���=  �h��֓  ����֓      C  , ,  ���֓  ����=  �����=  ����֓  ���֓      C  , ,  �Z��֓  �Z���=  ����=  ���֓  �Z��֓      C  , ,  Ũ��֓  Ũ���=  �R���=  �R��֓  Ũ��֓      C  , ,  ����֓  �����=  Ƞ���=  Ƞ��֓  ����֓      C  , ,  �D��֓  �D���=  �����=  ����֓  �D��֓      C  , ,  ̒��֓  ̒���=  �<���=  �<��֓  ̒��֓      C  , ,  ����֓  �����=  ϊ���=  ϊ��֓  ����֓      C  , ,  �.��֓  �.���=  �����=  ����֓  �.��֓      C  , ,  �����3  ������  ϊ����  ϊ���3  �����3      C  , ,  �.���3  �.����  ������  �����3  �.���3      C  , ,  �p���c  �p���  ����  ����c  �p���c      C  , ,  �����c  �����  �h���  �h���c  �����c      C  , ,  ����c  ����  �����  �����c  ����c      C  , ,  �Z���c  �Z���  ����  ����c  �Z���c      C  , ,  Ũ���c  Ũ���  �R���  �R���c  Ũ���c      C  , ,  �����c  �����  Ƞ���  Ƞ���c  �����c      C  , ,  �D���c  �D���  �����  �����c  �D���c      C  , ,  �p����  �p��إ  ���إ  �����  �p����      C  , ,  ������  ����إ  �h��إ  �h����  ������      C  , ,  �����  ���إ  ����إ  ������  �����      C  , ,  �Z����  �Z��إ  ���إ  �����  �Z����      C  , ,  Ũ����  Ũ��إ  �R��إ  �R����  Ũ����      C  , ,  ����ϕ  �����?  �����?  ����ϕ  ����ϕ      C  , ,  �P��ϕ  �P���?  �����?  ����ϕ  �P��ϕ      C  , ,  ����ϕ  �����?  �b���?  �b��ϕ  ����ϕ      C  , ,  � ��ϕ  � ���?  �����?  ����ϕ  � ��ϕ      C  , ,  ��ϕ  ���?  �2���?  �2��ϕ  ��ϕ      C  , ,  ����ϕ  �����?  Ě���?  Ě��ϕ  ����ϕ      C  , ,  �X��ϕ  �X���?  ����?  ���ϕ  �X��ϕ      C  , ,  ����ϕ  �����?  �j���?  �j��ϕ  ����ϕ      C  , ,  �(��ϕ  �(���?  �����?  ����ϕ  �(��ϕ      C  , ,  �p���+  �p����  �����  ����+  �p���+      C  , ,  �����+  ������  �h����  �h���+  �����+      C  , ,  ����+  �����  ������  �����+  ����+      C  , ,  �Z���+  �Z����  �����  ����+  �Z���+      C  , ,  Ũ���+  Ũ����  �R����  �R���+  Ũ���+      C  , ,  �����+  ������  Ƞ����  Ƞ���+  �����+      C  , ,  �D���+  �D����  ������  �����+  �D���+      C  , ,  ̒���+  ̒����  �<����  �<���+  ̒���+      C  , ,  �����+  ������  ϊ����  ϊ���+  �����+      C  , ,  �.���+  �.����  ������  �����+  �.���+      C  , ,  ɐ��ϕ  ɐ���?  �:���?  �:��ϕ  ɐ��ϕ      C  , ,  ����ϕ  �����?  ˢ���?  ˢ��ϕ  ����ϕ      C  , ,  �p����  �p���u  ����u  �����  �p����      C  , ,  ������  �����u  �h���u  �h����  ������      C  , ,  �����  ����u  �����u  ������  �����      C  , ,  �Z����  �Z���u  ����u  �����  �Z����      C  , ,  Ũ����  Ũ���u  �R���u  �R����  Ũ����      C  , ,  ������  �����u  Ƞ���u  Ƞ����  ������      C  , ,  �D����  �D���u  �����u  ������  �D����      C  , ,  ̒����  ̒���u  �<���u  �<����  ̒����      C  , ,  �0���%  �0����  ������  �����%  �0���%      C  , ,  И���%  И����  �B����  �B���%  И���%      C  , ,  � ���%  � ����  Ҫ����  Ҫ���%  � ���%      C  , ,  �����  ����ÿ  �h��ÿ  �h���  �����      C  , ,  ����  ���ÿ  ����ÿ  �����  ����      C  , ,  �����%  ������  ������  �����%  �����%      C  , ,  �p����  �p��Ə  ���Ə  �����  �p����      C  , ,  ������  ����·  ����·  ������  ������      C  , ,  �P����  �P��·  ����·  ������  �P����      C  , ,  ������  ����·  �b��·  �b����  ������      C  , ,  � ����  � ��·  ����·  ������  � ����      C  , ,  ����  ��·  �2��·  �2����  ����      C  , ,  ������  ����·  Ě��·  Ě����  ������      C  , ,  �X����  �X��·  ���·  �����  �X����      C  , ,  ������  ����·  �j��·  �j����  ������      C  , ,  �(����  �(��·  ����·  ������  �(����      C  , ,  ɐ����  ɐ��·  �:��·  �:����  ɐ����      C  , ,  ������  ����·  ˢ��·  ˢ����  ������      C  , ,  �`����  �`��·  �
��·  �
����  �`����      C  , ,  ������  ����·  �r��·  �r����  ������      C  , ,  �0����  �0��·  ����·  ������  �0����      C  , ,  И����  И��·  �B��·  �B����  И����      C  , ,  � ����  � ��·  Ҫ��·  Ҫ����  � ����      C  , ,  ������  ����Ə  �h��Ə  �h����  ������      C  , ,  �����  ���Ə  ����Ə  ������  �����      C  , ,  �p���}  �p���'  ����'  ����}  �p���}      C  , ,  �����}  �����'  �h���'  �h���}  �����}      C  , ,  ����}  ����'  �����'  �����}  ����}      C  , ,  �Z���}  �Z���'  ����'  ����}  �Z���}      C  , ,  Ũ���}  Ũ���'  �R���'  �R���}  Ũ���}      C  , ,  �����}  �����'  Ƞ���'  Ƞ���}  �����}      C  , ,  �D���}  �D���'  �����'  �����}  �D���}      C  , ,  ̒���}  ̒���'  �<���'  �<���}  ̒���}      C  , ,  �����}  �����'  ϊ���'  ϊ���}  �����}      C  , ,  �.���}  �.���'  �����'  �����}  �.���}      C  , ,  �Z����  �Z��Ə  ���Ə  �����  �Z����      C  , ,  Ũ����  Ũ��Ə  �R��Ə  �R����  Ũ����      C  , ,  ������  ����Ə  Ƞ��Ə  Ƞ����  ������      C  , ,  �P���%  �P����  ������  �����%  �P���%      C  , ,  �Z���  �Z��ÿ  ���ÿ  ����  �Z���      C  , ,  Ũ���  Ũ��ÿ  �R��ÿ  �R���  Ũ���      C  , ,  �����  ����ÿ  Ƞ��ÿ  Ƞ���  �����      C  , ,  �D���  �D��ÿ  ����ÿ  �����  �D���      C  , ,  ̒���  ̒��ÿ  �<��ÿ  �<���  ̒���      C  , ,  �����  ����ÿ  ϊ��ÿ  ϊ���  �����      C  , ,  �.���  �.��ÿ  ����ÿ  �����  �.���      C  , ,  ɐ���%  ɐ����  �:����  �:���%  ɐ���%      C  , ,  �.����  �.��Ə  ����Ə  ������  �.����      C  , ,  �D����  �D��Ə  ����Ə  ������  �D����      C  , ,  ̒����  ̒��Ə  �<��Ə  �<����  ̒����      C  , ,  ������  ����Ə  ϊ��Ə  ϊ����  ������      C  , ,  ���%  ����  �2����  �2���%  ���%      C  , ,  �����%  ������  Ě����  Ě���%  �����%      C  , ,  �X���%  �X����  �����  ����%  �X���%      C  , ,  �����%  ������  �j����  �j���%  �����%      C  , ,  �(���%  �(����  ������  �����%  �(���%      C  , ,  �p���  �p��ÿ  ���ÿ  ����  �p���      C  , ,  �����%  ������  ˢ����  ˢ���%  �����%      C  , ,  �`���%  �`����  �
����  �
���%  �`���%      C  , ,  �p����  �p���W  ����W  �����  �p����      C  , ,  ������  �����W  �h���W  �h����  ������      C  , ,  �����  ����W  �����W  ������  �����      C  , ,  �Z����  �Z���W  ����W  �����  �Z����      C  , ,  Ũ����  Ũ���W  �R���W  �R����  Ũ����      C  , ,  ������  �����W  Ƞ���W  Ƞ����  ������      C  , ,  �D����  �D���W  �����W  ������  �D����      C  , ,  ̒����  ̒���W  �<���W  �<����  ̒����      C  , ,  ������  �����W  ϊ���W  ϊ����  ������      C  , ,  �.����  �.���W  �����W  ������  �.����      C  , ,  �����%  ������  �b����  �b���%  �����%      C  , ,  � ���%  � ����  ������  �����%  � ���%      C  , ,  �����%  ������  �r����  �r���%  �����%      C  , ,  �X����  �X���5  ����5  �����  �X����      C  , ,  �X����  �X���}  ����}  �����  �X����      C  , ,  �X���  �X����  �����  ����  �X���      C  , ,  ]����  ]����)  ^����)  ^����  ]����      C  , ,  `@���  `@���)  `����)  `����  `@���      C  , ,  b����  b����)  c8���)  c8���  b����      C  , ,  d����  d����)  e����)  e����  d����      C  , ,  g*���  g*���)  g����)  g����  g*���      C  , ,  ix���  ix���)  j"���)  j"���  ix���      C  , ,  k����  k����)  lp���)  lp���  k����      C  , ,  n���  n���)  n����)  n����  n���      C  , ,  pb���  pb���)  q���)  q���  pb���      C  , ,  r����  r����)  sZ���)  sZ���  r����      C  , ,  t����  t����)  u����)  u����  t����      C  , ,  wL���  wL���)  w����)  w����  wL���      C  , ,  y����  y����)  zD���)  zD���  y����      C  , ,  {����  {����)  |����)  |����  {����      C  , ,  ~6���  ~6���)  ~����)  ~����  ~6���      C  , ,  �����  �����)  �.���)  �.���  �����      C  , ,  �����  �����)  �|���)  �|���  �����      C  , ,  � ���  � ���)  �����)  �����  � ���      C  , ,  �n���  �n���)  ����)  ����  �n���      C  , ,  �����  �����)  �f���)  �f���  �����      C  , ,  �
���  �
���)  �����)  �����  �
���      C  , ,  �X���  �X���)  ����)  ����  �X���      C  , ,  �����  �����)  �P���)  �P���  �����      C  , ,  �����  �����)  �����)  �����  �����      C  , ,  �B���  �B���)  �����)  �����  �B���      C  , ,  �����  �����)  �:���)  �:���  �����      C  , ,  �����  �����)  �����)  �����  �����      C  , ,  �,���  �,���)  �����)  �����  �,���      C  , ,  �z���  �z���)  �$���)  �$���  �z���      C  , ,  �����  �����)  �r���)  �r���  �����      C  , ,  ����  ����)  �����)  �����  ����      C  , ,  �d���  �d���)  ����)  ����  �d���      C  , ,  �����  �����)  �\���)  �\���  �����      C  , ,  � ���  � ���)  �����)  �����  � ���      C  , ,  �N���  �N���)  �����)  �����  �N���      C  , ,  �����  �����)  �F���)  �F���  �����      C  , ,  �����  �����)  �����)  �����  �����      C  , ,  �8���  �8���)  �����)  �����  �8���      C  , ,  �����  �����)  �0���)  �0���  �����      C  , ,  �����  �����)  �~���)  �~���  �����      C  , ,  �"���  �"���)  �����)  �����  �"���      C  , ,  �p���  �p���)  ����)  ����  �p���      C  , ,  �����  �����)  �h���)  �h���  �����      C  , ,  ����  ����)  �����)  �����  ����      C  , ,  �Z���  �Z���)  ����)  ����  �Z���      C  , ,  Ũ���  Ũ���)  �R���)  �R���  Ũ���      C  , ,  �����  �����)  Ƞ���)  Ƞ���  �����      C  , ,  �D���  �D���)  �����)  �����  �D���      C  , ,  ̒���  ̒���)  �<���)  �<���  ̒���      C  , ,  �����  �����)  ϊ���)  ϊ���  �����      C  , ,  �.���  �.���)  �����)  �����  �.���      C  , ,  �D����  �D���;  �����;  ������  �D����      C  , ,  ̒����  ̒���;  �<���;  �<����  ̒����      C  , ,  ������  �����;  ϊ���;  ϊ����  ������      C  , ,  �.����  �.���;  �����;  ������  �.����      C  , ,  �p���)  �p����  �����  ����)  �p���)      C  , ,  �����)  ������  �h����  �h���)  �����)      C  , ,  ����)  �����  ������  �����)  ����)      C  , ,  �Z���)  �Z����  �����  ����)  �Z���)      C  , ,  Ũ���)  Ũ����  �R����  �R���)  Ũ���)      C  , ,  �����)  ������  Ƞ����  Ƞ���)  �����)      C  , ,  �D���)  �D����  ������  �����)  �D���)      C  , ,  ̒���)  ̒����  �<����  �<���)  ̒���)      C  , ,  �����)  ������  ϊ����  ϊ���)  �����)      C  , ,  �.���)  �.����  ������  �����)  �.���)      C  , ,  �p����  �p���k  ����k  �����  �p����      C  , ,  ������  �����k  �h���k  �h����  ������      C  , ,  �����  ����k  �����k  ������  �����      C  , ,  �Z����  �Z���k  ����k  �����  �Z����      C  , ,  Ũ����  Ũ���k  �R���k  �R����  Ũ����      C  , ,  ������  �����k  Ƞ���k  Ƞ����  ������      C  , ,  �D����  �D���k  �����k  ������  �D����      C  , ,  ̒����  ̒���k  �<���k  �<����  ̒����      C  , ,  ������  �����k  ϊ���k  ϊ����  ������      C  , ,  �.����  �.���k  �����k  ������  �.����      C  , ,  �p����  �p����  �����  �����  �p����      C  , ,  ������  ������  �h����  �h����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �Z����  �Z����  �����  �����  �Z����      C  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      C  , ,  ������  ������  Ƞ����  Ƞ����  ������      C  , ,  �D����  �D����  ������  ������  �D����      C  , ,  ̒����  ̒����  �<����  �<����  ̒����      C  , ,  ������  ������  ϊ����  ϊ����  ������      C  , ,  �.����  �.����  ������  ������  �.����      C  , ,  �p���u  �p���  ����  ����u  �p���u      C  , ,  �����u  �����  �h���  �h���u  �����u      C  , ,  ����u  ����  �����  �����u  ����u      C  , ,  �Z���u  �Z���  ����  ����u  �Z���u      C  , ,  Ũ���u  Ũ���  �R���  �R���u  Ũ���u      C  , ,  �����u  �����  Ƞ���  Ƞ���u  �����u      C  , ,  �D���u  �D���  �����  �����u  �D���u      C  , ,  ̒���u  ̒���  �<���  �<���u  ̒���u      C  , ,  �����u  �����  ϊ���  ϊ���u  �����u      C  , ,  �.���u  �.���  �����  �����u  �.���u      C  , ,  �p���  �p����  �����  ����  �p���      C  , ,  �����  ������  �h����  �h���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �Z���  �Z����  �����  ����  �Z���      C  , ,  Ũ���  Ũ����  �R����  �R���  Ũ���      C  , ,  �����  ������  Ƞ����  Ƞ���  �����      C  , ,  �D���  �D����  ������  �����  �D���      C  , ,  ̒���  ̒����  �<����  �<���  ̒���      C  , ,  �����  ������  ϊ����  ϊ���  �����      C  , ,  �.���  �.����  ������  �����  �.���      C  , ,  ������  ������  �A����  �A����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �3����  �3����  ������  ������  �3����      C  , ,  ā����  ā����  �+����  �+����  ā����      C  , ,  ������  ������  �y����  �y����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �k����  �k����  �����  �����  �k����      C  , ,  ͹����  ͹����  �c����  �c����  ͹����      C  , ,  �����  �����  б����  б����  �����      C  , ,  ������  �����k  �A���k  �A����  ������      C  , ,  ������  �����k  �����k  ������  ������      C  , ,  �3����  �3���k  �����k  ������  �3����      C  , ,  ā����  ā���k  �+���k  �+����  ā����      C  , ,  ������  �����k  �y���k  �y����  ������      C  , ,  �����  ����k  �����k  ������  �����      C  , ,  �k����  �k���k  ����k  �����  �k����      C  , ,  ͹����  ͹���k  �c���k  �c����  ͹����      C  , ,  �����  ����k  б���k  б����  �����      C  , ,  �p����  �p���;  ����;  �����  �p����      C  , ,  ������  �����;  �h���;  �h����  ������      C  , ,  �����  ����;  �����;  ������  �����      C  , ,  �Z����  �Z���;  ����;  �����  �Z����      C  , ,  Ũ����  Ũ���;  �R���;  �R����  Ũ����      C  , ,  ������  �����;  Ƞ���;  Ƞ����  ������      C  , ,  ������  �����5  �����5  ������  ������      C  , ,  �`����  �`���5  �
���5  �
����  �`����      C  , ,  ������  �����5  �r���5  �r����  ������      C  , ,  �0����  �0���5  �����5  ������  �0����      C  , ,  Ƙ����  Ƙ���5  �B���5  �B����  Ƙ����      C  , ,  � ����  � ���5  Ȫ���5  Ȫ����  � ����      C  , ,  �h����  �h���5  ����5  �����  �h����      C  , ,  ������  �����5  �z���5  �z����  ������      C  , ,  �8����  �8���5  �����5  ������  �8����      C  , ,  ͠����  ͠���5  �J���5  �J����  ͠����      C  , ,  �����  ����5  ϲ���5  ϲ����  �����      C  , ,  �p����  �p���5  ����5  �����  �p����      C  , ,  ������  �����5  ҂���5  ҂����  ������      C  , ,  �����Y  �����  �h���  �h���Y  �����Y      C  , ,  ������  �����}  �j���}  �j����  ������      C  , ,  �(����  �(���}  �����}  ������  �(����      C  , ,  ������  �����}  �:���}  �:����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �`����  �`���}  �
���}  �
����  �`����      C  , ,  ������  �����}  �r���}  �r����  ������      C  , ,  �0����  �0���}  �����}  ������  �0����      C  , ,  Ƙ����  Ƙ���}  �B���}  �B����  Ƙ����      C  , ,  � ����  � ���}  Ȫ���}  Ȫ����  � ����      C  , ,  �h����  �h���}  ����}  �����  �h����      C  , ,  ������  �����}  �z���}  �z����  ������      C  , ,  �8����  �8���}  �����}  ������  �8����      C  , ,  ͠����  ͠���}  �J���}  �J����  ͠����      C  , ,  �����  ����}  ϲ���}  ϲ����  �����      C  , ,  �p����  �p���}  ����}  �����  �p����      C  , ,  ������  �����}  ҂���}  ҂����  ������      C  , ,  ����Y  ����  �����  �����Y  ����Y      C  , ,  �����  ������  �j����  �j���  �����      C  , ,  �(���  �(����  ������  �����  �(���      C  , ,  �����  ������  �:����  �:���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �`���  �`����  �
����  �
���  �`���      C  , ,  �����  ������  �r����  �r���  �����      C  , ,  �0���  �0����  ������  �����  �0���      C  , ,  Ƙ���  Ƙ����  �B����  �B���  Ƙ���      C  , ,  � ���  � ����  Ȫ����  Ȫ���  � ���      C  , ,  �h���  �h����  �����  ����  �h���      C  , ,  �����  ������  �z����  �z���  �����      C  , ,  �8���  �8����  ������  �����  �8���      C  , ,  ͠���  ͠����  �J����  �J���  ͠���      C  , ,  ����  �����  ϲ����  ϲ���  ����      C  , ,  �p���  �p����  �����  ����  �p���      C  , ,  �����  ������  ҂����  ҂���  �����      C  , ,  �Z���Y  �Z���  ����  ����Y  �Z���Y      C  , ,  Ũ���Y  Ũ���  �R���  �R���Y  Ũ���Y      C  , ,  �����Y  �����  Ƞ���  Ƞ���Y  �����Y      C  , ,  �D���Y  �D���  �����  �����Y  �D���Y      C  , ,  ̒���Y  ̒���  �<���  �<���Y  ̒���Y      C  , ,  �����Y  �����  ϊ���  ϊ���Y  �����Y      C  , ,  �.���Y  �.���  �����  �����Y  �.���Y      C  , ,  �p����  �p����  �����  �����  �p����      C  , ,  ������  ������  �h����  �h����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �Z����  �Z����  �����  �����  �Z����      C  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      C  , ,  ������  ������  Ƞ����  Ƞ����  ������      C  , ,  �D����  �D����  ������  ������  �D����      C  , ,  ̒����  ̒����  �<����  �<����  ̒����      C  , ,  ������  ������  ϊ����  ϊ����  ������      C  , ,  �.����  �.����  ������  ������  �.����      C  , ,  �p����  �p���3  ����3  �����  �p����      C  , ,  ������  �����3  �h���3  �h����  ������      C  , ,  �����  ����3  �����3  ������  �����      C  , ,  �Z����  �Z���3  ����3  �����  �Z����      C  , ,  Ũ����  Ũ���3  �R���3  �R����  Ũ����      C  , ,  ������  �����3  Ƞ���3  Ƞ����  ������      C  , ,  �D����  �D���3  �����3  ������  �D����      C  , ,  ̒����  ̒���3  �<���3  �<����  ̒����      C  , ,  ������  �����3  ϊ���3  ϊ����  ������      C  , ,  �.����  �.���3  �����3  ������  �.����      C  , ,  �p���!  �p����  �����  ����!  �p���!      C  , ,  �����!  ������  �h����  �h���!  �����!      C  , ,  ����!  �����  ������  �����!  ����!      C  , ,  �Z���!  �Z����  �����  ����!  �Z���!      C  , ,  Ũ���!  Ũ����  �R����  �R���!  Ũ���!      C  , ,  �����!  ������  Ƞ����  Ƞ���!  �����!      C  , ,  �D���!  �D����  ������  �����!  �D���!      C  , ,  ̒���!  ̒����  �<����  �<���!  ̒���!      C  , ,  �����!  ������  ϊ����  ϊ���!  �����!      C  , ,  �.���!  �.����  ������  �����!  �.���!      C  , ,  �p����  �p���c  ����c  �����  �p����      C  , ,  ������  �����c  �h���c  �h����  ������      C  , ,  �����  ����c  �����c  ������  �����      C  , ,  �Z����  �Z���c  ����c  �����  �Z����      C  , ,  Ũ����  Ũ���c  �R���c  �R����  Ũ����      C  , ,  ������  �����c  Ƞ���c  Ƞ����  ������      C  , ,  �D����  �D���c  �����c  ������  �D����      C  , ,  ̒����  ̒���c  �<���c  �<����  ̒����      C  , ,  ������  �����c  ϊ���c  ϊ����  ������      C  , ,  �.����  �.���c  �����c  ������  �.����      C  , ,  �p���Y  �p���  ����  ����Y  �p���Y      C  , ,  ������  �����5  �j���5  �j����  ������      C  , ,  �(����  �(���5  �����5  ������  �(����      C  , ,  ������  �����5  �:���5  �:����  ������      C  , ,  ������  �����}  �h���}  �h����  ������      C  , ,  �����  ����}  �����}  ������  �����      C  , ,  �Z����  �Z���}  ����}  �����  �Z����      C  , ,  Ũ����  Ũ���}  �R���}  �R����  Ũ����      C  , ,  ������  �����}  Ƞ���}  Ƞ����  ������      C  , ,  �D����  �D���}  �����}  ������  �D����      C  , ,  ̒����  ̒���}  �<���}  �<����  ̒����      C  , ,  ������  �����}  ϊ���}  ϊ����  ������      C  , ,  �.����  �.���}  �����}  ������  �.����      C  , ,  �p���k  �p���  ����  ����k  �p���k      C  , ,  �����k  �����  �h���  �h���k  �����k      C  , ,  ����k  ����  �����  �����k  ����k      C  , ,  �Z���k  �Z���  ����  ����k  �Z���k      C  , ,  Ũ���k  Ũ���  �R���  �R���k  Ũ���k      C  , ,  �����k  �����  Ƞ���  Ƞ���k  �����k      C  , ,  �D���k  �D���  �����  �����k  �D���k      C  , ,  ̒���k  ̒���  �<���  �<���k  ̒���k      C  , ,  �����k  �����  ϊ���  ϊ���k  �����k      C  , ,  �.���k  �.���  �����  �����k  �.���k      C  , ,  �p����  �p����  �����  �����  �p����      C  , ,  ������  ������  �h����  �h����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �Z����  �Z����  �����  �����  �Z����      C  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      C  , ,  ������  ������  Ƞ����  Ƞ����  ������      C  , ,  �D����  �D����  ������  ������  �D����      C  , ,  ̒����  ̒����  �<����  �<����  ̒����      C  , ,  ������  ������  ϊ����  ϊ����  ������      C  , ,  �.����  �.����  ������  ������  �.����      C  , ,  �p���s  �p���  ����  ����s  �p���s      C  , ,  �����s  �����  �h���  �h���s  �����s      C  , ,  ����s  ����  �����  �����s  ����s      C  , ,  �Z���s  �Z���  ����  ����s  �Z���s      C  , ,  Ũ���s  Ũ���  �R���  �R���s  Ũ���s      C  , ,  �����s  �����  Ƞ���  Ƞ���s  �����s      C  , ,  �D���s  �D���  �����  �����s  �D���s      C  , ,  ̒���s  ̒���  �<���  �<���s  ̒���s      C  , ,  �����s  �����  ϊ���  ϊ���s  �����s      C  , ,  �.���s  �.���  �����  �����s  �.���s      C  , ,  �p���  �p����  �����  ����  �p���      C  , ,  �����  ������  �h����  �h���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �Z���  �Z����  �����  ����  �Z���      C  , ,  Ũ���  Ũ����  �R����  �R���  Ũ���      C  , ,  �����  ������  Ƞ����  Ƞ���  �����      C  , ,  �D���  �D����  ������  �����  �D���      C  , ,  ̒���  ̒����  �<����  �<���  ̒���      C  , ,  �����  ������  ϊ����  ϊ���  �����      C  , ,  �.���  �.����  ������  �����  �.���      C  , ,  �p����  �p���M  ����M  �����  �p����      C  , ,  ������  �����M  �h���M  �h����  ������      C  , ,  �����  ����M  �����M  ������  �����      C  , ,  �Z����  �Z���M  ����M  �����  �Z����      C  , ,  Ũ����  Ũ���M  �R���M  �R����  Ũ����      C  , ,  ������  �����M  Ƞ���M  Ƞ����  ������      C  , ,  �D����  �D���M  �����M  ������  �D����      C  , ,  ̒����  ̒���M  �<���M  �<����  ̒����      C  , ,  ������  �����M  ϊ���M  ϊ����  ������      C  , ,  �.����  �.���M  �����M  ������  �.����      C  , ,  �p���;  �p����  �����  ����;  �p���;      C  , ,  �����;  ������  �h����  �h���;  �����;      C  , ,  ����;  �����  ������  �����;  ����;      C  , ,  �Z���;  �Z����  �����  ����;  �Z���;      C  , ,  Ũ���;  Ũ����  �R����  �R���;  Ũ���;      C  , ,  �����;  ������  Ƞ����  Ƞ���;  �����;      C  , ,  �D���;  �D����  ������  �����;  �D���;      C  , ,  ̒���;  ̒����  �<����  �<���;  ̒���;      C  , ,  �����;  ������  ϊ����  ϊ���;  �����;      C  , ,  �.���;  �.����  ������  �����;  �.���;      C  , ,  �p����  �p���}  ����}  �����  �p����      C  , ,  �Z����  �Z���a  ����a  �����  �Z����      C  , ,  Ũ����  Ũ���a  �R���a  �R����  Ũ����      C  , ,  ������  �����a  Ƞ���a  Ƞ����  ������      C  , ,  �D����  �D���a  �����a  ������  �D����      C  , ,  ̒����  ̒���a  �<���a  �<����  ̒����      C  , ,  ������  �����a  ϊ���a  ϊ����  ������      C  , ,  �.����  �.���a  �����a  ������  �.����      C  , ,  �p���O  �p����  �����  ����O  �p���O      C  , ,  �����O  ������  �h����  �h���O  �����O      C  , ,  ����O  �����  ������  �����O  ����O      C  , ,  �Z���O  �Z����  �����  ����O  �Z���O      C  , ,  Ũ���O  Ũ����  �R����  �R���O  Ũ���O      C  , ,  �����O  ������  Ƞ����  Ƞ���O  �����O      C  , ,  �D���O  �D����  ������  �����O  �D���O      C  , ,  ̒���O  ̒����  �<����  �<���O  ̒���O      C  , ,  �����O  ������  ϊ����  ϊ���O  �����O      C  , ,  �.���O  �.����  ������  �����O  �.���O      C  , ,  �p����  �p����  �����  �����  �p����      C  , ,  ������  ������  �h����  �h����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �Z����  �Z����  �����  �����  �Z����      C  , ,  Ũ����  Ũ����  �R����  �R����  Ũ����      C  , ,  ������  ������  Ƞ����  Ƞ����  ������      C  , ,  �D����  �D����  ������  ������  �D����      C  , ,  ̒����  ̒����  �<����  �<����  ̒����      C  , ,  ������  ������  ϊ����  ϊ����  ������      C  , ,  �.����  �.����  ������  ������  �.����      C  , ,  �p���  �p����  �����  ����  �p���      C  , ,  �����  ������  �h����  �h���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �Z���  �Z����  �����  ����  �Z���      C  , ,  Ũ���  Ũ����  �R����  �R���  Ũ���      C  , ,  �����  ������  Ƞ����  Ƞ���  �����      C  , ,  �D���  �D����  ������  �����  �D���      C  , ,  ̒���  ̒����  �<����  �<���  ̒���      C  , ,  �����  ������  ϊ����  ϊ���  �����      C  , ,  �.���  �.����  ������  �����  �.���      C  , ,  ������  �����}  �A���}  �A����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �3����  �3���}  �����}  ������  �3����      C  , ,  ā����  ā���}  �+���}  �+����  ā����      C  , ,  ������  �����}  �y���}  �y����  ������      C  , ,  �����  ����}  �����}  ������  �����      C  , ,  �k����  �k���}  ����}  �����  �k����      C  , ,  ͹����  ͹���}  �c���}  �c����  ͹����      C  , ,  �����  ����}  б���}  б����  �����      C  , ,  ������  �����a  �A���a  �A����  ������      C  , ,  ������  �����a  �����a  ������  ������      C  , ,  �3����  �3���a  �����a  ������  �3����      C  , ,  ā����  ā���a  �+���a  �+����  ā����      C  , ,  ������  �����a  �y���a  �y����  ������      C  , ,  �����  ����a  �����a  ������  �����      C  , ,  �k����  �k���a  ����a  �����  �k����      C  , ,  ͹����  ͹���a  �c���a  �c����  ͹����      C  , ,  �����  ����a  б���a  б����  �����      C  , ,  �p����  �p���1  ����1  �����  �p����      C  , ,  ������  �����1  �h���1  �h����  ������      C  , ,  �����  ����1  �����1  ������  �����      C  , ,  �Z����  �Z���1  ����1  �����  �Z����      C  , ,  Ũ����  Ũ���1  �R���1  �R����  Ũ����      C  , ,  ������  �����1  Ƞ���1  Ƞ����  ������      C  , ,  �D����  �D���1  �����1  ������  �D����      C  , ,  ̒����  ̒���1  �<���1  �<����  ̒����      C  , ,  ������  �����1  ϊ���1  ϊ����  ������      C  , ,  �.����  �.���1  �����1  ������  �.����      C  , ,  �p���  �p����  �����  ����  �p���      C  , ,  �����  ������  �h����  �h���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �Z���  �Z����  �����  ����  �Z���      C  , ,  Ũ���  Ũ����  �R����  �R���  Ũ���      C  , ,  �����  ������  Ƞ����  Ƞ���  �����      C  , ,  �D���  �D����  ������  �����  �D���      C  , ,  ̒���  ̒����  �<����  �<���  ̒���      C  , ,  �����  ������  ϊ����  ϊ���  �����      C  , ,  �.���  �.����  ������  �����  �.���      C  , ,  �p����  �p���a  ����a  �����  �p����      C  , ,  ������  �����a  �h���a  �h����  ������      C  , ,  �����  ����a  �����a  ������  �����      C  , ,  ������  ������  ������  ������  ������      C  , ,  ������  �����k  �����k  ������  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  ������  �����a  �����a  ������  ������      C  , ,  ����Y  ����  �����  �����Y  ����Y      C  , ,  �����  �����  ������  ������  �����      C  , ,  �����  ����3  �����3  ������  �����      C  , ,  ����!  �����  ������  �����!  ����!      C  , ,  ����  �����  ������  �����  ����      C  , ,  �����  ����c  �����c  ������  �����      C  , ,  �����  �����  ������  ������  �����      C  , ,  �p����  �p���5  ����5  �����  �p����      C  , ,  �p����  �p���}  ����}  �����  �p����      C  , ,  �p���  �p����  �����  ����  �p���      C  , ,  �����  ����;  �����;  ������  �����      C  , ,  ����u  ����  �����  �����u  ����u      C  , ,  ����)  �����  ������  �����)  ����)      C  , ,  �����  ����k  �����k  ������  �����      C  , ,  �d���  �d����  �����  ����  �d���      C  , ,  �"���  �"����  ������  �����  �"���      C  , ,  �����  ������  �\����  �\���  �����      C  , ,  �d����  �d����  �����  �����  �d����      C  , ,  ������  ������  �\����  �\����  ������      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �N���  �N����  ������  �����  �N���      C  , ,  �"����  �"����  ������  ������  �"����      C  , ,  �=����  �=����  ������  ������  �=����      C  , ,  ������  ������  �5����  �5����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �����  ������  �F����  �F���  �����      C  , ,  �'����  �'����  ������  ������  �'����      C  , ,  �u����  �u����  �����  �����  �u����      C  , ,  ������  ������  �m����  �m����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �_����  �_����  �	����  �	����  �_����      C  , ,  ������  ������  �W����  �W����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �I����  �I����  ������  ������  �I����      C  , ,  �=����  �=���k  �����k  ������  �=����      C  , ,  ������  �����k  �5���k  �5����  ������      C  , ,  ������  �����k  �����k  ������  ������      C  , ,  �'����  �'���k  �����k  ������  �'����      C  , ,  �u����  �u���k  ����k  �����  �u����      C  , ,  ������  �����k  �m���k  �m����  ������      C  , ,  �����  ����k  �����k  ������  �����      C  , ,  �_����  �_���k  �	���k  �	����  �_����      C  , ,  ������  �����k  �W���k  �W����  ������      C  , ,  ������  �����k  �����k  ������  ������      C  , ,  �I����  �I���k  �����k  ������  �I����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �d����  �d���;  ����;  �����  �d����      C  , ,  ������  �����;  �\���;  �\����  ������      C  , ,  � ����  � ���;  �����;  ������  � ����      C  , ,  �N����  �N���;  �����;  ������  �N����      C  , ,  ������  �����;  �F���;  �F����  ������      C  , ,  ������  �����;  �����;  ������  ������      C  , ,  �8����  �8���;  �����;  ������  �8����      C  , ,  ������  �����;  �0���;  �0����  ������      C  , ,  ������  �����;  �~���;  �~����  ������      C  , ,  �"����  �"���;  �����;  ������  �"����      C  , ,  �8���  �8����  ������  �����  �8���      C  , ,  �����  ������  �0����  �0���  �����      C  , ,  �d���)  �d����  �����  ����)  �d���)      C  , ,  �����)  ������  �\����  �\���)  �����)      C  , ,  � ���)  � ����  ������  �����)  � ���)      C  , ,  �N���)  �N����  ������  �����)  �N���)      C  , ,  �����)  ������  �F����  �F���)  �����)      C  , ,  �����)  ������  ������  �����)  �����)      C  , ,  �8���)  �8����  ������  �����)  �8���)      C  , ,  �����)  ������  �0����  �0���)  �����)      C  , ,  �����)  ������  �~����  �~���)  �����)      C  , ,  �"���)  �"����  ������  �����)  �"���)      C  , ,  �d���u  �d���  ����  ����u  �d���u      C  , ,  �����u  �����  �\���  �\���u  �����u      C  , ,  � ���u  � ���  �����  �����u  � ���u      C  , ,  �N���u  �N���  �����  �����u  �N���u      C  , ,  �����u  �����  �F���  �F���u  �����u      C  , ,  �����u  �����  �����  �����u  �����u      C  , ,  �8���u  �8���  �����  �����u  �8���u      C  , ,  �����u  �����  �0���  �0���u  �����u      C  , ,  �����u  �����  �~���  �~���u  �����u      C  , ,  �"���u  �"���  �����  �����u  �"���u      C  , ,  �����  ������  �~����  �~���  �����      C  , ,  �d����  �d���k  ����k  �����  �d����      C  , ,  ������  �����k  �\���k  �\����  ������      C  , ,  � ����  � ���k  �����k  ������  � ����      C  , ,  �N����  �N���k  �����k  ������  �N����      C  , ,  ������  �����k  �F���k  �F����  ������      C  , ,  ������  �����k  �����k  ������  ������      C  , ,  �8����  �8���k  �����k  ������  �8����      C  , ,  ������  �����k  �0���k  �0����  ������      C  , ,  ������  �����k  �~���k  �~����  ������      C  , ,  �"����  �"���k  �����k  ������  �"����      C  , ,  �N����  �N����  ������  ������  �N����      C  , ,  ������  ������  �F����  �F����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �8����  �8����  ������  ������  �8����      C  , ,  ������  ������  �0����  �0����  ������      C  , ,  ������  ������  �~����  �~����  ������      C  , ,  �z����  �z����  �$����  �$����  �z����      C  , ,  ������  ������  �r����  �r����  ������      C  , ,  �����  ������  ������  �����  �����      C  , ,  �B���  �B����  ������  �����  �B���      C  , ,  �����  ������  �:����  �:���  �����      C  , ,  ������  ������  ������  ������  ������      C  , ,  �����  ������  ������  �����  �����      C  , ,  �,���  �,����  ������  �����  �,���      C  , ,  �X���u  �X���  ����  ����u  �X���u      C  , ,  �����u  �����  �P���  �P���u  �����u      C  , ,  �����u  �����  �����  �����u  �����u      C  , ,  �B���u  �B���  �����  �����u  �B���u      C  , ,  �����u  �����  �:���  �:���u  �����u      C  , ,  �����u  �����  �����  �����u  �����u      C  , ,  �,���u  �,���  �����  �����u  �,���u      C  , ,  �z���u  �z���  �$���  �$���u  �z���u      C  , ,  �����u  �����  �r���  �r���u  �����u      C  , ,  �z���  �z����  �$����  �$���  �z���      C  , ,  �
���)  �
����  ������  �����)  �
���)      C  , ,  �X���)  �X����  �����  ����)  �X���)      C  , ,  �����)  ������  �P����  �P���)  �����)      C  , ,  �����)  ������  ������  �����)  �����)      C  , ,  �B���)  �B����  ������  �����)  �B���)      C  , ,  �����)  ������  �:����  �:���)  �����)      C  , ,  �����)  ������  ������  �����)  �����)      C  , ,  �,���)  �,����  ������  �����)  �,���)      C  , ,  �z���)  �z����  �$����  �$���)  �z���)      C  , ,  �����)  ������  �r����  �r���)  �����)      C  , ,  �B����  �B����  ������  ������  �B����      C  , ,  �1����  �1���k  �����k  ������  �1����      C  , ,  �����  ����k  �)���k  �)����  �����      C  , ,  ������  �����k  �w���k  �w����  ������      C  , ,  �����  ����k  �����k  ������  �����      C  , ,  �i����  �i���k  ����k  �����  �i����      C  , ,  ������  �����k  �a���k  �a����  ������      C  , ,  �����  ����k  �����k  ������  �����      C  , ,  �S����  �S���k  �����k  ������  �S����      C  , ,  ������  �����k  �K���k  �K����  ������      C  , ,  ������  �����k  �����k  ������  ������      C  , ,  �����  ������  �r����  �r���  �����      C  , ,  �1����  �1����  ������  ������  �1����      C  , ,  �����  �����  �)����  �)����  �����      C  , ,  ������  ������  �w����  �w����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �i����  �i����  �����  �����  �i����      C  , ,  ������  ������  �a����  �a����  ������      C  , ,  �����  �����  ������  ������  �����      C  , ,  �S����  �S����  ������  ������  �S����      C  , ,  ������  ������  �K����  �K����  ������      C  , ,  �
����  �
���k  �����k  ������  �
����      C  , ,  �X����  �X���k  ����k  �����  �X����      C  , ,  ������  �����k  �P���k  �P����  ������      C  , ,  ������  �����k  �����k  ������  ������      C  , ,  �B����  �B���k  �����k  ������  �B����      C  , ,  ������  �����k  �:���k  �:����  ������      C  , ,  ������  �����k  �����k  ������  ������      C  , ,  �,����  �,���k  �����k  ������  �,����      C  , ,  �z����  �z���k  �$���k  �$����  �z����      C  , ,  ������  �����k  �r���k  �r����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �
���u  �
���  �����  �����u  �
���u      C  , ,  �
����  �
���;  �����;  ������  �
����      C  , ,  �X����  �X���;  ����;  �����  �X����      C  , ,  ������  �����;  �P���;  �P����  ������      C  , ,  ������  �����;  �����;  ������  ������      C  , ,  �B����  �B���;  �����;  ������  �B����      C  , ,  ������  �����;  �:���;  �:����  ������      C  , ,  ������  �����;  �����;  ������  ������      C  , ,  �,����  �,���;  �����;  ������  �,����      C  , ,  �z����  �z���;  �$���;  �$����  �z����      C  , ,  ������  �����;  �r���;  �r����  ������      C  , ,  ������  ������  �:����  �:����  ������      C  , ,  �
���  �
����  ������  �����  �
���      C  , ,  �X���  �X����  �����  ����  �X���      C  , ,  �����  ������  �P����  �P���  �����      C  , ,  �,����  �,����  ������  ������  �,����      C  , ,  �
����  �
����  ������  ������  �
����      C  , ,  �X����  �X����  �����  �����  �X����      C  , ,  ������  ������  �P����  �P����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  ������  �����5  �r���5  �r����  ������      C  , ,  ������  �����}  �r���}  �r����  ������      C  , ,  �����  ������  �r����  �r���  �����      C  , ,  �z����  �z���3  �$���3  �$����  �z����      C  , ,  ������  �����3  �r���3  �r����  ������      C  , ,  ������  �����3  �:���3  �:����  ������      C  , ,  ������  �����3  �����3  ������  ������      C  , ,  �����Y  �����  �:���  �:���Y  �����Y      C  , ,  �����Y  �����  �����  �����Y  �����Y      C  , ,  �,���Y  �,���  �����  �����Y  �,���Y      C  , ,  �z���Y  �z���  �$���  �$���Y  �z���Y      C  , ,  �����Y  �����  �r���  �r���Y  �����Y      C  , ,  �����!  ������  �:����  �:���!  �����!      C  , ,  �,����  �,���3  �����3  ������  �,����      C  , ,  �����!  ������  ������  �����!  �����!      C  , ,  �,���!  �,����  ������  �����!  �,���!      C  , ,  �z���!  �z����  �$����  �$���!  �z���!      C  , ,  �����!  ������  �r����  �r���!  �����!      C  , ,  ������  ������  �:����  �:����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �,����  �,����  ������  ������  �,����      C  , ,  �z����  �z����  �$����  �$����  �z����      C  , ,  ������  ������  �r����  �r����  ������      C  , ,  ������  �����c  �:���c  �:����  ������      C  , ,  ������  �����c  �����c  ������  ������      C  , ,  �,����  �,���c  �����c  ������  �,����      C  , ,  �z����  �z���c  �$���c  �$����  �z����      C  , ,  ������  �����c  �r���c  �r����  ������      C  , ,  ������  �����3  �����3  ������  ������      C  , ,  �B���Y  �B���  �����  �����Y  �B���Y      C  , ,  �
���Y  �
���  �����  �����Y  �
���Y      C  , ,  ������  ������  �P����  �P����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �B����  �B����  ������  ������  �B����      C  , ,  �
����  �
����  ������  ������  �
����      C  , ,  �X����  �X����  �����  �����  �X����      C  , ,  �
���!  �
����  ������  �����!  �
���!      C  , ,  �X���!  �X����  �����  ����!  �X���!      C  , ,  �����!  ������  �P����  �P���!  �����!      C  , ,  �X���Y  �X���  ����  ����Y  �X���Y      C  , ,  �
����  �
���3  �����3  ������  �
����      C  , ,  �X����  �X���3  ����3  �����  �X����      C  , ,  �
����  �
���c  �����c  ������  �
����      C  , ,  �X����  �X���c  ����c  �����  �X����      C  , ,  ������  �����c  �P���c  �P����  ������      C  , ,  ������  �����c  �����c  ������  ������      C  , ,  �B����  �B���c  �����c  ������  �B����      C  , ,  �����!  ������  ������  �����!  �����!      C  , ,  �B���!  �B����  ������  �����!  �B���!      C  , ,  �����Y  �����  �P���  �P���Y  �����Y      C  , ,  �B����  �B���3  �����3  ������  �B����      C  , ,  �����Y  �����  �����  �����Y  �����Y      C  , ,  ������  �����3  �P���3  �P����  ������      C  , ,  ������  �����5  �:���5  �:����  ������      C  , ,  ������  �����5  �����5  ������  ������      C  , ,  �`����  �`���5  �
���5  �
����  �`����      C  , ,  ������  �����5  �2���5  �2����  ������      C  , ,  ������  �����5  �����5  ������  ������      C  , ,  ������  �����}  �2���}  �2����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �X����  �X���}  ����}  �����  �X����      C  , ,  ������  �����}  �j���}  �j����  ������      C  , ,  �(����  �(���}  �����}  ������  �(����      C  , ,  ������  �����}  �:���}  �:����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �`����  �`���}  �
���}  �
����  �`����      C  , ,  �����  ������  �2����  �2���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �X���  �X����  �����  ����  �X���      C  , ,  �����  ������  �j����  �j���  �����      C  , ,  �(���  �(����  ������  �����  �(���      C  , ,  �����  ������  �:����  �:���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �`���  �`����  �
����  �
���  �`���      C  , ,  �X����  �X���5  ����5  �����  �X����      C  , ,  ������  �����5  �j���5  �j����  ������      C  , ,  �(����  �(���5  �����5  ������  �(����      C  , ,  � ����  � ���}  �����}  ������  � ����      C  , ,  �h����  �h���}  ����}  �����  �h����      C  , ,  ������  �����}  �z���}  �z����  ������      C  , ,  �8����  �8���}  �����}  ������  �8����      C  , ,  ������  �����}  �J���}  �J����  ������      C  , ,  �����  ����}  �����}  ������  �����      C  , ,  � ����  � ���5  �����5  ������  � ����      C  , ,  �h����  �h���5  ����5  �����  �h����      C  , ,  ������  �����5  �z���5  �z����  ������      C  , ,  �8����  �8���5  �����5  ������  �8����      C  , ,  ������  �����5  �J���5  �J����  ������      C  , ,  �����  ����5  �����5  ������  �����      C  , ,  �0����  �0���5  �����5  ������  �0����      C  , ,  ������  �����5  �B���5  �B����  ������      C  , ,  �0���  �0����  ������  �����  �0���      C  , ,  �����  ������  �B����  �B���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �h���  �h����  �����  ����  �h���      C  , ,  �����  ������  �z����  �z���  �����      C  , ,  �8���  �8����  ������  �����  �8���      C  , ,  �����  ������  �J����  �J���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �0����  �0���}  �����}  ������  �0����      C  , ,  ������  �����}  �B���}  �B����  ������      C  , ,  � ���Y  � ���  �����  �����Y  � ���Y      C  , ,  �N���Y  �N���  �����  �����Y  �N���Y      C  , ,  �d����  �d���c  ����c  �����  �d����      C  , ,  ������  �����c  �\���c  �\����  ������      C  , ,  � ����  � ���c  �����c  ������  � ����      C  , ,  �N����  �N���c  �����c  ������  �N����      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �@����  �@���}  �����}  ������  �@����      C  , ,  ������  �����}  �R���}  �R����  ������      C  , ,  �����  ����}  �����}  ������  �����      C  , ,  �x����  �x���}  �"���}  �"����  �x����      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �H����  �H���}  �����}  ������  �H����      C  , ,  ������  �����}  �Z���}  �Z����  ������      C  , ,  �����  ����}  �����}  ������  �����      C  , ,  ������  �����}  �*���}  �*����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �P����  �P���}  �����}  ������  �P����      C  , ,  ������  �����}  �b���}  �b����  ������      C  , ,  � ����  � ���}  �����}  ������  � ����      C  , ,  ������  �����}  �2���}  �2����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  ������  �����c  �F���c  �F����  ������      C  , ,  ������  �����c  �����c  ������  ������      C  , ,  �8����  �8���c  �����c  ������  �8����      C  , ,  ������  �����c  �0���c  �0����  ������      C  , ,  ������  �����c  �~���c  �~����  ������      C  , ,  �"����  �"���c  �����c  ������  �"����      C  , ,  �����Y  �����  �F���  �F���Y  �����Y      C  , ,  �����Y  �����  �����  �����Y  �����Y      C  , ,  �8���Y  �8���  �����  �����Y  �8���Y      C  , ,  �����Y  �����  �0���  �0���Y  �����Y      C  , ,  �����Y  �����  �~���  �~���Y  �����Y      C  , ,  �"���Y  �"���  �����  �����Y  �"���Y      C  , ,  �d���Y  �d���  ����  ����Y  �d���Y      C  , ,  �d����  �d����  �����  �����  �d����      C  , ,  �d����  �d���3  ����3  �����  �d����      C  , ,  �d���!  �d����  �����  ����!  �d���!      C  , ,  �����!  ������  �\����  �\���!  �����!      C  , ,  � ���!  � ����  ������  �����!  � ���!      C  , ,  �N���!  �N����  ������  �����!  �N���!      C  , ,  �����!  ������  �F����  �F���!  �����!      C  , ,  �����!  ������  ������  �����!  �����!      C  , ,  �8���!  �8����  ������  �����!  �8���!      C  , ,  �����!  ������  �0����  �0���!  �����!      C  , ,  �����!  ������  �~����  �~���!  �����!      C  , ,  �"���!  �"����  ������  �����!  �"���!      C  , ,  ������  �����3  �\���3  �\����  ������      C  , ,  � ����  � ���3  �����3  ������  � ����      C  , ,  �N����  �N���3  �����3  ������  �N����      C  , ,  ������  �����3  �F���3  �F����  ������      C  , ,  ������  �����3  �����3  ������  ������      C  , ,  �8����  �8���3  �����3  ������  �8����      C  , ,  ������  �����3  �0���3  �0����  ������      C  , ,  �����  ������  ������  �����  �����      C  , ,  �@���  �@����  ������  �����  �@���      C  , ,  �����  ������  �R����  �R���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �x���  �x����  �"����  �"���  �x���      C  , ,  �����  ������  ������  �����  �����      C  , ,  �H���  �H����  ������  �����  �H���      C  , ,  �����  ������  �Z����  �Z���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �����  ������  �*����  �*���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �P���  �P����  ������  �����  �P���      C  , ,  �����  ������  �b����  �b���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �����  ������  �2����  �2���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  ������  �����5  �����5  ������  ������      C  , ,  �@����  �@���5  �����5  ������  �@����      C  , ,  ������  �����5  �R���5  �R����  ������      C  , ,  �����  ����5  �����5  ������  �����      C  , ,  �x����  �x���5  �"���5  �"����  �x����      C  , ,  ������  �����5  �����5  ������  ������      C  , ,  �H����  �H���5  �����5  ������  �H����      C  , ,  ������  �����5  �Z���5  �Z����  ������      C  , ,  �����  ����5  �����5  ������  �����      C  , ,  ������  �����5  �*���5  �*����  ������      C  , ,  ������  �����5  �����5  ������  ������      C  , ,  �P����  �P���5  �����5  ������  �P����      C  , ,  ������  �����5  �b���5  �b����  ������      C  , ,  � ����  � ���5  �����5  ������  � ����      C  , ,  ������  �����5  �2���5  �2����  ������      C  , ,  ������  �����5  �����5  ������  ������      C  , ,  ������  �����3  �~���3  �~����  ������      C  , ,  �"����  �"���3  �����3  ������  �"����      C  , ,  ������  ������  �\����  �\����  ������      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  �N����  �N����  ������  ������  �N����      C  , ,  ������  ������  �F����  �F����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �8����  �8����  ������  ������  �8����      C  , ,  ������  ������  �0����  �0����  ������      C  , ,  ������  ������  �~����  �~����  ������      C  , ,  �"����  �"����  ������  ������  �"����      C  , ,  �����Y  �����  �\���  �\���Y  �����Y      C  , ,  r8���  r8����  r�����  r����  r8���      C  , ,  r8����  r8���5  r����5  r�����  r8����      C  , ,  r8����  r8���}  r����}  r�����  r8����      C  , ,  {����  {�����  |�����  |����  {����      C  , ,  ~6���  ~6����  ~�����  ~����  ~6���      C  , ,  �����  ������  �.����  �.���  �����      C  , ,  �����  ������  �|����  �|���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �n���  �n����  �����  ����  �n���      C  , ,  ������  ������  ������  ������  ������      C  , ,  �G����  �G����  ������  ������  �G����      C  , ,  ������  ������  �?����  �?����  ������      C  , ,  �����  ������  �f����  �f���  �����      C  , ,  t����  t�����  u�����  u����  t����      C  , ,  r����  r�����  sZ����  sZ���  r����      C  , ,  r����u  r����  sZ���  sZ���u  r����u      C  , ,  t����u  t����  u����  u����u  t����u      C  , ,  wL���u  wL���  w����  w����u  wL���u      C  , ,  s�����  s����k  t����k  t�����  s�����      C  , ,  v%����  v%���k  v����k  v�����  v%����      C  , ,  xs����  xs���k  y���k  y����  xs����      C  , ,  z�����  z����k  {k���k  {k����  z�����      C  , ,  }����  }���k  }����k  }�����  }����      C  , ,  ]����  ]���k  ����k  �����  ]����      C  , ,  ������  �����k  �U���k  �U����  ������      C  , ,  ������  �����k  �����k  ������  ������      C  , ,  �G����  �G���k  �����k  ������  �G����      C  , ,  ������  �����k  �?���k  �?����  ������      C  , ,  wL���  wL����  w�����  w����  wL���      C  , ,  y����u  y����  zD���  zD���u  y����u      C  , ,  {����u  {����  |����  |����u  {����u      C  , ,  ~6���u  ~6���  ~����  ~����u  ~6���u      C  , ,  �����u  �����  �.���  �.���u  �����u      C  , ,  �����u  �����  �|���  �|���u  �����u      C  , ,  � ���u  � ���  �����  �����u  � ���u      C  , ,  �n���u  �n���  ����  ����u  �n���u      C  , ,  �����u  �����  �f���  �f���u  �����u      C  , ,  r�����  r����;  sZ���;  sZ����  r�����      C  , ,  t�����  t����;  u����;  u�����  t�����      C  , ,  wL����  wL���;  w����;  w�����  wL����      C  , ,  y�����  y����;  zD���;  zD����  y�����      C  , ,  {�����  {����;  |����;  |�����  {�����      C  , ,  ~6����  ~6���;  ~����;  ~�����  ~6����      C  , ,  ������  �����;  �.���;  �.����  ������      C  , ,  ������  �����;  �|���;  �|����  ������      C  , ,  � ����  � ���;  �����;  ������  � ����      C  , ,  �n����  �n���;  ����;  �����  �n����      C  , ,  ������  �����;  �f���;  �f����  ������      C  , ,  r����)  r�����  sZ����  sZ���)  r����)      C  , ,  t����)  t�����  u�����  u����)  t����)      C  , ,  wL���)  wL����  w�����  w����)  wL���)      C  , ,  y����)  y�����  zD����  zD���)  y����)      C  , ,  {����)  {�����  |�����  |����)  {����)      C  , ,  ~6���)  ~6����  ~�����  ~����)  ~6���)      C  , ,  �����)  ������  �.����  �.���)  �����)      C  , ,  �����)  ������  �|����  �|���)  �����)      C  , ,  � ���)  � ����  ������  �����)  � ���)      C  , ,  �n���)  �n����  �����  ����)  �n���)      C  , ,  �����)  ������  �f����  �f���)  �����)      C  , ,  s�����  s�����  t�����  t�����  s�����      C  , ,  v%����  v%����  v�����  v�����  v%����      C  , ,  xs����  xs����  y����  y����  xs����      C  , ,  z�����  z�����  {k����  {k����  z�����      C  , ,  }����  }����  }�����  }�����  }����      C  , ,  ]����  ]����  �����  �����  ]����      C  , ,  ������  ������  �U����  �U����  ������      C  , ,  r�����  r����k  sZ���k  sZ����  r�����      C  , ,  t�����  t����k  u����k  u�����  t�����      C  , ,  wL����  wL���k  w����k  w�����  wL����      C  , ,  y�����  y����k  zD���k  zD����  y�����      C  , ,  {�����  {����k  |����k  |�����  {�����      C  , ,  ~6����  ~6���k  ~����k  ~�����  ~6����      C  , ,  ������  �����k  �.���k  �.����  ������      C  , ,  ������  �����k  �|���k  �|����  ������      C  , ,  � ����  � ���k  �����k  ������  � ����      C  , ,  �n����  �n���k  ����k  �����  �n����      C  , ,  ������  �����k  �f���k  �f����  ������      C  , ,  y����  y�����  zD����  zD���  y����      C  , ,  r�����  r�����  sZ����  sZ����  r�����      C  , ,  t�����  t�����  u�����  u�����  t�����      C  , ,  wL����  wL����  w�����  w�����  wL����      C  , ,  y�����  y�����  zD����  zD����  y�����      C  , ,  {�����  {�����  |�����  |�����  {�����      C  , ,  ~6����  ~6����  ~�����  ~�����  ~6����      C  , ,  ������  ������  �.����  �.����  ������      C  , ,  ������  ������  �|����  �|����  ������      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  �n����  �n����  �����  �����  �n����      C  , ,  ������  ������  �f����  �f����  ������      C  , ,  k����)  k�����  lp����  lp���)  k����)      C  , ,  n���)  n����  n�����  n����)  n���)      C  , ,  pb���)  pb����  q����  q���)  pb���)      C  , ,  pb���  pb����  q����  q���  pb���      C  , ,  ]����  ]�����  ^�����  ^����  ]����      C  , ,  ]����u  ]����  ^����  ^����u  ]����u      C  , ,  `@���u  `@���  `����  `����u  `@���u      C  , ,  d����u  d����  e����  e����u  d����u      C  , ,  g*���u  g*���  g����  g����u  g*���u      C  , ,  ix���u  ix���  j"���  j"���u  ix���u      C  , ,  k����u  k����  lp���  lp���u  k����u      C  , ,  n���u  n���  n����  n����u  n���u      C  , ,  pb���u  pb���  q���  q���u  pb���u      C  , ,  `@���  `@����  `�����  `����  `@���      C  , ,  b����u  b����  c8���  c8���u  b����u      C  , ,  _����  _����  _�����  _�����  _����      C  , ,  ag����  ag����  b����  b����  ag����      C  , ,  c�����  c�����  d_����  d_����  c�����      C  , ,  f����  f����  f�����  f�����  f����      C  , ,  hQ����  hQ����  h�����  h�����  hQ����      C  , ,  j�����  j�����  kI����  kI����  j�����      C  , ,  l�����  l�����  m�����  m�����  l�����      C  , ,  o;����  o;����  o�����  o�����  o;����      C  , ,  q�����  q�����  r3����  r3����  q�����      C  , ,  b����  b�����  c8����  c8���  b����      C  , ,  d����  d�����  e�����  e����  d����      C  , ,  _����  _���k  _����k  _�����  _����      C  , ,  ag����  ag���k  b���k  b����  ag����      C  , ,  ]�����  ]����;  ^����;  ^�����  ]�����      C  , ,  `@����  `@���;  `����;  `�����  `@����      C  , ,  b�����  b����;  c8���;  c8����  b�����      C  , ,  ]�����  ]����k  ^����k  ^�����  ]�����      C  , ,  `@����  `@���k  `����k  `�����  `@����      C  , ,  b�����  b����k  c8���k  c8����  b�����      C  , ,  d�����  d����k  e����k  e�����  d�����      C  , ,  g*����  g*���k  g����k  g�����  g*����      C  , ,  ix����  ix���k  j"���k  j"����  ix����      C  , ,  k�����  k����k  lp���k  lp����  k�����      C  , ,  n����  n���k  n����k  n�����  n����      C  , ,  pb����  pb���k  q���k  q����  pb����      C  , ,  d�����  d����;  e����;  e�����  d�����      C  , ,  g*����  g*���;  g����;  g�����  g*����      C  , ,  ix����  ix���;  j"���;  j"����  ix����      C  , ,  k�����  k����;  lp���;  lp����  k�����      C  , ,  n����  n���;  n����;  n�����  n����      C  , ,  pb����  pb���;  q���;  q����  pb����      C  , ,  c�����  c����k  d_���k  d_����  c�����      C  , ,  f����  f���k  f����k  f�����  f����      C  , ,  hQ����  hQ���k  h����k  h�����  hQ����      C  , ,  j�����  j����k  kI���k  kI����  j�����      C  , ,  l�����  l����k  m����k  m�����  l�����      C  , ,  o;����  o;���k  o����k  o�����  o;����      C  , ,  ]�����  ]�����  ^�����  ^�����  ]�����      C  , ,  `@����  `@����  `�����  `�����  `@����      C  , ,  b�����  b�����  c8����  c8����  b�����      C  , ,  d�����  d�����  e�����  e�����  d�����      C  , ,  g*����  g*����  g�����  g�����  g*����      C  , ,  ix����  ix����  j"����  j"����  ix����      C  , ,  k�����  k�����  lp����  lp����  k�����      C  , ,  n����  n����  n�����  n�����  n����      C  , ,  pb����  pb����  q����  q����  pb����      C  , ,  q�����  q����k  r3���k  r3����  q�����      C  , ,  g*���  g*����  g�����  g����  g*���      C  , ,  ix���  ix����  j"����  j"���  ix���      C  , ,  k����  k�����  lp����  lp���  k����      C  , ,  n���  n����  n�����  n����  n���      C  , ,  ]����)  ]�����  ^�����  ^����)  ]����)      C  , ,  `@���)  `@����  `�����  `����)  `@���)      C  , ,  b����)  b�����  c8����  c8���)  b����)      C  , ,  d����)  d�����  e�����  e����)  d����)      C  , ,  g*���)  g*����  g�����  g����)  g*���)      C  , ,  ix���)  ix����  j"����  j"���)  ix���)      C  , ,  p����  p�����  qz����  qz���  p����      C  , ,  d����Y  d����  e����  e����Y  d����Y      C  , ,  b�����  b����3  c8���3  c8����  b�����      C  , ,  d�����  d����3  e����3  e�����  d�����      C  , ,  g*����  g*���3  g����3  g�����  g*����      C  , ,  ix����  ix���3  j"���3  j"����  ix����      C  , ,  k�����  k����3  lp���3  lp����  k�����      C  , ,  n����  n���3  n����3  n�����  n����      C  , ,  _�����  _����5  `����5  `�����  _�����      C  , ,  aX����  aX���5  b���5  b����  aX����      C  , ,  b�����  b����5  cj���5  cj����  b�����      C  , ,  d(����  d(���5  d����5  d�����  d(����      C  , ,  e�����  e����5  f:���5  f:����  e�����      C  , ,  ix���!  ix����  j"����  j"���!  ix���!      C  , ,  k����!  k�����  lp����  lp���!  k����!      C  , ,  n���!  n����  n�����  n����!  n���!      C  , ,  pb���!  pb����  q����  q���!  pb���!      C  , ,  f�����  f����5  g����5  g�����  f�����      C  , ,  h`����  h`���5  i
���5  i
����  h`����      C  , ,  i�����  i����5  jr���5  jr����  i�����      C  , ,  k0����  k0���5  k����5  k�����  k0����      C  , ,  l�����  l����5  mB���5  mB����  l�����      C  , ,  n ����  n ���5  n����5  n�����  n ����      C  , ,  oh����  oh���5  p���5  p����  oh����      C  , ,  p�����  p����5  qz���5  qz����  p�����      C  , ,  pb����  pb���3  q���3  q����  pb����      C  , ,  g*���Y  g*���  g����  g����Y  g*���Y      C  , ,  ix���Y  ix���  j"���  j"���Y  ix���Y      C  , ,  k����Y  k����  lp���  lp���Y  k����Y      C  , ,  n���Y  n���  n����  n����Y  n���Y      C  , ,  pb���Y  pb���  q���  q���Y  pb���Y      C  , ,  ]����Y  ]����  ^����  ^����Y  ]����Y      C  , ,  ]�����  ]����3  ^����3  ^�����  ]�����      C  , ,  `@����  `@���3  `����3  `�����  `@����      C  , ,  ] ����  ] ���}  ]����}  ]�����  ] ����      C  , ,  ^�����  ^����}  _2���}  _2����  ^�����      C  , ,  _�����  _����}  `����}  `�����  _�����      C  , ,  aX����  aX���}  b���}  b����  aX����      C  , ,  b�����  b����}  cj���}  cj����  b�����      C  , ,  ]�����  ]����c  ^����c  ^�����  ]�����      C  , ,  ]�����  ]�����  ^�����  ^�����  ]�����      C  , ,  `@����  `@����  `�����  `�����  `@����      C  , ,  `@����  `@���c  `����c  `�����  `@����      C  , ,  b�����  b����c  c8���c  c8����  b�����      C  , ,  ] ����  ] ���5  ]����5  ]�����  ] ����      C  , ,  ^�����  ^����5  _2���5  _2����  ^�����      C  , ,  d�����  d����c  e����c  e�����  d�����      C  , ,  g*����  g*���c  g����c  g�����  g*����      C  , ,  ix����  ix���c  j"���c  j"����  ix����      C  , ,  k�����  k����c  lp���c  lp����  k�����      C  , ,  n����  n���c  n����c  n�����  n����      C  , ,  pb����  pb���c  q���c  q����  pb����      C  , ,  ] ���  ] ����  ]�����  ]����  ] ���      C  , ,  ^����  ^�����  _2����  _2���  ^����      C  , ,  _����  _�����  `�����  `����  _����      C  , ,  aX���  aX����  b����  b���  aX���      C  , ,  b����  b�����  cj����  cj���  b����      C  , ,  d(���  d(����  d�����  d����  d(���      C  , ,  e����  e�����  f:����  f:���  e����      C  , ,  d(����  d(���}  d����}  d�����  d(����      C  , ,  e�����  e����}  f:���}  f:����  e�����      C  , ,  f�����  f����}  g����}  g�����  f�����      C  , ,  h`����  h`���}  i
���}  i
����  h`����      C  , ,  i�����  i����}  jr���}  jr����  i�����      C  , ,  k0����  k0���}  k����}  k�����  k0����      C  , ,  l�����  l����}  mB���}  mB����  l�����      C  , ,  n ����  n ���}  n����}  n�����  n ����      C  , ,  oh����  oh���}  p���}  p����  oh����      C  , ,  p�����  p����}  qz���}  qz����  p�����      C  , ,  b�����  b�����  c8����  c8����  b�����      C  , ,  d�����  d�����  e�����  e�����  d�����      C  , ,  g*����  g*����  g�����  g�����  g*����      C  , ,  ix����  ix����  j"����  j"����  ix����      C  , ,  k�����  k�����  lp����  lp����  k�����      C  , ,  n����  n����  n�����  n�����  n����      C  , ,  pb����  pb����  q����  q����  pb����      C  , ,  `@���Y  `@���  `����  `����Y  `@���Y      C  , ,  b����Y  b����  c8���  c8���Y  b����Y      C  , ,  ]����!  ]�����  ^�����  ^����!  ]����!      C  , ,  `@���!  `@����  `�����  `����!  `@���!      C  , ,  b����!  b�����  c8����  c8���!  b����!      C  , ,  d����!  d�����  e�����  e����!  d����!      C  , ,  g*���!  g*����  g�����  g����!  g*���!      C  , ,  f����  f�����  g�����  g����  f����      C  , ,  h`���  h`����  i
����  i
���  h`���      C  , ,  i����  i�����  jr����  jr���  i����      C  , ,  k0���  k0����  k�����  k����  k0���      C  , ,  l����  l�����  mB����  mB���  l����      C  , ,  n ���  n ����  n�����  n����  n ���      C  , ,  oh���  oh����  p����  p���  oh���      C  , ,  ~6����  ~6���c  ~����c  ~�����  ~6����      C  , ,  ~6����  ~6����  ~�����  ~�����  ~6����      C  , ,  ~6����  ~6���3  ~����3  ~�����  ~6����      C  , ,  ~6���Y  ~6���  ~����  ~����Y  ~6���Y      C  , ,  ~6���!  ~6����  ~�����  ~����!  ~6���!      C  , ,  ������  �����c  �|���c  �|����  ������      C  , ,  � ����  � ���c  �����c  ������  � ����      C  , ,  �n����  �n���c  ����c  �����  �n����      C  , ,  ������  �����c  �f���c  �f����  ������      C  , ,  �n���Y  �n���  ����  ����Y  �n���Y      C  , ,  �����Y  �����  �f���  �f���Y  �����Y      C  , ,  � ���!  � ����  ������  �����!  � ���!      C  , ,  �n���!  �n����  �����  ����!  �n���!      C  , ,  �����Y  �����  �|���  �|���Y  �����Y      C  , ,  ������  ������  �.����  �.����  ������      C  , ,  ������  ������  �|����  �|����  ������      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  �n����  �n����  �����  �����  �n����      C  , ,  ������  ������  �f����  �f����  ������      C  , ,  �����!  ������  �f����  �f���!  �����!      C  , ,  � ���Y  � ���  �����  �����Y  � ���Y      C  , ,  ������  �����3  �.���3  �.����  ������      C  , ,  ������  �����3  �|���3  �|����  ������      C  , ,  � ����  � ���3  �����3  ������  � ����      C  , ,  �n����  �n���3  ����3  �����  �n����      C  , ,  ������  �����3  �f���3  �f����  ������      C  , ,  �����Y  �����  �.���  �.���Y  �����Y      C  , ,  ������  �����c  �.���c  �.����  ������      C  , ,  �����!  ������  �.����  �.���!  �����!      C  , ,  �����!  ������  �|����  �|���!  �����!      C  , ,  r����!  r�����  sZ����  sZ���!  r����!      C  , ,  t����!  t�����  u�����  u����!  t����!      C  , ,  wL���!  wL����  w�����  w����!  wL���!      C  , ,  y����!  y�����  zD����  zD���!  y����!      C  , ,  {����!  {�����  |�����  |����!  {����!      C  , ,  r����Y  r����  sZ���  sZ���Y  r����Y      C  , ,  t����Y  t����  u����  u����Y  t����Y      C  , ,  r�����  r����3  sZ���3  sZ����  r�����      C  , ,  t�����  t����3  u����3  u�����  t�����      C  , ,  wL����  wL���3  w����3  w�����  wL����      C  , ,  y�����  y����3  zD���3  zD����  y�����      C  , ,  {�����  {����3  |����3  |�����  {�����      C  , ,  wL����  wL���c  w����c  w�����  wL����      C  , ,  y�����  y����c  zD���c  zD����  y�����      C  , ,  {�����  {����c  |����c  |�����  {�����      C  , ,  r�����  r�����  sZ����  sZ����  r�����      C  , ,  t�����  t�����  u�����  u�����  t�����      C  , ,  wL����  wL����  w�����  w�����  wL����      C  , ,  wL���Y  wL���  w����  w����Y  wL���Y      C  , ,  y����Y  y����  zD���  zD���Y  y����Y      C  , ,  {����Y  {����  |����  |����Y  {����Y      C  , ,  y�����  y�����  zD����  zD����  y�����      C  , ,  {�����  {�����  |�����  |�����  {�����      C  , ,  r�����  r����c  sZ���c  sZ����  r�����      C  , ,  t�����  t����c  u����c  u�����  t�����      C  , ,  }x����  }x���}  ~"���}  ~"����  }x����      C  , ,  vp���  vp����  w����  w���  vp���      C  , ,  w����  w�����  x�����  x����  w����      C  , ,  y@���  y@����  y�����  y����  y@���      C  , ,  z����  z�����  {R����  {R���  z����      C  , ,  |���  |����  |�����  |����  |���      C  , ,  }x���  }x����  ~"����  ~"���  }x���      C  , ,  |����  |���5  |����5  |�����  |����      C  , ,  }x����  }x���5  ~"���5  ~"����  }x����      C  , ,  z�����  z����5  {R���5  {R����  z�����      C  , ,  s����  s�����  tJ����  tJ���  s����      C  , ,  u���  u����  u�����  u����  u���      C  , ,  s�����  s����}  tJ���}  tJ����  s�����      C  , ,  u����  u���}  u����}  u�����  u����      C  , ,  vp����  vp���}  w���}  w����  vp����      C  , ,  w�����  w����}  x����}  x�����  w�����      C  , ,  s�����  s����5  tJ���5  tJ����  s�����      C  , ,  u����  u���5  u����5  u�����  u����      C  , ,  vp����  vp���5  w���5  w����  vp����      C  , ,  w�����  w����5  x����5  x�����  w�����      C  , ,  y@����  y@���5  y����5  y�����  y@����      C  , ,  y@����  y@���}  y����}  y�����  y@����      C  , ,  z�����  z����}  {R���}  {R����  z�����      C  , ,  |����  |���}  |����}  |�����  |����      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �P����  �P���}  �����}  ������  �P����      C  , ,  ������  �����}  �b���}  �b����  ������      C  , ,  ������  �����5  �Z���5  �Z����  ������      C  , ,  �����  ����5  �����5  ������  �����      C  , ,  ������  �����5  �*���5  �*����  ������      C  , ,  ������  �����5  �����5  ������  ������      C  , ,  �P����  �P���5  �����5  ������  �P����      C  , ,  ������  �����5  �b���5  �b����  ������      C  , ,  � ����  � ���5  �����5  ������  � ����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �P���  �P����  ������  �����  �P���      C  , ,  �����  ������  �b����  �b���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  ~�����  ~����5  ����5  �����  ~�����      C  , ,  ~����  ~�����  �����  ����  ~����      C  , ,  �H���  �H����  ������  �����  �H���      C  , ,  �����  ������  �Z����  �Z���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �����  ������  �*����  �*���  �����      C  , ,  �H����  �H���5  �����5  ������  �H����      C  , ,  ~�����  ~����}  ����}  �����  ~�����      C  , ,  �H����  �H���}  �����}  ������  �H����      C  , ,  � ����  � ���}  �����}  ������  � ����      C  , ,  ������  �����}  �Z���}  �Z����  ������      C  , ,  �����  ����}  �����}  ������  �����      C  , ,  ������  �����}  �*���}  �*����  ������      C  , ,  t�����  t�����  u�����  u�����  t�����      C  , ,  wL����  wL����  w�����  w�����  wL����      C  , ,  r�����  r����M  sZ���M  sZ����  r�����      C  , ,  t�����  t����M  u����M  u�����  t�����      C  , ,  wL����  wL���M  w����M  w�����  wL����      C  , ,  y�����  y����M  zD���M  zD����  y�����      C  , ,  {�����  {����M  |����M  |�����  {�����      C  , ,  ~6����  ~6���M  ~����M  ~�����  ~6����      C  , ,  ������  �����M  �.���M  �.����  ������      C  , ,  ������  �����M  �|���M  �|����  ������      C  , ,  � ����  � ���M  �����M  ������  � ����      C  , ,  �n����  �n���M  ����M  �����  �n����      C  , ,  ������  �����M  �f���M  �f����  ������      C  , ,  r����s  r����  sZ���  sZ���s  r����s      C  , ,  t����s  t����  u����  u����s  t����s      C  , ,  wL���s  wL���  w����  w����s  wL���s      C  , ,  y����s  y����  zD���  zD���s  y����s      C  , ,  {����s  {����  |����  |����s  {����s      C  , ,  r����;  r�����  sZ����  sZ���;  r����;      C  , ,  t����;  t�����  u�����  u����;  t����;      C  , ,  wL���;  wL����  w�����  w����;  wL���;      C  , ,  y����;  y�����  zD����  zD���;  y����;      C  , ,  {����;  {�����  |�����  |����;  {����;      C  , ,  ~6���;  ~6����  ~�����  ~����;  ~6���;      C  , ,  �����;  ������  �.����  �.���;  �����;      C  , ,  �����;  ������  �|����  �|���;  �����;      C  , ,  � ���;  � ����  ������  �����;  � ���;      C  , ,  �n���;  �n����  �����  ����;  �n���;      C  , ,  �����;  ������  �f����  �f���;  �����;      C  , ,  ~6���s  ~6���  ~����  ~����s  ~6���s      C  , ,  �����s  �����  �.���  �.���s  �����s      C  , ,  �����s  �����  �|���  �|���s  �����s      C  , ,  � ���s  � ���  �����  �����s  � ���s      C  , ,  �n���s  �n���  ����  ����s  �n���s      C  , ,  �����s  �����  �f���  �f���s  �����s      C  , ,  y�����  y�����  zD����  zD����  y�����      C  , ,  {�����  {�����  |�����  |�����  {�����      C  , ,  ~6����  ~6����  ~�����  ~�����  ~6����      C  , ,  ������  ������  �.����  �.����  ������      C  , ,  r�����  r����}  sZ���}  sZ����  r�����      C  , ,  t�����  t����}  u����}  u�����  t�����      C  , ,  wL����  wL���}  w����}  w�����  wL����      C  , ,  y�����  y����}  zD���}  zD����  y�����      C  , ,  {�����  {����}  |����}  |�����  {�����      C  , ,  ~6����  ~6���}  ~����}  ~�����  ~6����      C  , ,  ������  �����}  �.���}  �.����  ������      C  , ,  ������  �����}  �|���}  �|����  ������      C  , ,  � ����  � ���}  �����}  ������  � ����      C  , ,  �n����  �n���}  ����}  �����  �n����      C  , ,  ������  �����}  �f���}  �f����  ������      C  , ,  ������  ������  �|����  �|����  ������      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  �n����  �n����  �����  �����  �n����      C  , ,  ������  ������  �f����  �f����  ������      C  , ,  r����k  r����  sZ���  sZ���k  r����k      C  , ,  t����k  t����  u����  u����k  t����k      C  , ,  wL���k  wL���  w����  w����k  wL���k      C  , ,  y����k  y����  zD���  zD���k  y����k      C  , ,  {����k  {����  |����  |����k  {����k      C  , ,  ~6���k  ~6���  ~����  ~����k  ~6���k      C  , ,  �����k  �����  �.���  �.���k  �����k      C  , ,  �����k  �����  �|���  �|���k  �����k      C  , ,  � ���k  � ���  �����  �����k  � ���k      C  , ,  �n���k  �n���  ����  ����k  �n���k      C  , ,  �����k  �����  �f���  �f���k  �����k      C  , ,  r����  r�����  sZ����  sZ���  r����      C  , ,  t����  t�����  u�����  u����  t����      C  , ,  wL���  wL����  w�����  w����  wL���      C  , ,  y����  y�����  zD����  zD���  y����      C  , ,  {����  {�����  |�����  |����  {����      C  , ,  ~6���  ~6����  ~�����  ~����  ~6���      C  , ,  �����  ������  �.����  �.���  �����      C  , ,  �����  ������  �|����  �|���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �n���  �n����  �����  ����  �n���      C  , ,  �����  ������  �f����  �f���  �����      C  , ,  r�����  r�����  sZ����  sZ����  r�����      C  , ,  d�����  d����M  e����M  e�����  d�����      C  , ,  g*����  g*���M  g����M  g�����  g*����      C  , ,  ix����  ix���M  j"���M  j"����  ix����      C  , ,  k�����  k����M  lp���M  lp����  k�����      C  , ,  b����;  b�����  c8����  c8���;  b����;      C  , ,  b�����  b�����  c8����  c8����  b�����      C  , ,  d�����  d�����  e�����  e�����  d�����      C  , ,  b����  b�����  c8����  c8���  b����      C  , ,  d����  d�����  e�����  e����  d����      C  , ,  g*���  g*����  g�����  g����  g*���      C  , ,  ix���  ix����  j"����  j"���  ix���      C  , ,  b����k  b����  c8���  c8���k  b����k      C  , ,  d����k  d����  e����  e����k  d����k      C  , ,  g*���k  g*���  g����  g����k  g*���k      C  , ,  ix���k  ix���  j"���  j"���k  ix���k      C  , ,  k����k  k����  lp���  lp���k  k����k      C  , ,  n���k  n���  n����  n����k  n���k      C  , ,  pb���k  pb���  q���  q���k  pb���k      C  , ,  d����;  d�����  e�����  e����;  d����;      C  , ,  g*���;  g*����  g�����  g����;  g*���;      C  , ,  ix���;  ix����  j"����  j"���;  ix���;      C  , ,  k����;  k�����  lp����  lp���;  k����;      C  , ,  n���;  n����  n�����  n����;  n���;      C  , ,  pb���;  pb����  q����  q���;  pb���;      C  , ,  b�����  b����}  c8���}  c8����  b�����      C  , ,  d�����  d����}  e����}  e�����  d�����      C  , ,  g*����  g*���}  g����}  g�����  g*����      C  , ,  ix����  ix���}  j"���}  j"����  ix����      C  , ,  k�����  k����}  lp���}  lp����  k�����      C  , ,  k����  k�����  lp����  lp���  k����      C  , ,  n���  n����  n�����  n����  n���      C  , ,  pb���  pb����  q����  q���  pb���      C  , ,  n����  n���}  n����}  n�����  n����      C  , ,  pb����  pb���}  q���}  q����  pb����      C  , ,  n����  n���M  n����M  n�����  n����      C  , ,  pb����  pb���M  q���M  q����  pb����      C  , ,  b����s  b����  c8���  c8���s  b����s      C  , ,  d����s  d����  e����  e����s  d����s      C  , ,  g*���s  g*���  g����  g����s  g*���s      C  , ,  ix���s  ix���  j"���  j"���s  ix���s      C  , ,  k����s  k����  lp���  lp���s  k����s      C  , ,  n���s  n���  n����  n����s  n���s      C  , ,  pb���s  pb���  q���  q���s  pb���s      C  , ,  g*����  g*����  g�����  g�����  g*����      C  , ,  ix����  ix����  j"����  j"����  ix����      C  , ,  k�����  k�����  lp����  lp����  k�����      C  , ,  n����  n����  n�����  n�����  n����      C  , ,  pb����  pb����  q����  q����  pb����      C  , ,  b�����  b����M  c8���M  c8����  b�����      C  , ,  pb���  pb����  q����  q���  pb���      C  , ,  l�����  l����}  m����}  m�����  l�����      C  , ,  o;����  o;���}  o����}  o�����  o;����      C  , ,  q�����  q����}  r3���}  r3����  q�����      C  , ,  ag����  ag���}  b���}  b����  ag����      C  , ,  c�����  c����}  d_���}  d_����  c�����      C  , ,  _����  _���a  _����a  _�����  _����      C  , ,  ag����  ag���a  b���a  b����  ag����      C  , ,  ]�����  ]����1  ^����1  ^�����  ]�����      C  , ,  `@����  `@���1  `����1  `�����  `@����      C  , ,  b�����  b����1  c8���1  c8����  b�����      C  , ,  ]�����  ]����a  ^����a  ^�����  ]�����      C  , ,  `@����  `@���a  `����a  `�����  `@����      C  , ,  b�����  b����a  c8���a  c8����  b�����      C  , ,  d�����  d����a  e����a  e�����  d�����      C  , ,  g*����  g*���a  g����a  g�����  g*����      C  , ,  ix����  ix���a  j"���a  j"����  ix����      C  , ,  k�����  k����a  lp���a  lp����  k�����      C  , ,  n����  n���a  n����a  n�����  n����      C  , ,  pb����  pb���a  q���a  q����  pb����      C  , ,  d�����  d����1  e����1  e�����  d�����      C  , ,  g*����  g*���1  g����1  g�����  g*����      C  , ,  ix����  ix���1  j"���1  j"����  ix����      C  , ,  k�����  k����1  lp���1  lp����  k�����      C  , ,  n����  n���1  n����1  n�����  n����      C  , ,  pb����  pb���1  q���1  q����  pb����      C  , ,  c�����  c����a  d_���a  d_����  c�����      C  , ,  f����  f���a  f����a  f�����  f����      C  , ,  hQ����  hQ���a  h����a  h�����  hQ����      C  , ,  j�����  j����a  kI���a  kI����  j�����      C  , ,  ]����O  ]�����  ^�����  ^����O  ]����O      C  , ,  `@���O  `@����  `�����  `����O  `@���O      C  , ,  b����O  b�����  c8����  c8���O  b����O      C  , ,  d����O  d�����  e�����  e����O  d����O      C  , ,  g*���O  g*����  g�����  g����O  g*���O      C  , ,  ix���O  ix����  j"����  j"���O  ix���O      C  , ,  k����O  k�����  lp����  lp���O  k����O      C  , ,  n���O  n����  n�����  n����O  n���O      C  , ,  pb���O  pb����  q����  q���O  pb���O      C  , ,  l�����  l����a  m����a  m�����  l�����      C  , ,  o;����  o;���a  o����a  o�����  o;����      C  , ,  q�����  q����a  r3���a  r3����  q�����      C  , ,  f����  f���}  f����}  f�����  f����      C  , ,  hQ����  hQ���}  h����}  h�����  hQ����      C  , ,  j�����  j����}  kI���}  kI����  j�����      C  , ,  ]����  ]�����  ^�����  ^����  ]����      C  , ,  `@���  `@����  `�����  `����  `@���      C  , ,  b����  b�����  c8����  c8���  b����      C  , ,  d����  d�����  e�����  e����  d����      C  , ,  ]�����  ]�����  ^�����  ^�����  ]�����      C  , ,  `@����  `@����  `�����  `�����  `@����      C  , ,  b�����  b�����  c8����  c8����  b�����      C  , ,  b����  b�����  c8����  c8���  b����      C  , ,  d����  d�����  e�����  e����  d����      C  , ,  g*���  g*����  g�����  g����  g*���      C  , ,  ix���  ix����  j"����  j"���  ix���      C  , ,  k����  k�����  lp����  lp���  k����      C  , ,  n���  n����  n�����  n����  n���      C  , ,  pb���  pb����  q����  q���  pb���      C  , ,  d�����  d�����  e�����  e�����  d�����      C  , ,  g*����  g*����  g�����  g�����  g*����      C  , ,  ix����  ix����  j"����  j"����  ix����      C  , ,  k�����  k�����  lp����  lp����  k�����      C  , ,  n����  n����  n�����  n�����  n����      C  , ,  pb����  pb����  q����  q����  pb����      C  , ,  g*���  g*����  g�����  g����  g*���      C  , ,  ix���  ix����  j"����  j"���  ix���      C  , ,  k����  k�����  lp����  lp���  k����      C  , ,  n���  n����  n�����  n����  n���      C  , ,  _����  _���}  _����}  _�����  _����      C  , ,  ������  ������  �f����  �f����  ������      C  , ,  v%����  v%���}  v����}  v�����  v%����      C  , ,  xs����  xs���}  y���}  y����  xs����      C  , ,  z�����  z����}  {k���}  {k����  z�����      C  , ,  }����  }���}  }����}  }�����  }����      C  , ,  r�����  r����a  sZ���a  sZ����  r�����      C  , ,  t�����  t����a  u����a  u�����  t�����      C  , ,  wL����  wL���a  w����a  w�����  wL����      C  , ,  y�����  y����a  zD���a  zD����  y�����      C  , ,  {�����  {����a  |����a  |�����  {�����      C  , ,  ~6����  ~6���a  ~����a  ~�����  ~6����      C  , ,  ������  �����a  �.���a  �.����  ������      C  , ,  ������  �����a  �|���a  �|����  ������      C  , ,  � ����  � ���a  �����a  ������  � ����      C  , ,  �n����  �n���a  ����a  �����  �n����      C  , ,  ������  �����a  �f���a  �f����  ������      C  , ,  ]����  ]���}  ����}  �����  ]����      C  , ,  ������  �����}  �U���}  �U����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �G����  �G���}  �����}  ������  �G����      C  , ,  s�����  s����a  t����a  t�����  s�����      C  , ,  v%����  v%���a  v����a  v�����  v%����      C  , ,  xs����  xs���a  y���a  y����  xs����      C  , ,  z�����  z����a  {k���a  {k����  z�����      C  , ,  }����  }���a  }����a  }�����  }����      C  , ,  ]����  ]���a  ����a  �����  ]����      C  , ,  ������  �����a  �U���a  �U����  ������      C  , ,  ������  �����a  �����a  ������  ������      C  , ,  r����  r�����  sZ����  sZ���  r����      C  , ,  t����  t�����  u�����  u����  t����      C  , ,  wL���  wL����  w�����  w����  wL���      C  , ,  y����  y�����  zD����  zD���  y����      C  , ,  {����  {�����  |�����  |����  {����      C  , ,  ~6���  ~6����  ~�����  ~����  ~6���      C  , ,  �����  ������  �.����  �.���  �����      C  , ,  r����O  r�����  sZ����  sZ���O  r����O      C  , ,  t����O  t�����  u�����  u����O  t����O      C  , ,  wL���O  wL����  w�����  w����O  wL���O      C  , ,  y����O  y�����  zD����  zD���O  y����O      C  , ,  {����O  {�����  |�����  |����O  {����O      C  , ,  ~6���O  ~6����  ~�����  ~����O  ~6���O      C  , ,  �����O  ������  �.����  �.���O  �����O      C  , ,  �����O  ������  �|����  �|���O  �����O      C  , ,  � ���O  � ����  ������  �����O  � ���O      C  , ,  �n���O  �n����  �����  ����O  �n���O      C  , ,  �����O  ������  �f����  �f���O  �����O      C  , ,  �����  ������  �|����  �|���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �n���  �n����  �����  ����  �n���      C  , ,  �����  ������  �f����  �f���  �����      C  , ,  �G����  �G���a  �����a  ������  �G����      C  , ,  r�����  r����1  sZ���1  sZ����  r�����      C  , ,  t�����  t����1  u����1  u�����  t�����      C  , ,  wL����  wL���1  w����1  w�����  wL����      C  , ,  y�����  y����1  zD���1  zD����  y�����      C  , ,  {�����  {����1  |����1  |�����  {�����      C  , ,  ~6����  ~6���1  ~����1  ~�����  ~6����      C  , ,  ������  �����1  �.���1  �.����  ������      C  , ,  ������  �����1  �|���1  �|����  ������      C  , ,  � ����  � ���1  �����1  ������  � ����      C  , ,  �n����  �n���1  ����1  �����  �n����      C  , ,  ������  �����1  �f���1  �f����  ������      C  , ,  ������  �����a  �?���a  �?����  ������      C  , ,  ������  �����}  �?���}  �?����  ������      C  , ,  r����  r�����  sZ����  sZ���  r����      C  , ,  t����  t�����  u�����  u����  t����      C  , ,  wL���  wL����  w�����  w����  wL���      C  , ,  y����  y�����  zD����  zD���  y����      C  , ,  {����  {�����  |�����  |����  {����      C  , ,  ~6���  ~6����  ~�����  ~����  ~6���      C  , ,  �����  ������  �.����  �.���  �����      C  , ,  �����  ������  �|����  �|���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �n���  �n����  �����  ����  �n���      C  , ,  �����  ������  �f����  �f���  �����      C  , ,  s�����  s����}  t����}  t�����  s�����      C  , ,  r�����  r�����  sZ����  sZ����  r�����      C  , ,  t�����  t�����  u�����  u�����  t�����      C  , ,  wL����  wL����  w�����  w�����  wL����      C  , ,  y�����  y�����  zD����  zD����  y�����      C  , ,  {�����  {�����  |�����  |�����  {�����      C  , ,  ~6����  ~6����  ~�����  ~�����  ~6����      C  , ,  ������  ������  �.����  �.����  ������      C  , ,  ������  ������  �|����  �|����  ������      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  �n����  �n����  �����  �����  �n����      C  , ,  �����  ����M  �����M  ������  �����      C  , ,  �����  ����1  �����1  ������  �����      C  , ,  ����k  ����  �����  �����k  ����k      C  , ,  ����  �����  ������  �����  ����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �����  ����a  �����a  ������  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  ����O  �����  ������  �����O  ����O      C  , ,  ����;  �����  ������  �����;  ����;      C  , ,  �����  �����  ������  ������  �����      C  , ,  ����s  ����  �����  �����s  ����s      C  , ,  �����  �����  ������  ������  �����      C  , ,  �����  ����}  �����}  ������  �����      C  , ,  �d���k  �d���  ����  ����k  �d���k      C  , ,  �����k  �����  �\���  �\���k  �����k      C  , ,  � ���k  � ���  �����  �����k  � ���k      C  , ,  �N���k  �N���  �����  �����k  �N���k      C  , ,  �����k  �����  �F���  �F���k  �����k      C  , ,  �����k  �����  �����  �����k  �����k      C  , ,  �8���k  �8���  �����  �����k  �8���k      C  , ,  �����k  �����  �0���  �0���k  �����k      C  , ,  �����k  �����  �~���  �~���k  �����k      C  , ,  ������  �����M  �\���M  �\����  ������      C  , ,  �"���k  �"���  �����  �����k  �"���k      C  , ,  � ����  � ���M  �����M  ������  � ����      C  , ,  �d���  �d����  �����  ����  �d���      C  , ,  �����  ������  �\����  �\���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �N����  �N���M  �����M  ������  �N����      C  , ,  ������  �����M  �F���M  �F����  ������      C  , ,  ������  �����M  �����M  ������  ������      C  , ,  �8����  �8���M  �����M  ������  �8����      C  , ,  �d���;  �d����  �����  ����;  �d���;      C  , ,  �����;  ������  �\����  �\���;  �����;      C  , ,  � ���;  � ����  ������  �����;  � ���;      C  , ,  �N���;  �N����  ������  �����;  �N���;      C  , ,  �����;  ������  �F����  �F���;  �����;      C  , ,  �����;  ������  ������  �����;  �����;      C  , ,  �8���;  �8����  ������  �����;  �8���;      C  , ,  �����;  ������  �0����  �0���;  �����;      C  , ,  �����;  ������  �~����  �~���;  �����;      C  , ,  �"���;  �"����  ������  �����;  �"���;      C  , ,  �N���  �N����  ������  �����  �N���      C  , ,  �����  ������  �F����  �F���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �8���  �8����  ������  �����  �8���      C  , ,  �����  ������  �0����  �0���  �����      C  , ,  �����  ������  �~����  �~���  �����      C  , ,  �"���  �"����  ������  �����  �"���      C  , ,  ������  �����M  �0���M  �0����  ������      C  , ,  ������  �����M  �~���M  �~����  ������      C  , ,  �d���s  �d���  ����  ����s  �d���s      C  , ,  �����s  �����  �\���  �\���s  �����s      C  , ,  � ���s  � ���  �����  �����s  � ���s      C  , ,  �N���s  �N���  �����  �����s  �N���s      C  , ,  �����s  �����  �F���  �F���s  �����s      C  , ,  �����s  �����  �����  �����s  �����s      C  , ,  �8���s  �8���  �����  �����s  �8���s      C  , ,  �����s  �����  �0���  �0���s  �����s      C  , ,  �����s  �����  �~���  �~���s  �����s      C  , ,  �"���s  �"���  �����  �����s  �"���s      C  , ,  �"����  �"���M  �����M  ������  �"����      C  , ,  �d����  �d����  �����  �����  �d����      C  , ,  ������  ������  �\����  �\����  ������      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  �d����  �d���M  ����M  �����  �d����      C  , ,  �d����  �d���}  ����}  �����  �d����      C  , ,  ������  �����}  �\���}  �\����  ������      C  , ,  � ����  � ���}  �����}  ������  � ����      C  , ,  �N����  �N���}  �����}  ������  �N����      C  , ,  ������  �����}  �F���}  �F����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �8����  �8���}  �����}  ������  �8����      C  , ,  ������  �����}  �0���}  �0����  ������      C  , ,  ������  �����}  �~���}  �~����  ������      C  , ,  �"����  �"���}  �����}  ������  �"����      C  , ,  �N����  �N����  ������  ������  �N����      C  , ,  ������  ������  �F����  �F����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �8����  �8����  ������  ������  �8����      C  , ,  ������  ������  �0����  �0����  ������      C  , ,  ������  ������  �~����  �~����  ������      C  , ,  �"����  �"����  ������  ������  �"����      C  , ,  �����k  �����  �:���  �:���k  �����k      C  , ,  �����k  �����  �����  �����k  �����k      C  , ,  �,���k  �,���  �����  �����k  �,���k      C  , ,  �
����  �
����  ������  ������  �
����      C  , ,  �X����  �X����  �����  �����  �X����      C  , ,  ������  ������  �P����  �P����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �B����  �B����  ������  ������  �B����      C  , ,  ������  ������  �:����  �:����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �
���s  �
���  �����  �����s  �
���s      C  , ,  �X���s  �X���  ����  ����s  �X���s      C  , ,  �����s  �����  �P���  �P���s  �����s      C  , ,  �����s  �����  �����  �����s  �����s      C  , ,  �,���s  �,���  �����  �����s  �,���s      C  , ,  �z���s  �z���  �$���  �$���s  �z���s      C  , ,  �B���s  �B���  �����  �����s  �B���s      C  , ,  �����s  �����  �r���  �r���s  �����s      C  , ,  �����s  �����  �:���  �:���s  �����s      C  , ,  �����s  �����  �����  �����s  �����s      C  , ,  �
���  �
����  ������  �����  �
���      C  , ,  �X���  �X����  �����  ����  �X���      C  , ,  �����  ������  �P����  �P���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �B���  �B����  ������  �����  �B���      C  , ,  �����  ������  �:����  �:���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �,���  �,����  ������  �����  �,���      C  , ,  �z���  �z����  �$����  �$���  �z���      C  , ,  �,����  �,����  ������  ������  �,����      C  , ,  �z����  �z����  �$����  �$����  �z����      C  , ,  ������  ������  �r����  �r����  ������      C  , ,  �����  ������  �r����  �r���  �����      C  , ,  �z���k  �z���  �$���  �$���k  �z���k      C  , ,  �����k  �����  �r���  �r���k  �����k      C  , ,  ������  �����M  �����M  ������  ������      C  , ,  �
����  �
���}  �����}  ������  �
����      C  , ,  �X����  �X���}  ����}  �����  �X����      C  , ,  ������  �����}  �P���}  �P����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �B����  �B���}  �����}  ������  �B����      C  , ,  ������  �����}  �:���}  �:����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �,����  �,���}  �����}  ������  �,����      C  , ,  �z����  �z���}  �$���}  �$����  �z����      C  , ,  ������  �����}  �r���}  �r����  ������      C  , ,  �,����  �,���M  �����M  ������  �,����      C  , ,  �z����  �z���M  �$���M  �$����  �z����      C  , ,  ������  �����M  �r���M  �r����  ������      C  , ,  �
���;  �
����  ������  �����;  �
���;      C  , ,  �X���;  �X����  �����  ����;  �X���;      C  , ,  �����;  ������  �P����  �P���;  �����;      C  , ,  �����;  ������  ������  �����;  �����;      C  , ,  �B���;  �B����  ������  �����;  �B���;      C  , ,  �����;  ������  �:����  �:���;  �����;      C  , ,  �����;  ������  ������  �����;  �����;      C  , ,  �,���;  �,����  ������  �����;  �,���;      C  , ,  �z���;  �z����  �$����  �$���;  �z���;      C  , ,  �����;  ������  �r����  �r���;  �����;      C  , ,  �
���k  �
���  �����  �����k  �
���k      C  , ,  �X���k  �X���  ����  ����k  �X���k      C  , ,  �����k  �����  �P���  �P���k  �����k      C  , ,  �����k  �����  �����  �����k  �����k      C  , ,  �B���k  �B���  �����  �����k  �B���k      C  , ,  �
����  �
���M  �����M  ������  �
����      C  , ,  �X����  �X���M  ����M  �����  �X����      C  , ,  ������  �����M  �P���M  �P����  ������      C  , ,  ������  �����M  �����M  ������  ������      C  , ,  �B����  �B���M  �����M  ������  �B����      C  , ,  ������  �����M  �:���M  �:����  ������      C  , ,  �i����  �i���}  ����}  �����  �i����      C  , ,  ������  �����}  �a���}  �a����  ������      C  , ,  �����  ����}  �����}  ������  �����      C  , ,  �S����  �S���}  �����}  ������  �S����      C  , ,  ������  �����}  �K���}  �K����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �
����  �
����  ������  ������  �
����      C  , ,  �X����  �X����  �����  �����  �X����      C  , ,  ������  ������  �P����  �P����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �B����  �B����  ������  ������  �B����      C  , ,  ������  ������  �:����  �:����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �,����  �,����  ������  ������  �,����      C  , ,  �z����  �z����  �$����  �$����  �z����      C  , ,  ������  ������  �r����  �r����  ������      C  , ,  �����  ������  �P����  �P���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �B���  �B����  ������  �����  �B���      C  , ,  �����  ������  �:����  �:���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �,���  �,����  ������  �����  �,���      C  , ,  �z���  �z����  �$����  �$���  �z���      C  , ,  �����  ������  �r����  �r���  �����      C  , ,  �X���  �X����  �����  ����  �X���      C  , ,  �����  ������  �P����  �P���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �B���  �B����  ������  �����  �B���      C  , ,  �����  ������  �:����  �:���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �,���  �,����  ������  �����  �,���      C  , ,  �z���  �z����  �$����  �$���  �z���      C  , ,  �����  ������  �r����  �r���  �����      C  , ,  �X����  �X���1  ����1  �����  �X����      C  , ,  ������  �����1  �P���1  �P����  ������      C  , ,  �
���O  �
����  ������  �����O  �
���O      C  , ,  �X���O  �X����  �����  ����O  �X���O      C  , ,  �����O  ������  �P����  �P���O  �����O      C  , ,  �����O  ������  ������  �����O  �����O      C  , ,  �B���O  �B����  ������  �����O  �B���O      C  , ,  �����O  ������  �:����  �:���O  �����O      C  , ,  �����O  ������  ������  �����O  �����O      C  , ,  �,���O  �,����  ������  �����O  �,���O      C  , ,  �z���O  �z����  �$����  �$���O  �z���O      C  , ,  �����O  ������  �r����  �r���O  �����O      C  , ,  ������  �����1  �����1  ������  ������      C  , ,  �1����  �1���a  �����a  ������  �1����      C  , ,  �����  ����a  �)���a  �)����  �����      C  , ,  ������  �����a  �w���a  �w����  ������      C  , ,  �����  ����a  �����a  ������  �����      C  , ,  �i����  �i���a  ����a  �����  �i����      C  , ,  ������  �����a  �a���a  �a����  ������      C  , ,  �����  ����a  �����a  ������  �����      C  , ,  �S����  �S���a  �����a  ������  �S����      C  , ,  ������  �����a  �K���a  �K����  ������      C  , ,  ������  �����a  �����a  ������  ������      C  , ,  �B����  �B���1  �����1  ������  �B����      C  , ,  ������  �����1  �:���1  �:����  ������      C  , ,  ������  �����1  �����1  ������  ������      C  , ,  �,����  �,���1  �����1  ������  �,����      C  , ,  �z����  �z���1  �$���1  �$����  �z����      C  , ,  ������  �����1  �r���1  �r����  ������      C  , ,  �
����  �
���1  �����1  ������  �
����      C  , ,  �
���  �
����  ������  �����  �
���      C  , ,  �
����  �
���a  �����a  ������  �
����      C  , ,  �X����  �X���a  ����a  �����  �X����      C  , ,  ������  �����a  �P���a  �P����  ������      C  , ,  ������  �����a  �����a  ������  ������      C  , ,  �B����  �B���a  �����a  ������  �B����      C  , ,  ������  �����a  �:���a  �:����  ������      C  , ,  ������  �����a  �����a  ������  ������      C  , ,  �,����  �,���a  �����a  ������  �,����      C  , ,  �z����  �z���a  �$���a  �$����  �z����      C  , ,  ������  �����a  �r���a  �r����  ������      C  , ,  �
���  �
����  ������  �����  �
���      C  , ,  �X���  �X����  �����  ����  �X���      C  , ,  �1����  �1���}  �����}  ������  �1����      C  , ,  �����  ����}  �)���}  �)����  �����      C  , ,  ������  �����}  �w���}  �w����  ������      C  , ,  �����  ����}  �����}  ������  �����      C  , ,  �'����  �'���}  �����}  ������  �'����      C  , ,  �u����  �u���}  ����}  �����  �u����      C  , ,  ������  �����}  �m���}  �m����  ������      C  , ,  �����  ����}  �����}  ������  �����      C  , ,  �_����  �_���}  �	���}  �	����  �_����      C  , ,  ������  �����}  �W���}  �W����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  �I����  �I���}  �����}  ������  �I����      C  , ,  �����O  ������  �\����  �\���O  �����O      C  , ,  � ���O  � ����  ������  �����O  � ���O      C  , ,  �N���O  �N����  ������  �����O  �N���O      C  , ,  �����O  ������  �F����  �F���O  �����O      C  , ,  �����O  ������  ������  �����O  �����O      C  , ,  �8���O  �8����  ������  �����O  �8���O      C  , ,  �����O  ������  �0����  �0���O  �����O      C  , ,  �����O  ������  �~����  �~���O  �����O      C  , ,  �"���O  �"����  ������  �����O  �"���O      C  , ,  �N����  �N���1  �����1  ������  �N����      C  , ,  ������  �����1  �F���1  �F����  ������      C  , ,  ������  �����1  �����1  ������  ������      C  , ,  �8����  �8���1  �����1  ������  �8����      C  , ,  ������  �����1  �0���1  �0����  ������      C  , ,  ������  �����1  �~���1  �~����  ������      C  , ,  �"����  �"���1  �����1  ������  �"����      C  , ,  �d����  �d���1  ����1  �����  �d����      C  , ,  �d���  �d����  �����  ����  �d���      C  , ,  �d���  �d����  �����  ����  �d���      C  , ,  �����  ������  �\����  �\���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �N���  �N����  ������  �����  �N���      C  , ,  �����  ������  �F����  �F���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �8���  �8����  ������  �����  �8���      C  , ,  �����  ������  �0����  �0���  �����      C  , ,  �����  ������  �~����  �~���  �����      C  , ,  �"���  �"����  ������  �����  �"���      C  , ,  �����  ������  �\����  �\���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �N���  �N����  ������  �����  �N���      C  , ,  �����  ������  �F����  �F���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �8���  �8����  ������  �����  �8���      C  , ,  �����  ������  �0����  �0���  �����      C  , ,  �����  ������  �~����  �~���  �����      C  , ,  �"���  �"����  ������  �����  �"���      C  , ,  ������  �����1  �\���1  �\����  ������      C  , ,  �d����  �d���a  ����a  �����  �d����      C  , ,  �=����  �=���a  �����a  ������  �=����      C  , ,  ������  �����a  �5���a  �5����  ������      C  , ,  ������  �����a  �����a  ������  ������      C  , ,  �'����  �'���a  �����a  ������  �'����      C  , ,  �u����  �u���a  ����a  �����  �u����      C  , ,  ������  �����a  �m���a  �m����  ������      C  , ,  �����  ����a  �����a  ������  �����      C  , ,  �_����  �_���a  �	���a  �	����  �_����      C  , ,  ������  �����a  �W���a  �W����  ������      C  , ,  ������  �����a  �����a  ������  ������      C  , ,  �I����  �I���a  �����a  ������  �I����      C  , ,  ������  �����a  �\���a  �\����  ������      C  , ,  � ����  � ���a  �����a  ������  � ����      C  , ,  �N����  �N���a  �����a  ������  �N����      C  , ,  ������  �����a  �F���a  �F����  ������      C  , ,  ������  �����a  �����a  ������  ������      C  , ,  �8����  �8���a  �����a  ������  �8����      C  , ,  ������  �����a  �0���a  �0����  ������      C  , ,  ������  �����a  �~���a  �~����  ������      C  , ,  �"����  �"���a  �����a  ������  �"����      C  , ,  � ����  � ���1  �����1  ������  � ����      C  , ,  �d���O  �d����  �����  ����O  �d���O      C  , ,  �d����  �d����  �����  �����  �d����      C  , ,  ������  ������  �\����  �\����  ������      C  , ,  � ����  � ����  ������  ������  � ����      C  , ,  �N����  �N����  ������  ������  �N����      C  , ,  ������  ������  �F����  �F����  ������      C  , ,  ������  ������  ������  ������  ������      C  , ,  �8����  �8����  ������  ������  �8����      C  , ,  ������  ������  �0����  �0����  ������      C  , ,  ������  ������  �~����  �~����  ������      C  , ,  �"����  �"����  ������  ������  �"����      C  , ,  �=����  �=���}  �����}  ������  �=����      C  , ,  ������  �����}  �5���}  �5����  ������      C  , ,  ������  �����}  �����}  ������  ������      C  , ,  ����f1  ����f�  ����f�  ����f1  ����f1      C  , ,  ����d  ����d�  ����d�  ����d  ����d      C  , ,  ����  �����  ������  �����  ����      C  , ,  �����  ����Y  �����Y  ������  �����      C  , ,  ���r  ���r�  ����r�  ����r  ���r      C  , ,  ���p�  ���qN  ����qN  ����p�  ���p�      C  , ,  ���o<  ���o�  ����o�  ����o<  ���o<      C  , ,  ���m�  ���n~  ����n~  ����m�  ���m�      C  , ,  ���ll  ���m  ����m  ����ll  ���ll      C  , ,  ���k  ���k�  ����k�  ����k  ���k      C  , ,  ���i�  ���jF  ����jF  ����i�  ���i�      C  , ,  �����  ������  �~����  �~���  �����      C  , ,  �"���  �"����  ������  �����  �"���      C  , ,  �d���  �d����  �����  ����  �d���      C  , ,  �d����  �d���Y  ����Y  �����  �d����      C  , ,  ������  �����Y  �\���Y  �\����  ������      C  , ,  � ����  � ���Y  �����Y  ������  � ����      C  , ,  �N����  �N���Y  �����Y  ������  �N����      C  , ,  ������  �����Y  �F���Y  �F����  ������      C  , ,  ������  �����Y  �����Y  ������  ������      C  , ,  �8����  �8���Y  �����Y  ������  �8����      C  , ,  ������  �����Y  �0���Y  �0����  ������      C  , ,  ������  �����Y  �~���Y  �~����  ������      C  , ,  �"����  �"���Y  �����Y  ������  �"����      C  , ,  �����  ������  �\����  �\���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �N���  �N����  ������  �����  �N���      C  , ,  �����  ������  �F����  �F���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �8���  �8����  ������  �����  �8���      C  , ,  �����  ������  �0����  �0���  �����      C  , ,  �
����  �
���Y  �����Y  ������  �
����      C  , ,  �X����  �X���Y  ����Y  �����  �X����      C  , ,  ������  �����Y  �P���Y  �P����  ������      C  , ,  ������  �����Y  �����Y  ������  ������      C  , ,  �B����  �B���Y  �����Y  ������  �B����      C  , ,  ������  �����Y  �:���Y  �:����  ������      C  , ,  ������  �����Y  �����Y  ������  ������      C  , ,  �,����  �,���Y  �����Y  ������  �,����      C  , ,  �z����  �z���Y  �$���Y  �$����  �z����      C  , ,  ������  �����Y  �r���Y  �r����  ������      C  , ,  �����  ������  �r����  �r���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  �,���  �,����  ������  �����  �,���      C  , ,  �z���  �z����  �$����  �$���  �z���      C  , ,  �B���  �B����  ������  �����  �B���      C  , ,  �����  ������  �:����  �:���  �����      C  , ,  �
���  �
����  ������  �����  �
���      C  , ,  �X���  �X����  �����  ����  �X���      C  , ,  �����  ������  �P����  �P���  �����      C  , ,  �����  ������  ������  �����  �����      C  , ,  ���p�  ���qN  ����qN  ����p�  ���p�      C  , ,  �V��p�  �V��qN  � ��qN  � ��p�  �V��p�      C  , ,  ����p�  ����qN  �t��qN  �t��p�  ����p�      C  , ,  ���p�  ���qN  ����qN  ����p�  ���p�      C  , ,  �f��p�  �f��qN  ���qN  ���p�  �f��p�      C  , ,  ����p�  ����qN  �^��qN  �^��p�  ����p�      C  , ,  �l��r  �l��r�  ���r�  ���r  �l��r      C  , ,  ���o<  ���o�  ����o�  ����o<  ���o<      C  , ,  �l��o<  �l��o�  ���o�  ���o<  �l��o<      C  , ,  ����o<  ����o�  �d��o�  �d��o<  ����o<      C  , ,  ���o<  ���o�  ����o�  ����o<  ���o<      C  , ,  �V��o<  �V��o�  � ��o�  � ��o<  �V��o<      C  , ,  ����o<  ����o�  �t��o�  �t��o<  ����o<      C  , ,  ���o<  ���o�  ����o�  ����o<  ���o<      C  , ,  �f��o<  �f��o�  ���o�  ���o<  �f��o<      C  , ,  ����o<  ����o�  �^��o�  �^��o<  ����o<      C  , ,  ����r  ����r�  �d��r�  �d��r  ����r      C  , ,  ���m�  ���n~  ����n~  ����m�  ���m�      C  , ,  �l��m�  �l��n~  ���n~  ���m�  �l��m�      C  , ,  ����m�  ����n~  �d��n~  �d��m�  ����m�      C  , ,  ���m�  ���n~  ����n~  ����m�  ���m�      C  , ,  �V��m�  �V��n~  � ��n~  � ��m�  �V��m�      C  , ,  ����m�  ����n~  �t��n~  �t��m�  ����m�      C  , ,  ���m�  ���n~  ����n~  ����m�  ���m�      C  , ,  �f��m�  �f��n~  ���n~  ���m�  �f��m�      C  , ,  ����m�  ����n~  �^��n~  �^��m�  ����m�      C  , ,  ���r  ���r�  ����r�  ����r  ���r      C  , ,  ���ll  ���m  ����m  ����ll  ���ll      C  , ,  �l��ll  �l��m  ���m  ���ll  �l��ll      C  , ,  ����ll  ����m  �d��m  �d��ll  ����ll      C  , ,  ���ll  ���m  ����m  ����ll  ���ll      C  , ,  �V��ll  �V��m  � ��m  � ��ll  �V��ll      C  , ,  ����ll  ����m  �t��m  �t��ll  ����ll      C  , ,  ���ll  ���m  ����m  ����ll  ���ll      C  , ,  �f��ll  �f��m  ���m  ���ll  �f��ll      C  , ,  ����ll  ����m  �^��m  �^��ll  ����ll      C  , ,  �V��r  �V��r�  � ��r�  � ��r  �V��r      C  , ,  ���k  ���k�  ����k�  ����k  ���k      C  , ,  �l��k  �l��k�  ���k�  ���k  �l��k      C  , ,  ����k  ����k�  �d��k�  �d��k  ����k      C  , ,  ���k  ���k�  ����k�  ����k  ���k      C  , ,  �V��k  �V��k�  � ��k�  � ��k  �V��k      C  , ,  ����k  ����k�  �t��k�  �t��k  ����k      C  , ,  ���k  ���k�  ����k�  ����k  ���k      C  , ,  �f��k  �f��k�  ���k�  ���k  �f��k      C  , ,  ����k  ����k�  �^��k�  �^��k  ����k      C  , ,  ����r  ����r�  �t��r�  �t��r  ����r      C  , ,  ���i�  ���jF  ����jF  ����i�  ���i�      C  , ,  �l��i�  �l��jF  ���jF  ���i�  �l��i�      C  , ,  ����i�  ����jF  �d��jF  �d��i�  ����i�      C  , ,  ���i�  ���jF  ����jF  ����i�  ���i�      C  , ,  �V��i�  �V��jF  � ��jF  � ��i�  �V��i�      C  , ,  ����i�  ����jF  �t��jF  �t��i�  ����i�      C  , ,  ���i�  ���jF  ����jF  ����i�  ���i�      C  , ,  �f��i�  �f��jF  ���jF  ���i�  �f��i�      C  , ,  ����i�  ����jF  �^��jF  �^��i�  ����i�      C  , ,  ���r  ���r�  ����r�  ����r  ���r      C  , ,  �f��r  �f��r�  ���r�  ���r  �f��r      C  , ,  ����r  ����r�  �^��r�  �^��r  ����r      C  , ,  ���r  ���r�  ����r�  ����r  ���r      C  , ,  ���p�  ���qN  ����qN  ����p�  ���p�      C  , ,  �l��p�  �l��qN  ���qN  ���p�  �l��p�      C  , ,  ����p�  ����qN  �d��qN  �d��p�  ����p�      C  , ,  �$��m�  �$��n~  ����n~  ����m�  �$��m�      C  , ,  �r��m�  �r��n~  ���n~  ���m�  �r��m�      C  , ,  ����m�  ����n~  �j��n~  �j��m�  ����m�      C  , ,  ���m�  ���n~  ����n~  ����m�  ���m�      C  , ,  �P��r  �P��r�  ����r�  ����r  �P��r      C  , ,  ����r  ����r�  �H��r�  �H��r  ����r      C  , ,  ����r  ����r�  ����r�  ����r  ����r      C  , ,  �:��r  �:��r�  ����r�  ����r  �:��r      C  , ,  ����r  ����r�  �2��r�  �2��r  ����r      C  , ,  ����r  ����r�  ����r�  ����r  ����r      C  , ,  �$��r  �$��r�  ����r�  ����r  �$��r      C  , ,  �r��r  �r��r�  ���r�  ���r  �r��r      C  , ,  ����r  ����r�  �j��r�  �j��r  ����r      C  , ,  ���r  ���r�  ����r�  ����r  ���r      C  , ,  �P��ll  �P��m  ����m  ����ll  �P��ll      C  , ,  ����ll  ����m  �H��m  �H��ll  ����ll      C  , ,  ����ll  ����m  ����m  ����ll  ����ll      C  , ,  �:��ll  �:��m  ����m  ����ll  �:��ll      C  , ,  ����ll  ����m  �2��m  �2��ll  ����ll      C  , ,  ����ll  ����m  ����m  ����ll  ����ll      C  , ,  �$��ll  �$��m  ����m  ����ll  �$��ll      C  , ,  �r��ll  �r��m  ���m  ���ll  �r��ll      C  , ,  ����ll  ����m  �j��m  �j��ll  ����ll      C  , ,  ���ll  ���m  ����m  ����ll  ���ll      C  , ,  �P��o<  �P��o�  ����o�  ����o<  �P��o<      C  , ,  ����o<  ����o�  �H��o�  �H��o<  ����o<      C  , ,  ����o<  ����o�  ����o�  ����o<  ����o<      C  , ,  �:��o<  �:��o�  ����o�  ����o<  �:��o<      C  , ,  ����o<  ����o�  �2��o�  �2��o<  ����o<      C  , ,  ����o<  ����o�  ����o�  ����o<  ����o<      C  , ,  �$��o<  �$��o�  ����o�  ����o<  �$��o<      C  , ,  �r��o<  �r��o�  ���o�  ���o<  �r��o<      C  , ,  ����o<  ����o�  �j��o�  �j��o<  ����o<      C  , ,  ���o<  ���o�  ����o�  ����o<  ���o<      C  , ,  �P��k  �P��k�  ����k�  ����k  �P��k      C  , ,  ����k  ����k�  �H��k�  �H��k  ����k      C  , ,  ����k  ����k�  ����k�  ����k  ����k      C  , ,  �:��k  �:��k�  ����k�  ����k  �:��k      C  , ,  ����k  ����k�  �2��k�  �2��k  ����k      C  , ,  ����k  ����k�  ����k�  ����k  ����k      C  , ,  �$��k  �$��k�  ����k�  ����k  �$��k      C  , ,  �r��k  �r��k�  ���k�  ���k  �r��k      C  , ,  ����k  ����k�  �j��k�  �j��k  ����k      C  , ,  ���k  ���k�  ����k�  ����k  ���k      C  , ,  �P��p�  �P��qN  ����qN  ����p�  �P��p�      C  , ,  ����p�  ����qN  �H��qN  �H��p�  ����p�      C  , ,  ����p�  ����qN  ����qN  ����p�  ����p�      C  , ,  �:��p�  �:��qN  ����qN  ����p�  �:��p�      C  , ,  ����p�  ����qN  �2��qN  �2��p�  ����p�      C  , ,  ����p�  ����qN  ����qN  ����p�  ����p�      C  , ,  �$��p�  �$��qN  ����qN  ����p�  �$��p�      C  , ,  �r��p�  �r��qN  ���qN  ���p�  �r��p�      C  , ,  ����p�  ����qN  �j��qN  �j��p�  ����p�      C  , ,  ���p�  ���qN  ����qN  ����p�  ���p�      C  , ,  �P��i�  �P��jF  ����jF  ����i�  �P��i�      C  , ,  ����i�  ����jF  �H��jF  �H��i�  ����i�      C  , ,  ����i�  ����jF  ����jF  ����i�  ����i�      C  , ,  �:��i�  �:��jF  ����jF  ����i�  �:��i�      C  , ,  ����i�  ����jF  �2��jF  �2��i�  ����i�      C  , ,  ����i�  ����jF  ����jF  ����i�  ����i�      C  , ,  �$��i�  �$��jF  ����jF  ����i�  �$��i�      C  , ,  �r��i�  �r��jF  ���jF  ���i�  �r��i�      C  , ,  ����i�  ����jF  �j��jF  �j��i�  ����i�      C  , ,  ���i�  ���jF  ����jF  ����i�  ���i�      C  , ,  �P��m�  �P��n~  ����n~  ����m�  �P��m�      C  , ,  ����m�  ����n~  �H��n~  �H��m�  ����m�      C  , ,  ����m�  ����n~  ����n~  ����m�  ����m�      C  , ,  �:��m�  �:��n~  ����n~  ����m�  �:��m�      C  , ,  ����m�  ����n~  �2��n~  �2��m�  ����m�      C  , ,  ����m�  ����n~  ����n~  ����m�  ����m�      C  , ,  y�����  y����Y  zD���Y  zD����  y�����      C  , ,  {�����  {����Y  |����Y  |�����  {�����      C  , ,  ~6����  ~6���Y  ~����Y  ~�����  ~6����      C  , ,  ������  �����Y  �.���Y  �.����  ������      C  , ,  ������  �����Y  �|���Y  �|����  ������      C  , ,  � ����  � ���Y  �����Y  ������  � ����      C  , ,  �n����  �n���Y  ����Y  �����  �n����      C  , ,  ������  �����Y  �f���Y  �f����  ������      C  , ,  r�����  r����Y  sZ���Y  sZ����  r�����      C  , ,  t�����  t����Y  u����Y  u�����  t�����      C  , ,  wL����  wL���Y  w����Y  w�����  wL����      C  , ,  r����  r�����  sZ����  sZ���  r����      C  , ,  t����  t�����  u�����  u����  t����      C  , ,  wL���  wL����  w�����  w����  wL���      C  , ,  y����  y�����  zD����  zD���  y����      C  , ,  {����  {�����  |�����  |����  {����      C  , ,  ~6���  ~6����  ~�����  ~����  ~6���      C  , ,  �����  ������  �.����  �.���  �����      C  , ,  �����  ������  �|����  �|���  �����      C  , ,  � ���  � ����  ������  �����  � ���      C  , ,  �n���  �n����  �����  ����  �n���      C  , ,  �����  ������  �f����  �f���  �����      C  , ,  ]����  ]�����  ^�����  ^����  ]����      C  , ,  g*���  g*����  g�����  g����  g*���      C  , ,  `@���  `@����  `�����  `����  `@���      C  , ,  d����  d�����  e�����  e����  d����      C  , ,  k����  k�����  lp����  lp���  k����      C  , ,  n���  n����  n�����  n����  n���      C  , ,  pb���  pb����  q����  q���  pb���      C  , ,  b����  b�����  c8����  c8���  b����      C  , ,  ix���  ix����  j"����  j"���  ix���      C  , ,  `@����  `@���Y  `����Y  `�����  `@����      C  , ,  b�����  b����Y  c8���Y  c8����  b�����      C  , ,  d�����  d����Y  e����Y  e�����  d�����      C  , ,  g*����  g*���Y  g����Y  g�����  g*����      C  , ,  ix����  ix���Y  j"���Y  j"����  ix����      C  , ,  k�����  k����Y  lp���Y  lp����  k�����      C  , ,  n����  n���Y  n����Y  n�����  n����      C  , ,  pb����  pb���Y  q���Y  q����  pb����      C  , ,  ]�����  ]����Y  ^����Y  ^�����  ]�����      C  , ,  ����p�  ����qN  �z��qN  �z��p�  ����p�      C  , ,  w`��r  w`��r�  x
��r�  x
��r  w`��r      C  , ,  ����o<  ����o�  �z��o�  �z��o<  ����o<      C  , ,  w`��m�  w`��n~  x
��n~  x
��m�  w`��m�      C  , ,  y���m�  y���n~  zX��n~  zX��m�  y���m�      C  , ,  {���m�  {���n~  |���n~  |���m�  {���m�      C  , ,  ~J��m�  ~J��n~  ~���n~  ~���m�  ~J��m�      C  , ,  ����m�  ����n~  �B��n~  �B��m�  ����m�      C  , ,  ����m�  ����n~  ����n~  ����m�  ����m�      C  , ,  �4��m�  �4��n~  ����n~  ����m�  �4��m�      C  , ,  ����m�  ����n~  �,��n~  �,��m�  ����m�      C  , ,  ����m�  ����n~  �z��n~  �z��m�  ����m�      C  , ,  y���r  y���r�  zX��r�  zX��r  y���r      C  , ,  �4��ll  �4��m  ����m  ����ll  �4��ll      C  , ,  w`��i�  w`��jF  x
��jF  x
��i�  w`��i�      C  , ,  y���i�  y���jF  zX��jF  zX��i�  y���i�      C  , ,  {���i�  {���jF  |���jF  |���i�  {���i�      C  , ,  ~J��i�  ~J��jF  ~���jF  ~���i�  ~J��i�      C  , ,  ����i�  ����jF  �B��jF  �B��i�  ����i�      C  , ,  ����i�  ����jF  ����jF  ����i�  ����i�      C  , ,  �4��i�  �4��jF  ����jF  ����i�  �4��i�      C  , ,  ����i�  ����jF  �,��jF  �,��i�  ����i�      C  , ,  ����i�  ����jF  �z��jF  �z��i�  ����i�      C  , ,  {���r  {���r�  |���r�  |���r  {���r      C  , ,  ~J��r  ~J��r�  ~���r�  ~���r  ~J��r      C  , ,  ����r  ����r�  �B��r�  �B��r  ����r      C  , ,  ����r  ����r�  ����r�  ����r  ����r      C  , ,  �4��r  �4��r�  ����r�  ����r  �4��r      C  , ,  ����r  ����r�  �,��r�  �,��r  ����r      C  , ,  ����r  ����r�  �z��r�  �z��r  ����r      C  , ,  ����ll  ����m  �,��m  �,��ll  ����ll      C  , ,  ����ll  ����m  �z��m  �z��ll  ����ll      C  , ,  w`��o<  w`��o�  x
��o�  x
��o<  w`��o<      C  , ,  y���o<  y���o�  zX��o�  zX��o<  y���o<      C  , ,  {���o<  {���o�  |���o�  |���o<  {���o<      C  , ,  ~J��o<  ~J��o�  ~���o�  ~���o<  ~J��o<      C  , ,  ����o<  ����o�  �B��o�  �B��o<  ����o<      C  , ,  ����o<  ����o�  ����o�  ����o<  ����o<      C  , ,  �4��o<  �4��o�  ����o�  ����o<  �4��o<      C  , ,  w`��p�  w`��qN  x
��qN  x
��p�  w`��p�      C  , ,  ����o<  ����o�  �,��o�  �,��o<  ����o<      C  , ,  w`��k  w`��k�  x
��k�  x
��k  w`��k      C  , ,  y���k  y���k�  zX��k�  zX��k  y���k      C  , ,  {���k  {���k�  |���k�  |���k  {���k      C  , ,  ~J��k  ~J��k�  ~���k�  ~���k  ~J��k      C  , ,  w`��ll  w`��m  x
��m  x
��ll  w`��ll      C  , ,  ����k  ����k�  �B��k�  �B��k  ����k      C  , ,  ����k  ����k�  ����k�  ����k  ����k      C  , ,  y���ll  y���m  zX��m  zX��ll  y���ll      C  , ,  �4��k  �4��k�  ����k�  ����k  �4��k      C  , ,  ����k  ����k�  �,��k�  �,��k  ����k      C  , ,  ����k  ����k�  �z��k�  �z��k  ����k      C  , ,  y���p�  y���qN  zX��qN  zX��p�  y���p�      C  , ,  {���p�  {���qN  |���qN  |���p�  {���p�      C  , ,  ~J��p�  ~J��qN  ~���qN  ~���p�  ~J��p�      C  , ,  ����p�  ����qN  �B��qN  �B��p�  ����p�      C  , ,  ����p�  ����qN  ����qN  ����p�  ����p�      C  , ,  �4��p�  �4��qN  ����qN  ����p�  �4��p�      C  , ,  ����p�  ����qN  �,��qN  �,��p�  ����p�      C  , ,  {���ll  {���m  |���m  |���ll  {���ll      C  , ,  ~J��ll  ~J��m  ~���m  ~���ll  ~J��ll      C  , ,  ����ll  ����m  �B��m  �B��ll  ����ll      C  , ,  ����ll  ����m  ����m  ����ll  ����ll      C  , ,  r���[
  r���[�  sn��[�  sn��[
  r���[
      C  , ,  u��[
  u��[�  u���[�  u���[
  u��[
      C  , ,  w`��[
  w`��[�  x
��[�  x
��[
  w`��[
      C  , ,  y���[
  y���[�  zX��[�  zX��[
  y���[
      C  , ,  {���[
  {���[�  |���[�  |���[
  {���[
      C  , ,  ~J��[
  ~J��[�  ~���[�  ~���[
  ~J��[
      C  , ,  ����[
  ����[�  �B��[�  �B��[
  ����[
      C  , ,  ����[
  ����[�  ����[�  ����[
  ����[
      C  , ,  �4��[
  �4��[�  ����[�  ����[
  �4��[
      C  , ,  ����[
  ����[�  �,��[�  �,��[
  ����[
      C  , ,  ����[
  ����[�  �z��[�  �z��[
  ����[
      C  , ,  ���d  ���d�  ����d�  ����d  ���d      C  , ,  �[��d  �[��d�  ���d�  ���d  �[��d      C  , ,  ����d  ����d�  �S��d�  �S��d  ����d      C  , ,  ����h4  ����h�  �B��h�  �B��h4  ����h4      C  , ,  ����h4  ����h�  ����h�  ����h4  ����h4      C  , ,  r���b  r���b�  sn��b�  sn��b  r���b      C  , ,  u��b  u��b�  u���b�  u���b  u��b      C  , ,  w`��b  w`��b�  x
��b�  x
��b  w`��b      C  , ,  y���b  y���b�  zX��b�  zX��b  y���b      C  , ,  {���b  {���b�  |���b�  |���b  {���b      C  , ,  ~J��b  ~J��b�  ~���b�  ~���b  ~J��b      C  , ,  ����b  ����b�  �B��b�  �B��b  ����b      C  , ,  ����b  ����b�  ����b�  ����b  ����b      C  , ,  �4��b  �4��b�  ����b�  ����b  �4��b      C  , ,  ����b  ����b�  �,��b�  �,��b  ����b      C  , ,  ����b  ����b�  �z��b�  �z��b  ����b      C  , ,  �4��h4  �4��h�  ����h�  ����h4  �4��h4      C  , ,  r���`�  r���aT  sn��aT  sn��`�  r���`�      C  , ,  u��`�  u��aT  u���aT  u���`�  u��`�      C  , ,  w`��`�  w`��aT  x
��aT  x
��`�  w`��`�      C  , ,  y���`�  y���aT  zX��aT  zX��`�  y���`�      C  , ,  {���`�  {���aT  |���aT  |���`�  {���`�      C  , ,  ~J��`�  ~J��aT  ~���aT  ~���`�  ~J��`�      C  , ,  ����`�  ����aT  �B��aT  �B��`�  ����`�      C  , ,  ����`�  ����aT  ����aT  ����`�  ����`�      C  , ,  �4��`�  �4��aT  ����aT  ����`�  �4��`�      C  , ,  ����`�  ����aT  �,��aT  �,��`�  ����`�      C  , ,  ����`�  ����aT  �z��aT  �z��`�  ����`�      C  , ,  r���_B  r���_�  sn��_�  sn��_B  r���_B      C  , ,  u��_B  u��_�  u���_�  u���_B  u��_B      C  , ,  w`��_B  w`��_�  x
��_�  x
��_B  w`��_B      C  , ,  y���_B  y���_�  zX��_�  zX��_B  y���_B      C  , ,  {���_B  {���_�  |���_�  |���_B  {���_B      C  , ,  ~J��_B  ~J��_�  ~���_�  ~���_B  ~J��_B      C  , ,  ����_B  ����_�  �B��_�  �B��_B  ����_B      C  , ,  ����_B  ����_�  ����_�  ����_B  ����_B      C  , ,  �4��_B  �4��_�  ����_�  ����_B  �4��_B      C  , ,  ����_B  ����_�  �,��_�  �,��_B  ����_B      C  , ,  ����_B  ����_�  �z��_�  �z��_B  ����_B      C  , ,  r���]�  r���^�  sn��^�  sn��]�  r���]�      C  , ,  u��]�  u��^�  u���^�  u���]�  u��]�      C  , ,  w`��]�  w`��^�  x
��^�  x
��]�  w`��]�      C  , ,  y���]�  y���^�  zX��^�  zX��]�  y���]�      C  , ,  {���]�  {���^�  |���^�  |���]�  {���]�      C  , ,  ~J��]�  ~J��^�  ~���^�  ~���]�  ~J��]�      C  , ,  ����]�  ����^�  �B��^�  �B��]�  ����]�      C  , ,  ����]�  ����^�  ����^�  ����]�  ����]�      C  , ,  �4��]�  �4��^�  ����^�  ����]�  �4��]�      C  , ,  ����]�  ����^�  �,��^�  �,��]�  ����]�      C  , ,  ����]�  ����^�  �z��^�  �z��]�  ����]�      C  , ,  r���\r  r���]  sn��]  sn��\r  r���\r      C  , ,  u��\r  u��]  u���]  u���\r  u��\r      C  , ,  w`��\r  w`��]  x
��]  x
��\r  w`��\r      C  , ,  y���\r  y���]  zX��]  zX��\r  y���\r      C  , ,  {���\r  {���]  |���]  |���\r  {���\r      C  , ,  ~J��\r  ~J��]  ~���]  ~���\r  ~J��\r      C  , ,  ����\r  ����]  �B��]  �B��\r  ����\r      C  , ,  ����\r  ����]  ����]  ����\r  ����\r      C  , ,  �4��\r  �4��]  ����]  ����\r  �4��\r      C  , ,  ����\r  ����]  �,��]  �,��\r  ����\r      C  , ,  ����\r  ����]  �z��]  �z��\r  ����\r      C  , ,  ����h4  ����h�  �,��h�  �,��h4  ����h4      C  , ,  ����f1  ����f�  �S��f�  �S��f1  ����f1      C  , ,  y���h4  y���h�  zX��h�  zX��h4  y���h4      C  , ,  {���h4  {���h�  |���h�  |���h4  {���h4      C  , ,  ~J��h4  ~J��h�  ~���h�  ~���h4  ~J��h4      C  , ,  s���d  s���d�  t���d�  t���d  s���d      C  , ,  v9��d  v9��d�  v���d�  v���d  v9��d      C  , ,  x���d  x���d�  y1��d�  y1��d  x���d      C  , ,  z���d  z���d�  {��d�  {��d  z���d      C  , ,  }#��d  }#��d�  }���d�  }���d  }#��d      C  , ,  q��d  q��d�  ���d�  ���d  q��d      C  , ,  ����d  ����d�  �i��d�  �i��d  ����d      C  , ,  ����h4  ����h�  �z��h�  �z��h4  ����h4      C  , ,  w`��h4  w`��h�  x
��h�  x
��h4  w`��h4      C  , ,  s���f1  s���f�  t���f�  t���f1  s���f1      C  , ,  v9��f1  v9��f�  v���f�  v���f1  v9��f1      C  , ,  x���f1  x���f�  y1��f�  y1��f1  x���f1      C  , ,  z���f1  z���f�  {��f�  {��f1  z���f1      C  , ,  }#��f1  }#��f�  }���f�  }���f1  }#��f1      C  , ,  q��f1  q��f�  ���f�  ���f1  q��f1      C  , ,  ����f1  ����f�  �i��f�  �i��f1  ����f1      C  , ,  ���f1  ���f�  ����f�  ����f1  ���f1      C  , ,  �[��f1  �[��f�  ���f�  ���f1  �[��f1      C  , ,  ����Y�  ����ZL  �z��ZL  �z��Y�  ����Y�      C  , ,  r���Y�  r���ZL  sn��ZL  sn��Y�  r���Y�      C  , ,  r���X:  r���X�  sn��X�  sn��X:  r���X:      C  , ,  u��X:  u��X�  u���X�  u���X:  u��X:      C  , ,  w`��X:  w`��X�  x
��X�  x
��X:  w`��X:      C  , ,  y���X:  y���X�  zX��X�  zX��X:  y���X:      C  , ,  {���X:  {���X�  |���X�  |���X:  {���X:      C  , ,  ~J��X:  ~J��X�  ~���X�  ~���X:  ~J��X:      C  , ,  ����X:  ����X�  �B��X�  �B��X:  ����X:      C  , ,  ����X:  ����X�  ����X�  ����X:  ����X:      C  , ,  �4��X:  �4��X�  ����X�  ����X:  �4��X:      C  , ,  ����X:  ����X�  �,��X�  �,��X:  ����X:      C  , ,  ����X:  ����X�  �z��X�  �z��X:  ����X:      C  , ,  u��Y�  u��ZL  u���ZL  u���Y�  u��Y�      C  , ,  w`��Y�  w`��ZL  x
��ZL  x
��Y�  w`��Y�      C  , ,  y���Y�  y���ZL  zX��ZL  zX��Y�  y���Y�      C  , ,  {���Y�  {���ZL  |���ZL  |���Y�  {���Y�      C  , ,  ~J��Y�  ~J��ZL  ~���ZL  ~���Y�  ~J��Y�      C  , ,  ����Y�  ����ZL  �B��ZL  �B��Y�  ����Y�      C  , ,  ����Y�  ����ZL  ����ZL  ����Y�  ����Y�      C  , ,  �4��Y�  �4��ZL  ����ZL  ����Y�  �4��Y�      C  , ,  ����Y�  ����ZL  �,��ZL  �,��Y�  ����Y�      C  , ,  ���`�  ���aT  ����aT  ����`�  ���`�      C  , ,  ���_B  ���_�  ����_�  ����_B  ���_B      C  , ,  ���]�  ���^�  ����^�  ����]�  ���]�      C  , ,  ���\r  ���]  ����]  ����\r  ���\r      C  , ,  ���h4  ���h�  ����h�  ����h4  ���h4      C  , ,  ���[
  ���[�  ����[�  ����[
  ���[
      C  , ,  �l��[
  �l��[�  ���[�  ���[
  �l��[
      C  , ,  ����[
  ����[�  �d��[�  �d��[
  ����[
      C  , ,  ���[
  ���[�  ����[�  ����[
  ���[
      C  , ,  �V��[
  �V��[�  � ��[�  � ��[
  �V��[
      C  , ,  ����[
  ����[�  �t��[�  �t��[
  ����[
      C  , ,  ���[
  ���[�  ����[�  ����[
  ���[
      C  , ,  �f��[
  �f��[�  ���[�  ���[
  �f��[
      C  , ,  ����[
  ����[�  �^��[�  �^��[
  ����[
      C  , ,  ���[
  ���[�  ����[�  ����[
  ���[
      C  , ,  �P��[
  �P��[�  ����[�  ����[
  �P��[
      C  , ,  ����[
  ����[�  �H��[�  �H��[
  ����[
      C  , ,  ����[
  ����[�  ����[�  ����[
  ����[
      C  , ,  �:��[
  �:��[�  ����[�  ����[
  �:��[
      C  , ,  ����[
  ����[�  �2��[�  �2��[
  ����[
      C  , ,  ����[
  ����[�  ����[�  ����[
  ����[
      C  , ,  �$��[
  �$��[�  ����[�  ����[
  �$��[
      C  , ,  �r��[
  �r��[�  ���[�  ���[
  �r��[
      C  , ,  ����[
  ����[�  �j��[�  �j��[
  ����[
      C  , ,  ���[
  ���[�  ����[�  ����[
  ���[
      C  , ,  ���b  ���b�  ����b�  ����b  ���b      C  , ,  ���Y�  ���ZL  ����ZL  ����Y�  ���Y�      C  , ,  ���X:  ���X�  ����X�  ����X:  ���X:      C  , ,  �$��_B  �$��_�  ����_�  ����_B  �$��_B      C  , ,  �r��_B  �r��_�  ���_�  ���_B  �r��_B      C  , ,  ����_B  ����_�  �j��_�  �j��_B  ����_B      C  , ,  ���_B  ���_�  ����_�  ����_B  ���_B      C  , ,  ����`�  ����aT  �H��aT  �H��`�  ����`�      C  , ,  �P��]�  �P��^�  ����^�  ����]�  �P��]�      C  , ,  ����]�  ����^�  �H��^�  �H��]�  ����]�      C  , ,  ����]�  ����^�  ����^�  ����]�  ����]�      C  , ,  �:��]�  �:��^�  ����^�  ����]�  �:��]�      C  , ,  ����]�  ����^�  �2��^�  �2��]�  ����]�      C  , ,  ����]�  ����^�  ����^�  ����]�  ����]�      C  , ,  �$��]�  �$��^�  ����^�  ����]�  �$��]�      C  , ,  �r��]�  �r��^�  ���^�  ���]�  �r��]�      C  , ,  ����]�  ����^�  �j��^�  �j��]�  ����]�      C  , ,  ���]�  ���^�  ����^�  ����]�  ���]�      C  , ,  �)��d  �)��d�  ����d�  ����d  �)��d      C  , ,  �w��d  �w��d�  �!��d�  �!��d  �w��d      C  , ,  ����d  ����d�  �o��d�  �o��d  ����d      C  , ,  ���d  ���d�  ����d�  ����d  ���d      C  , ,  �a��d  �a��d�  ���d�  ���d  �a��d      C  , ,  ����d  ����d�  �Y��d�  �Y��d  ����d      C  , ,  ����d  ����d�  ����d�  ����d  ����d      C  , ,  �K��d  �K��d�  ����d�  ����d  �K��d      C  , ,  ����d  ����d�  �C��d�  �C��d  ����d      C  , ,  ����d  ����d�  ����d�  ����d  ����d      C  , ,  ����`�  ����aT  ����aT  ����`�  ����`�      C  , ,  �P��\r  �P��]  ����]  ����\r  �P��\r      C  , ,  ����\r  ����]  �H��]  �H��\r  ����\r      C  , ,  ����\r  ����]  ����]  ����\r  ����\r      C  , ,  �:��\r  �:��]  ����]  ����\r  �:��\r      C  , ,  ����\r  ����]  �2��]  �2��\r  ����\r      C  , ,  ����\r  ����]  ����]  ����\r  ����\r      C  , ,  �$��\r  �$��]  ����]  ����\r  �$��\r      C  , ,  �r��\r  �r��]  ���]  ���\r  �r��\r      C  , ,  ����\r  ����]  �j��]  �j��\r  ����\r      C  , ,  ���\r  ���]  ����]  ����\r  ���\r      C  , ,  �5��d  �5��d�  ����d�  ����d  �5��d      C  , ,  �:��`�  �:��aT  ����aT  ����`�  �:��`�      C  , ,  �P��h4  �P��h�  ����h�  ����h4  �P��h4      C  , ,  ����h4  ����h�  �H��h�  �H��h4  ����h4      C  , ,  ����`�  ����aT  �2��aT  �2��`�  ����`�      C  , ,  ����`�  ����aT  ����aT  ����`�  ����`�      C  , ,  �$��`�  �$��aT  ����aT  ����`�  �$��`�      C  , ,  �r��`�  �r��aT  ���aT  ���`�  �r��`�      C  , ,  ����`�  ����aT  �j��aT  �j��`�  ����`�      C  , ,  ���`�  ���aT  ����aT  ����`�  ���`�      C  , ,  ����f1  ����f�  ����f�  ����f1  ����f1      C  , ,  �5��f1  �5��f�  ����f�  ����f1  �5��f1      C  , ,  ����h4  ����h�  ����h�  ����h4  ����h4      C  , ,  �:��h4  �:��h�  ����h�  ����h4  �:��h4      C  , ,  ����h4  ����h�  �2��h�  �2��h4  ����h4      C  , ,  ����h4  ����h�  ����h�  ����h4  ����h4      C  , ,  �$��h4  �$��h�  ����h�  ����h4  �$��h4      C  , ,  �r��h4  �r��h�  ���h�  ���h4  �r��h4      C  , ,  ����h4  ����h�  �j��h�  �j��h4  ����h4      C  , ,  ���h4  ���h�  ����h�  ����h4  ���h4      C  , ,  �P��`�  �P��aT  ����aT  ����`�  �P��`�      C  , ,  �P��_B  �P��_�  ����_�  ����_B  �P��_B      C  , ,  ����_B  ����_�  �H��_�  �H��_B  ����_B      C  , ,  ����_B  ����_�  ����_�  ����_B  ����_B      C  , ,  �:��_B  �:��_�  ����_�  ����_B  �:��_B      C  , ,  �P��b  �P��b�  ����b�  ����b  �P��b      C  , ,  ����_B  ����_�  �2��_�  �2��_B  ����_B      C  , ,  ����b  ����b�  �H��b�  �H��b  ����b      C  , ,  ����b  ����b�  ����b�  ����b  ����b      C  , ,  �:��b  �:��b�  ����b�  ����b  �:��b      C  , ,  ����b  ����b�  �2��b�  �2��b  ����b      C  , ,  ����b  ����b�  ����b�  ����b  ����b      C  , ,  �$��b  �$��b�  ����b�  ����b  �$��b      C  , ,  �r��b  �r��b�  ���b�  ���b  �r��b      C  , ,  ����b  ����b�  �j��b�  �j��b  ����b      C  , ,  ���b  ���b�  ����b�  ����b  ���b      C  , ,  ����_B  ����_�  ����_�  ����_B  ����_B      C  , ,  �)��f1  �)��f�  ����f�  ����f1  �)��f1      C  , ,  �w��f1  �w��f�  �!��f�  �!��f1  �w��f1      C  , ,  ����f1  ����f�  �o��f�  �o��f1  ����f1      C  , ,  ���f1  ���f�  ����f�  ����f1  ���f1      C  , ,  �a��f1  �a��f�  ���f�  ���f1  �a��f1      C  , ,  ����f1  ����f�  �Y��f�  �Y��f1  ����f1      C  , ,  ����f1  ����f�  ����f�  ����f1  ����f1      C  , ,  �K��f1  �K��f�  ����f�  ����f1  �K��f1      C  , ,  ����f1  ����f�  �C��f�  �C��f1  ����f1      C  , ,  ����d  ����d�  �7��d�  �7��d  ����d      C  , ,  ���]�  ���^�  ����^�  ����]�  ���]�      C  , ,  �l��]�  �l��^�  ���^�  ���]�  �l��]�      C  , ,  ����]�  ����^�  �d��^�  �d��]�  ����]�      C  , ,  ����h4  ����h�  �t��h�  �t��h4  ����h4      C  , ,  ���h4  ���h�  ����h�  ����h4  ���h4      C  , ,  �f��h4  �f��h�  ���h�  ���h4  �f��h4      C  , ,  ����h4  ����h�  �^��h�  �^��h4  ����h4      C  , ,  ���]�  ���^�  ����^�  ����]�  ���]�      C  , ,  �V��]�  �V��^�  � ��^�  � ��]�  �V��]�      C  , ,  ����]�  ����^�  �t��^�  �t��]�  ����]�      C  , ,  �E��f1  �E��f�  ����f�  ����f1  �E��f1      C  , ,  ����f1  ����f�  �=��f�  �=��f1  ����f1      C  , ,  ����f1  ����f�  ����f�  ����f1  ����f1      C  , ,  �/��f1  �/��f�  ����f�  ����f1  �/��f1      C  , ,  ���]�  ���^�  ����^�  ����]�  ���]�      C  , ,  �f��]�  �f��^�  ���^�  ���]�  �f��]�      C  , ,  ����]�  ����^�  �^��^�  �^��]�  ����]�      C  , ,  �l��_B  �l��_�  ���_�  ���_B  �l��_B      C  , ,  ����_B  ����_�  �d��_�  �d��_B  ����_B      C  , ,  ���_B  ���_�  ����_�  ����_B  ���_B      C  , ,  �V��_B  �V��_�  � ��_�  � ��_B  �V��_B      C  , ,  ����_B  ����_�  �t��_�  �t��_B  ����_B      C  , ,  ���_B  ���_�  ����_�  ����_B  ���_B      C  , ,  �f��_B  �f��_�  ���_�  ���_B  �f��_B      C  , ,  ����_B  ����_�  �^��_�  �^��_B  ����_B      C  , ,  ���`�  ���aT  ����aT  ����`�  ���`�      C  , ,  �V��`�  �V��aT  � ��aT  � ��`�  �V��`�      C  , ,  ����`�  ����aT  �t��aT  �t��`�  ����`�      C  , ,  ����d  ����d�  ����d�  ����d  ����d      C  , ,  ���`�  ���aT  ����aT  ����`�  ���`�      C  , ,  �f��`�  �f��aT  ���aT  ���`�  �f��`�      C  , ,  ����`�  ����aT  �^��aT  �^��`�  ����`�      C  , ,  ���`�  ���aT  ����aT  ����`�  ���`�      C  , ,  �l��`�  �l��aT  ���aT  ���`�  �l��`�      C  , ,  ����f1  ����f�  ����f�  ����f1  ����f1      C  , ,  ���b  ���b�  ����b�  ����b  ���b      C  , ,  �l��b  �l��b�  ���b�  ���b  �l��b      C  , ,  ����b  ����b�  �d��b�  �d��b  ����b      C  , ,  ���b  ���b�  ����b�  ����b  ���b      C  , ,  �V��b  �V��b�  � ��b�  � ��b  �V��b      C  , ,  ����b  ����b�  �t��b�  �t��b  ����b      C  , ,  ���b  ���b�  ����b�  ����b  ���b      C  , ,  �f��b  �f��b�  ���b�  ���b  �f��b      C  , ,  ����b  ����b�  �^��b�  �^��b  ����b      C  , ,  ����`�  ����aT  �d��aT  �d��`�  ����`�      C  , ,  ���h4  ���h�  ����h�  ����h4  ���h4      C  , ,  ���_B  ���_�  ����_�  ����_B  ���_B      C  , ,  �l��h4  �l��h�  ���h�  ���h4  �l��h4      C  , ,  ����h4  ����h�  �d��h�  �d��h4  ����h4      C  , ,  ���\r  ���]  ����]  ����\r  ���\r      C  , ,  �l��\r  �l��]  ���]  ���\r  �l��\r      C  , ,  ����\r  ����]  �d��]  �d��\r  ����\r      C  , ,  ���\r  ���]  ����]  ����\r  ���\r      C  , ,  �V��\r  �V��]  � ��]  � ��\r  �V��\r      C  , ,  ����\r  ����]  �t��]  �t��\r  ����\r      C  , ,  ���\r  ���]  ����]  ����\r  ���\r      C  , ,  �?��f1  �?��f�  ����f�  ����f1  �?��f1      C  , ,  ����f1  ����f�  �7��f�  �7��f1  ����f1      C  , ,  ����f1  ����f�  ����f�  ����f1  ����f1      C  , ,  �f��\r  �f��]  ���]  ���\r  �f��\r      C  , ,  ����\r  ����]  �^��]  �^��\r  ����\r      C  , ,  ���h4  ���h�  ����h�  ����h4  ���h4      C  , ,  �V��h4  �V��h�  � ��h�  � ��h4  �V��h4      C  , ,  �E��d  �E��d�  ����d�  ����d  �E��d      C  , ,  ����d  ����d�  �=��d�  �=��d  ����d      C  , ,  ����d  ����d�  ����d�  ����d  ����d      C  , ,  �/��d  �/��d�  ����d�  ����d  �/��d      C  , ,  ����d  ����d�  ����d�  ����d  ����d      C  , ,  �?��d  �?��d�  ����d�  ����d  �?��d      C  , ,  �l��X:  �l��X�  ���X�  ���X:  �l��X:      C  , ,  ����X:  ����X�  �d��X�  �d��X:  ����X:      C  , ,  ���X:  ���X�  ����X�  ����X:  ���X:      C  , ,  �V��X:  �V��X�  � ��X�  � ��X:  �V��X:      C  , ,  ����X:  ����X�  �t��X�  �t��X:  ����X:      C  , ,  ���X:  ���X�  ����X�  ����X:  ���X:      C  , ,  �f��X:  �f��X�  ���X�  ���X:  �f��X:      C  , ,  ����X:  ����X�  �^��X�  �^��X:  ����X:      C  , ,  �V��Y�  �V��ZL  � ��ZL  � ��Y�  �V��Y�      C  , ,  ����Y�  ����ZL  �t��ZL  �t��Y�  ����Y�      C  , ,  ���Y�  ���ZL  ����ZL  ����Y�  ���Y�      C  , ,  �f��Y�  �f��ZL  ���ZL  ���Y�  �f��Y�      C  , ,  ����Y�  ����ZL  �^��ZL  �^��Y�  ����Y�      C  , ,  ���Y�  ���ZL  ����ZL  ����Y�  ���Y�      C  , ,  �l��Y�  �l��ZL  ���ZL  ���Y�  �l��Y�      C  , ,  ����Y�  ����ZL  �d��ZL  �d��Y�  ����Y�      C  , ,  ���Y�  ���ZL  ����ZL  ����Y�  ���Y�      C  , ,  ���X:  ���X�  ����X�  ����X:  ���X:      C  , ,  ����Y�  ����ZL  �H��ZL  �H��Y�  ����Y�      C  , ,  �P��X:  �P��X�  ����X�  ����X:  �P��X:      C  , ,  ����X:  ����X�  �H��X�  �H��X:  ����X:      C  , ,  ����X:  ����X�  ����X�  ����X:  ����X:      C  , ,  �:��X:  �:��X�  ����X�  ����X:  �:��X:      C  , ,  ����X:  ����X�  �2��X�  �2��X:  ����X:      C  , ,  ����X:  ����X�  ����X�  ����X:  ����X:      C  , ,  �$��X:  �$��X�  ����X�  ����X:  �$��X:      C  , ,  �r��X:  �r��X�  ���X�  ���X:  �r��X:      C  , ,  ����X:  ����X�  �j��X�  �j��X:  ����X:      C  , ,  ���X:  ���X�  ����X�  ����X:  ���X:      C  , ,  ����Y�  ����ZL  ����ZL  ����Y�  ����Y�      C  , ,  �:��Y�  �:��ZL  ����ZL  ����Y�  �:��Y�      C  , ,  ����Y�  ����ZL  �2��ZL  �2��Y�  ����Y�      C  , ,  ����Y�  ����ZL  ����ZL  ����Y�  ����Y�      C  , ,  �$��Y�  �$��ZL  ����ZL  ����Y�  �$��Y�      C  , ,  �r��Y�  �r��ZL  ���ZL  ���Y�  �r��Y�      C  , ,  ����Y�  ����ZL  �j��ZL  �j��Y�  ����Y�      C  , ,  ���Y�  ���ZL  ����ZL  ����Y�  ���Y�      C  , ,  �P��Y�  �P��ZL  ����ZL  ����Y�  �P��Y�      C  , ,  �Z��h�  �Z��i�  ���i�  ���h�  �Z��h�      C  , ,  ����h�  ����i�  �l��i�  �l��h�  ����h�      C  , ,  �*��h�  �*��i�  ����i�  ����h�  �*��h�      C  , ,  ђ��h�  ђ��i�  �<��i�  �<��h�  ђ��h�      C  , ,  ����h�  ����i�  Ӥ��i�  Ӥ��h�  ����h�      C  , ,  �b��h�  �b��i�  ���i�  ���h�  �b��h�      C  , ,  ����h�  ����i�  �t��i�  �t��h�  ����h�      C  , ,  �2��h�  �2��i�  ����i�  ����h�  �2��h�      C  , ,  ؚ��h�  ؚ��i�  �D��i�  �D��h�  ؚ��h�      C  , ,  ���h�  ���i�  ڬ��i�  ڬ��h�  ���h�      C  , ,  �j��h�  �j��i�  ���i�  ���h�  �j��h�      C  , ,  ����i~  ����j(  �x��j(  �x��i~  ����i~      C  , ,  ����i~  ����j(  �\��j(  �\��i~  ����i~      C  , ,  ����i~  ����j(  �@��j(  �@��i~  ����i~      C  , ,  �z��i~  �z��j(  �$��j(  �$��i~  �z��i~      C  , ,  ^��i~  ^��j( ��j( ��i~  ^��i~      C  , , B��i~ B��j( ���j( ���i~ B��i~      C  , , &��i~ &��j( ���j( ���i~ &��i~      C  , , 	
��i~ 	
��j( 	���j( 	���i~ 	
��i~      C  , , ���i~ ���j( ���j( ���i~ ���i~      C  , , ���i~ ���j( |��j( |��i~ ���i~      C  , , ���i~ ���j( `��j( `��i~ ���i~      C  , , ���i~ ���j( D��j( D��i~ ���i~      C  , , ~��i~ ~��j( (��j( (��i~ ~��i~      C  , , b��i~ b��j( ��j( ��i~ b��i~      C  , , ���o ���o� |��o� |��o ���o      C  , , ���o ���o� `��o� `��o ���o      C  , , ���o ���o� D��o� D��o ���o      C  , , ~��o ~��o� (��o� (��o ~��o      C  , , b��o b��o� ��o� ��o b��o      C  , , ~��lN ~��l� (��l� (��lN ~��lN      C  , , b��lN b��l� ��l� ��lN b��lN      C  , ,  ����o  ����o�  �x��o�  �x��o  ����o      C  , ,  ����o  ����o�  �\��o�  �\��o  ����o      C  , ,  ����o  ����o�  �@��o�  �@��o  ����o      C  , ,  �z��o  �z��o�  �$��o�  �$��o  �z��o      C  , ,  ^��o  ^��o� ��o� ��o  ^��o      C  , , B��o B��o� ���o� ���o B��o      C  , ,  ����j�  ����k�  �x��k�  �x��j�  ����j�      C  , ,  ����j�  ����k�  �\��k�  �\��j�  ����j�      C  , ,  ����j�  ����k�  �@��k�  �@��j�  ����j�      C  , ,  �z��j�  �z��k�  �$��k�  �$��j�  �z��j�      C  , ,  ^��j�  ^��k� ��k� ��j�  ^��j�      C  , , B��j� B��k� ���k� ���j� B��j�      C  , , &��j� &��k� ���k� ���j� &��j�      C  , , 	
��j� 	
��k� 	���k� 	���j� 	
��j�      C  , , ���j� ���k� ���k� ���j� ���j�      C  , , ���j� ���k� |��k� |��j� ���j�      C  , , ���j� ���k� `��k� `��j� ���j�      C  , , ���j� ���k� D��k� D��j� ���j�      C  , , ~��j� ~��k� (��k� (��j� ~��j�      C  , , b��j� b��k� ��k� ��j� b��j�      C  , , &��o &��o� ���o� ���o &��o      C  , , 	
��o 	
��o� 	���o� 	���o 	
��o      C  , , ���o ���o� ���o� ���o ���o      C  , ,  ����p�  ����q0  �x��q0  �x��p�  ����p�      C  , ,  ����p�  ����q0  �\��q0  �\��p�  ����p�      C  , ,  ����m�  ����n`  �x��n`  �x��m�  ����m�      C  , ,  ����m�  ����n`  �\��n`  �\��m�  ����m�      C  , ,  ����m�  ����n`  �@��n`  �@��m�  ����m�      C  , ,  �z��m�  �z��n`  �$��n`  �$��m�  �z��m�      C  , ,  ^��m�  ^��n` ��n` ��m�  ^��m�      C  , , B��m� B��n` ���n` ���m� B��m�      C  , , &��m� &��n` ���n` ���m� &��m�      C  , , 	
��m� 	
��n` 	���n` 	���m� 	
��m�      C  , , ���m� ���n` ���n` ���m� ���m�      C  , , ���m� ���n` |��n` |��m� ���m�      C  , , ���m� ���n` `��n` `��m� ���m�      C  , , ���m� ���n` D��n` D��m� ���m�      C  , , ~��m� ~��n` (��n` (��m� ~��m�      C  , , b��m� b��n` ��n` ��m� b��m�      C  , ,  ����p�  ����q0  �@��q0  �@��p�  ����p�      C  , ,  �z��p�  �z��q0  �$��q0  �$��p�  �z��p�      C  , ,  ^��p�  ^��q0 ��q0 ��p�  ^��p�      C  , , B��p� B��q0 ���q0 ���p� B��p�      C  , , &��p� &��q0 ���q0 ���p� &��p�      C  , , 	
��p� 	
��q0 	���q0 	���p� 	
��p�      C  , , ���p� ���q0 ���q0 ���p� ���p�      C  , , ���p� ���q0 |��q0 |��p� ���p�      C  , , ���p� ���q0 `��q0 `��p� ���p�      C  , , ���p� ���q0 D��q0 D��p� ���p�      C  , , ~��p� ~��q0 (��q0 (��p� ~��p�      C  , , b��p� b��q0 ��q0 ��p� b��p�      C  , ,  ����q�  ����r�  �x��r�  �x��q�  ����q�      C  , ,  ����q�  ����r�  �\��r�  �\��q�  ����q�      C  , ,  ����q�  ����r�  �@��r�  �@��q�  ����q�      C  , ,  �z��q�  �z��r�  �$��r�  �$��q�  �z��q�      C  , ,  ^��q�  ^��r� ��r� ��q�  ^��q�      C  , , B��q� B��r� ���r� ���q� B��q�      C  , , &��q� &��r� ���r� ���q� &��q�      C  , , 	
��q� 	
��r� 	���r� 	���q� 	
��q�      C  , , ���q� ���r� ���r� ���q� ���q�      C  , , ���q� ���r� |��r� |��q� ���q�      C  , , ���q� ���r� `��r� `��q� ���q�      C  , , ���q� ���r� D��r� D��q� ���q�      C  , , ~��q� ~��r� (��r� (��q� ~��q�      C  , , b��q� b��r� ��r� ��q� b��q�      C  , ,  ����lN  ����l�  �x��l�  �x��lN  ����lN      C  , ,  ����lN  ����l�  �\��l�  �\��lN  ����lN      C  , ,  ����lN  ����l�  �@��l�  �@��lN  ����lN      C  , ,  �z��lN  �z��l�  �$��l�  �$��lN  �z��lN      C  , ,  ^��lN  ^��l� ��l� ��lN  ^��lN      C  , , B��lN B��l� ���l� ���lN B��lN      C  , , &��lN &��l� ���l� ���lN &��lN      C  , , 	
��lN 	
��l� 	���l� 	���lN 	
��lN      C  , , ���lN ���l� ���l� ���lN ���lN      C  , , ���lN ���l� |��l� |��lN ���lN      C  , , ���lN ���l� `��l� `��lN ���lN      C  , , ���lN ���l� D��l� D��lN ���lN      C  , ,  �\��o<  �\��o�  ���o�  ���o<  �\��o<      C  , ,  �Z��n�  �Z��od  ���od  ���n�  �Z��n�      C  , ,  ����n�  ����od  �l��od  �l��n�  ����n�      C  , ,  �*��n�  �*��od  ����od  ����n�  �*��n�      C  , ,  ђ��n�  ђ��od  �<��od  �<��n�  ђ��n�      C  , ,  �b��p,  �b��p�  ���p�  ���p,  �b��p,      C  , ,  ����p,  ����p�  �t��p�  �t��p,  ����p,      C  , ,  �2��p,  �2��p�  ����p�  ����p,  �2��p,      C  , ,  ؚ��p,  ؚ��p�  �D��p�  �D��p,  ؚ��p,      C  , ,  ���p,  ���p�  ڬ��p�  ڬ��p,  ���p,      C  , ,  �j��p,  �j��p�  ���p�  ���p,  �j��p,      C  , ,  ����n�  ����od  Ӥ��od  Ӥ��n�  ����n�      C  , ,  �b��n�  �b��od  ���od  ���n�  �b��n�      C  , ,  �\��m�  �\��n~  ���n~  ���m�  �\��m�      C  , ,  �Z��mH  �Z��m�  ���m�  ���mH  �Z��mH      C  , ,  ����mH  ����m�  �l��m�  �l��mH  ����mH      C  , ,  �*��mH  �*��m�  ����m�  ����mH  �*��mH      C  , ,  ђ��mH  ђ��m�  �<��m�  �<��mH  ђ��mH      C  , ,  ����mH  ����m�  Ӥ��m�  Ӥ��mH  ����mH      C  , ,  �b��mH  �b��m�  ���m�  ���mH  �b��mH      C  , ,  ����mH  ����m�  �t��m�  �t��mH  ����mH      C  , ,  �2��mH  �2��m�  ����m�  ����mH  �2��mH      C  , ,  ؚ��mH  ؚ��m�  �D��m�  �D��mH  ؚ��mH      C  , ,  ���mH  ���m�  ڬ��m�  ڬ��mH  ���mH      C  , ,  �j��mH  �j��m�  ���m�  ���mH  �j��mH      C  , ,  ����n�  ����od  �t��od  �t��n�  ����n�      C  , ,  �2��n�  �2��od  ����od  ����n�  �2��n�      C  , ,  ؚ��n�  ؚ��od  �D��od  �D��n�  ؚ��n�      C  , ,  ���n�  ���od  ڬ��od  ڬ��n�  ���n�      C  , ,  �j��n�  �j��od  ���od  ���n�  �j��n�      C  , ,  ������  �����Y  �h���Y  �h����  ������      C  , ,  �����  ����Y  �����Y  ������  �����      C  , ,  �Z����  �Z���Y  ����Y  �����  �Z����      C  , ,  Ũ����  Ũ���Y  �R���Y  �R����  Ũ����      C  , ,  Ũ���  Ũ����  �R����  �R���  Ũ���      C  , ,  �����  ������  Ƞ����  Ƞ���  �����      C  , ,  �D���  �D����  ������  �����  �D���      C  , ,  ̒���  ̒����  �<����  �<���  ̒���      C  , ,  �����  ������  ϊ����  ϊ���  �����      C  , ,  �.���  �.����  ������  �����  �.���      C  , ,  �\��r  �\��r�  ���r�  ���r  �\��r      C  , ,  �Z��q�  �Z��rH  ���rH  ���q�  �Z��q�      C  , ,  ����q�  ����rH  �l��rH  �l��q�  ����q�      C  , ,  �*��q�  �*��rH  ����rH  ����q�  �*��q�      C  , ,  ђ��q�  ђ��rH  �<��rH  �<��q�  ђ��q�      C  , ,  ����q�  ����rH  Ӥ��rH  Ӥ��q�  ����q�      C  , ,  �b��q�  �b��rH  ���rH  ���q�  �b��q�      C  , ,  ����q�  ����rH  �t��rH  �t��q�  ����q�      C  , ,  �2��q�  �2��rH  ����rH  ����q�  �2��q�      C  , ,  ؚ��q�  ؚ��rH  �D��rH  �D��q�  ؚ��q�      C  , ,  �\��p�  �\��qN  ���qN  ���p�  �\��p�      C  , ,  ���q�  ���rH  ڬ��rH  ڬ��q�  ���q�      C  , ,  �j��q�  �j��rH  ���rH  ���q�  �j��q�      C  , ,  �Z��p,  �Z��p�  ���p�  ���p,  �Z��p,      C  , ,  ����p,  ����p�  �l��p�  �l��p,  ����p,      C  , ,  �*��p,  �*��p�  ����p�  ����p,  �*��p,      C  , ,  ђ��p,  ђ��p�  �<��p�  �<��p,  ђ��p,      C  , ,  ����p,  ����p�  Ӥ��p�  Ӥ��p,  ����p,      C  , ,  �\��i�  �\��jF  ���jF  ���i�  �\��i�      C  , ,  ������  �����Y  Ƞ���Y  Ƞ����  ������      C  , ,  �D����  �D���Y  �����Y  ������  �D����      C  , ,  �\��k  �\��k�  ���k�  ���k  �\��k      C  , ,  �Z��jd  �Z��k  ���k  ���jd  �Z��jd      C  , ,  ����jd  ����k  �l��k  �l��jd  ����jd      C  , ,  �*��jd  �*��k  ����k  ����jd  �*��jd      C  , ,  ђ��jd  ђ��k  �<��k  �<��jd  ђ��jd      C  , ,  ����jd  ����k  Ӥ��k  Ӥ��jd  ����jd      C  , ,  �p���  �p����  �����  ����  �p���      C  , ,  �p����  �p���Y  ����Y  �����  �p����      C  , ,  �\��ll  �\��m  ���m  ���ll  �\��ll      C  , ,  �Z��k�  �Z��l�  ���l�  ���k�  �Z��k�      C  , ,  ����k�  ����l�  �l��l�  �l��k�  ����k�      C  , ,  �*��k�  �*��l�  ����l�  ����k�  �*��k�      C  , ,  ђ��k�  ђ��l�  �<��l�  �<��k�  ђ��k�      C  , ,  ����k�  ����l�  Ӥ��l�  Ӥ��k�  ����k�      C  , ,  �b��k�  �b��l�  ���l�  ���k�  �b��k�      C  , ,  ����k�  ����l�  �t��l�  �t��k�  ����k�      C  , ,  �2��k�  �2��l�  ����l�  ����k�  �2��k�      C  , ,  ؚ��k�  ؚ��l�  �D��l�  �D��k�  ؚ��k�      C  , ,  ���k�  ���l�  ڬ��l�  ڬ��k�  ���k�      C  , ,  �j��k�  �j��l�  ���l�  ���k�  �j��k�      C  , ,  �b��jd  �b��k  ���k  ���jd  �b��jd      C  , ,  ����jd  ����k  �t��k  �t��jd  ����jd      C  , ,  �2��jd  �2��k  ����k  ����jd  �2��jd      C  , ,  ؚ��jd  ؚ��k  �D��k  �D��jd  ؚ��jd      C  , ,  ���jd  ���k  ڬ��k  ڬ��jd  ���jd      C  , ,  �j��jd  �j��k  ���k  ���jd  �j��jd      C  , ,  ̒����  ̒���Y  �<���Y  �<����  ̒����      C  , ,  ������  �����Y  ϊ���Y  ϊ����  ������      C  , ,  �.����  �.���Y  �����Y  ������  �.����      C  , ,  �����  ������  �h����  �h���  �����      C  , ,  ����  �����  ������  �����  ����      C  , ,  �Z���  �Z����  �����  ����  �Z���      C  , ,  �b��d�  �b��eF  ���eF  ���d�  �b��d�      C  , ,  �b��g�  �b��h*  ���h*  ���g�  �b��g�      C  , ,  �b��[�  �b��\�  ���\�  ���[�  �b��[�      C  , ,  �b��^�  �b��_~  ���_~  ���^�  �b��^�      C  , ,  �b��a�  �b��bb  ���bb  ���a�  �b��a�      C  , ,  �b��`F  �b��`�  ���`�  ���`F  �b��`F      C  , ,  �\��[
  �\��[�  ���[�  ���[
  �\��[
      C  , ,  �Z��Z~  �Z��[(  ���[(  ���Z~  �Z��Z~      C  , ,  ����Z~  ����[(  �l��[(  �l��Z~  ����Z~      C  , ,  �*��Z~  �*��[(  ����[(  ����Z~  �*��Z~      C  , ,  ђ��Z~  ђ��[(  �<��[(  �<��Z~  ђ��Z~      C  , ,  ����Z~  ����[(  Ӥ��[(  Ӥ��Z~  ����Z~      C  , ,  �b��Z~  �b��[(  ���[(  ���Z~  �b��Z~      C  , ,  ����Z~  ����[(  �t��[(  �t��Z~  ����Z~      C  , ,  �2��Z~  �2��[(  ����[(  ����Z~  �2��Z~      C  , ,  ؚ��Z~  ؚ��[(  �D��[(  �D��Z~  ؚ��Z~      C  , ,  ���Z~  ���[(  ڬ��[(  ڬ��Z~  ���Z~      C  , ,  �j��Z~  �j��[(  ���[(  ���Z~  �j��Z~      C  , ,  �b��f  �b��f�  ���f�  ���f  �b��f      C  , ,  �b��Y  �b��Y�  ���Y�  ���Y  �b��Y      C  , ,  �b��c*  �b��c�  ���c�  ���c*  �b��c*      C  , ,  �b��W�  �b��XD  ���XD  ���W�  �b��W�      C  , ,  �b��V(  �b��V�  ���V�  ���V(  �b��V(      C  , ,  �b��]b  �b��^  ���^  ���]b  �b��]b      C  , ,  ���d�  ���eF  ڬ��eF  ڬ��d�  ���d�      C  , ,  ����a�  ����bb  �t��bb  �t��a�  ����a�      C  , ,  �2��a�  �2��bb  ����bb  ����a�  �2��a�      C  , ,  �j��d�  �j��eF  ���eF  ���d�  �j��d�      C  , ,  ����d�  ����eF  �t��eF  �t��d�  ����d�      C  , ,  ����g�  ����h*  �t��h*  �t��g�  ����g�      C  , ,  �2��g�  �2��h*  ����h*  ����g�  �2��g�      C  , ,  ؚ��g�  ؚ��h*  �D��h*  �D��g�  ؚ��g�      C  , ,  ���g�  ���h*  ڬ��h*  ڬ��g�  ���g�      C  , ,  �j��g�  �j��h*  ���h*  ���g�  �j��g�      C  , ,  �2��d�  �2��eF  ����eF  ����d�  �2��d�      C  , ,  ����[�  ����\�  �t��\�  �t��[�  ����[�      C  , ,  �2��[�  �2��\�  ����\�  ����[�  �2��[�      C  , ,  ؚ��[�  ؚ��\�  �D��\�  �D��[�  ؚ��[�      C  , ,  ���[�  ���\�  ڬ��\�  ڬ��[�  ���[�      C  , ,  �j��[�  �j��\�  ���\�  ���[�  �j��[�      C  , ,  ����`F  ����`�  �t��`�  �t��`F  ����`F      C  , ,  �2��`F  �2��`�  ����`�  ����`F  �2��`F      C  , ,  ؚ��`F  ؚ��`�  �D��`�  �D��`F  ؚ��`F      C  , ,  ���`F  ���`�  ڬ��`�  ڬ��`F  ���`F      C  , ,  �j��`F  �j��`�  ���`�  ���`F  �j��`F      C  , ,  ؚ��a�  ؚ��bb  �D��bb  �D��a�  ؚ��a�      C  , ,  ���a�  ���bb  ڬ��bb  ڬ��a�  ���a�      C  , ,  ؚ��d�  ؚ��eF  �D��eF  �D��d�  ؚ��d�      C  , ,  ����f  ����f�  �t��f�  �t��f  ����f      C  , ,  �2��f  �2��f�  ����f�  ����f  �2��f      C  , ,  ؚ��f  ؚ��f�  �D��f�  �D��f  ؚ��f      C  , ,  ���f  ���f�  ڬ��f�  ڬ��f  ���f      C  , ,  �j��f  �j��f�  ���f�  ���f  �j��f      C  , ,  ����^�  ����_~  �t��_~  �t��^�  ����^�      C  , ,  �j��a�  �j��bb  ���bb  ���a�  �j��a�      C  , ,  �2��^�  �2��_~  ����_~  ����^�  �2��^�      C  , ,  ����c*  ����c�  �t��c�  �t��c*  ����c*      C  , ,  �2��c*  �2��c�  ����c�  ����c*  �2��c*      C  , ,  ؚ��c*  ؚ��c�  �D��c�  �D��c*  ؚ��c*      C  , ,  ���c*  ���c�  ڬ��c�  ڬ��c*  ���c*      C  , ,  �j��c*  �j��c�  ���c�  ���c*  �j��c*      C  , ,  ؚ��^�  ؚ��_~  �D��_~  �D��^�  ؚ��^�      C  , ,  ���^�  ���_~  ڬ��_~  ڬ��^�  ���^�      C  , ,  �j��^�  �j��_~  ���_~  ���^�  �j��^�      C  , ,  ����]b  ����^  �t��^  �t��]b  ����]b      C  , ,  �2��]b  �2��^  ����^  ����]b  �2��]b      C  , ,  ؚ��]b  ؚ��^  �D��^  �D��]b  ؚ��]b      C  , ,  ���]b  ���^  ڬ��^  ڬ��]b  ���]b      C  , ,  �j��]b  �j��^  ���^  ���]b  �j��]b      C  , ,  ����a�  ����bb  Ӥ��bb  Ӥ��a�  ����a�      C  , ,  �\��_B  �\��_�  ���_�  ���_B  �\��_B      C  , ,  �Z��^�  �Z��_~  ���_~  ���^�  �Z��^�      C  , ,  ����^�  ����_~  �l��_~  �l��^�  ����^�      C  , ,  �*��^�  �*��_~  ����_~  ����^�  �*��^�      C  , ,  ђ��^�  ђ��_~  �<��_~  �<��^�  ђ��^�      C  , ,  ����^�  ����_~  Ӥ��_~  Ӥ��^�  ����^�      C  , ,  ђ��d�  ђ��eF  �<��eF  �<��d�  ђ��d�      C  , ,  �\��b  �\��b�  ���b�  ���b  �\��b      C  , ,  ����d�  ����eF  Ӥ��eF  Ӥ��d�  ����d�      C  , ,  �Z��f  �Z��f�  ���f�  ���f  �Z��f      C  , ,  ����f  ����f�  �l��f�  �l��f  ����f      C  , ,  �*��f  �*��f�  ����f�  ����f  �*��f      C  , ,  ђ��f  ђ��f�  �<��f�  �<��f  ђ��f      C  , ,  ����f  ����f�  Ӥ��f�  Ӥ��f  ����f      C  , ,  �Z��a�  �Z��bb  ���bb  ���a�  �Z��a�      C  , ,  ����a�  ����bb  �l��bb  �l��a�  ����a�      C  , ,  �*��a�  �*��bb  ����bb  ����a�  �*��a�      C  , ,  �\��\r  �\��]  ���]  ���\r  �\��\r      C  , ,  �Z��[�  �Z��\�  ���\�  ���[�  �Z��[�      C  , ,  ����[�  ����\�  �l��\�  �l��[�  ����[�      C  , ,  �\��`�  �\��aT  ���aT  ���`�  �\��`�      C  , ,  �Z��`F  �Z��`�  ���`�  ���`F  �Z��`F      C  , ,  �Z��d�  �Z��eF  ���eF  ���d�  �Z��d�      C  , ,  �Z��c*  �Z��c�  ���c�  ���c*  �Z��c*      C  , ,  ����c*  ����c�  �l��c�  �l��c*  ����c*      C  , ,  �*��c*  �*��c�  ����c�  ����c*  �*��c*      C  , ,  ђ��c*  ђ��c�  �<��c�  �<��c*  ђ��c*      C  , ,  ����c*  ����c�  Ӥ��c�  Ӥ��c*  ����c*      C  , ,  ����`F  ����`�  �l��`�  �l��`F  ����`F      C  , ,  �*��`F  �*��`�  ����`�  ����`F  �*��`F      C  , ,  ђ��`F  ђ��`�  �<��`�  �<��`F  ђ��`F      C  , ,  ����`F  ����`�  Ӥ��`�  Ӥ��`F  ����`F      C  , ,  �*��[�  �*��\�  ����\�  ����[�  �*��[�      C  , ,  ђ��[�  ђ��\�  �<��\�  �<��[�  ђ��[�      C  , ,  ����d�  ����eF  �l��eF  �l��d�  ����d�      C  , ,  �\��]�  �\��^�  ���^�  ���]�  �\��]�      C  , ,  �Z��]b  �Z��^  ���^  ���]b  �Z��]b      C  , ,  ����]b  ����^  �l��^  �l��]b  ����]b      C  , ,  �*��]b  �*��^  ����^  ����]b  �*��]b      C  , ,  ����[�  ����\�  Ӥ��\�  Ӥ��[�  ����[�      C  , ,  ђ��]b  ђ��^  �<��^  �<��]b  ђ��]b      C  , ,  �\��h4  �\��h�  ���h�  ���h4  �\��h4      C  , ,  ����]b  ����^  Ӥ��^  Ӥ��]b  ����]b      C  , ,  �Z��g�  �Z��h*  ���h*  ���g�  �Z��g�      C  , ,  ����g�  ����h*  �l��h*  �l��g�  ����g�      C  , ,  �*��g�  �*��h*  ����h*  ����g�  �*��g�      C  , ,  ђ��g�  ђ��h*  �<��h*  �<��g�  ђ��g�      C  , ,  ����g�  ����h*  Ӥ��h*  Ӥ��g�  ����g�      C  , ,  ђ��a�  ђ��bb  �<��bb  �<��a�  ђ��a�      C  , ,  �*��d�  �*��eF  ����eF  ����d�  �*��d�      C  , ,  ����W�  ����XD  Ӥ��XD  Ӥ��W�  ����W�      C  , ,  �Z��Y  �Z��Y�  ���Y�  ���Y  �Z��Y      C  , ,  ����Y  ����Y�  �l��Y�  �l��Y  ����Y      C  , ,  �Z��V(  �Z��V�  ���V�  ���V(  �Z��V(      C  , ,  ����V(  ����V�  �l��V�  �l��V(  ����V(      C  , ,  �*��V(  �*��V�  ����V�  ����V(  �*��V(      C  , ,  ђ��V(  ђ��V�  �<��V�  �<��V(  ђ��V(      C  , ,  ����V(  ����V�  Ӥ��V�  Ӥ��V(  ����V(      C  , ,  �*��Y  �*��Y�  ����Y�  ����Y  �*��Y      C  , ,  ђ��Y  ђ��Y�  �<��Y�  �<��Y  ђ��Y      C  , ,  ����Y  ����Y�  Ӥ��Y�  Ӥ��Y  ����Y      C  , ,  �\��Y�  �\��ZL  ���ZL  ���Y�  �\��Y�      C  , ,  �\��X:  �\��X�  ���X�  ���X:  �\��X:      C  , ,  �Z��W�  �Z��XD  ���XD  ���W�  �Z��W�      C  , ,  ����W�  ����XD  �l��XD  �l��W�  ����W�      C  , ,  �*��W�  �*��XD  ����XD  ����W�  �*��W�      C  , ,  ђ��W�  ђ��XD  �<��XD  �<��W�  ђ��W�      C  , ,  ����W�  ����XD  �t��XD  �t��W�  ����W�      C  , ,  �2��W�  �2��XD  ����XD  ����W�  �2��W�      C  , ,  ����V(  ����V�  �t��V�  �t��V(  ����V(      C  , ,  �2��V(  �2��V�  ����V�  ����V(  �2��V(      C  , ,  ؚ��V(  ؚ��V�  �D��V�  �D��V(  ؚ��V(      C  , ,  ���V(  ���V�  ڬ��V�  ڬ��V(  ���V(      C  , ,  �j��V(  �j��V�  ���V�  ���V(  �j��V(      C  , ,  ؚ��W�  ؚ��XD  �D��XD  �D��W�  ؚ��W�      C  , ,  ���W�  ���XD  ڬ��XD  ڬ��W�  ���W�      C  , ,  �j��W�  �j��XD  ���XD  ���W�  �j��W�      C  , ,  ����Y  ����Y�  �t��Y�  �t��Y  ����Y      C  , ,  �2��Y  �2��Y�  ����Y�  ����Y  �2��Y      C  , ,  ؚ��Y  ؚ��Y�  �D��Y�  �D��Y  ؚ��Y      C  , ,  ���Y  ���Y�  ڬ��Y�  ڬ��Y  ���Y      C  , ,  �j��Y  �j��Y�  ���Y�  ���Y  �j��Y      C  , ,  ����Z�  ����[Z  �x��[Z  �x��Z�  ����Z�      C  , ,  ����Z�  ����[Z  �\��[Z  �\��Z�  ����Z�      C  , ,  ����Z�  ����[Z  �@��[Z  �@��Z�  ����Z�      C  , ,  �z��Z�  �z��[Z  �$��[Z  �$��Z�  �z��Z�      C  , ,  ^��Z�  ^��[Z ��[Z ��Z�  ^��Z�      C  , , B��Z� B��[Z ���[Z ���Z� B��Z�      C  , , &��Z� &��[Z ���[Z ���Z� &��Z�      C  , , 	
��Z� 	
��[Z 	���[Z 	���Z� 	
��Z�      C  , , ���Z� ���[Z ���[Z ���Z� ���Z�      C  , , ���Z� ���[Z |��[Z |��Z� ���Z�      C  , , ���Z� ���[Z `��[Z `��Z� ���Z�      C  , , ���Z� ���[Z D��[Z D��Z� ���Z�      C  , , ~��Z� ~��[Z (��[Z (��Z� ~��Z�      C  , , b��Z� b��[Z ��[Z ��Z� b��Z�      C  , , &��bv &��c  ���c  ���bv &��bv      C  , , 	
��bv 	
��c  	���c  	���bv 	
��bv      C  , , ���bv ���c  ���c  ���bv ���bv      C  , , ���bv ���c  |��c  |��bv ���bv      C  , , ���bv ���c  `��c  `��bv ���bv      C  , , ���bv ���c  D��c  D��bv ���bv      C  , , ~��bv ~��c  (��c  (��bv ~��bv      C  , , ���`U ���`� B��`� B��`U ���`U      C  , , &��f� &��gX ���gX ���f� &��f�      C  , , 	
��f� 	
��gX 	���gX 	���f� 	
��f�      C  , , ���f� ���gX ���gX ���f� ���f�      C  , , ���f� ���gX |��gX |��f� ���f�      C  , , ���f� ���gX `��gX `��f� ���f�      C  , , ���f� ���gX D��gX D��f� ���f�      C  , , ~��f� ~��gX (��gX (��f� ~��f�      C  , , b��f� b��gX ��gX ��f� b��f�      C  , , ���^9 ���^� B��^� B��^9 ���^9      C  , , 
|��^9 
|��^� &��^� &��^9 
|��^9      C  , , &��\ &��\� ���\� ���\ &��\      C  , , &��eF &��e� ���e� ���eF &��eF      C  , , 	
��eF 	
��e� 	���e� 	���eF 	
��eF      C  , , ���eF ���e� ���e� ���eF ���eF      C  , , ���eF ���e� |��e� |��eF ���eF      C  , , ���eF ���e� `��e� `��eF ���eF      C  , , ���eF ���e� D��e� D��eF ���eF      C  , , ~��eF ~��e� (��e� (��eF ~��eF      C  , , b��eF b��e� ��e� ��eF b��eF      C  , , 	
��\ 	
��\� 	���\� 	���\ 	
��\      C  , , ���\ ���\� ���\� ���\ ���\      C  , , ���\ ���\� |��\� |��\ ���\      C  , , ���\ ���\� `��\� `��\ ���\      C  , , ���\ ���\� D��\� D��\ ���\      C  , , ~��\ ~��\� (��\� (��\ ~��\      C  , , b��\ b��\� ��\� ��\ b��\      C  , , &��h &��h� ���h� ���h &��h      C  , , 	
��h 	
��h� 	���h� 	���h 	
��h      C  , , ���h ���h� ���h� ���h ���h      C  , , ���h ���h� |��h� |��h ���h      C  , , ���h ���h� `��h� `��h ���h      C  , , ���h ���h� D��h� D��h ���h      C  , , ~��h ~��h� (��h� (��h ~��h      C  , , b��h b��h� ��h� ��h b��h      C  , , `��^9 `��^� 
��^� 
��^9 `��^9      C  , , D��^9 D��^� ���^� ���^9 D��^9      C  , , (��^9 (��^� ���^� ���^9 (��^9      C  , , ��^9 ��^� ���^� ���^9 ��^9      C  , , ���^9 ���^� ���^� ���^9 ���^9      C  , , ���^9 ���^� ~��^� ~��^9 ���^9      C  , , 
|��`U 
|��`� &��`� &��`U 
|��`U      C  , , `��`U `��`� 
��`� 
��`U `��`U      C  , , D��`U D��`� ���`� ���`U D��`U      C  , , (��`U (��`� ���`� ���`U (��`U      C  , , ��`U ��`� ���`� ���`U ��`U      C  , , ���`U ���`� ���`� ���`U ���`U      C  , , ���`U ���`� ~��`� ~��`U ���`U      C  , , b��bv b��c  ��c  ��bv b��bv      C  , , &��c� &��d� ���d� ���c� &��c�      C  , , 	
��c� 	
��d� 	���d� 	���c� 	
��c�      C  , , ���c� ���d� ���d� ���c� ���c�      C  , , ���c� ���d� |��d� |��c� ���c�      C  , , ���c� ���d� `��d� `��c� ���c�      C  , , ���c� ���d� D��d� D��c� ���c�      C  , , ~��c� ~��d� (��d� (��c� ~��c�      C  , , b��c� b��d� ��d� ��c� b��c�      C  , ,  ^��h  ^��h� ��h� ��h  ^��h      C  , , B��h B��h� ���h� ���h B��h      C  , ,  ���`U  ���`�  ����`�  ����`U  ���`U      C  , ,  ����`U  ����`�  ����`�  ����`U  ����`U      C  , ,  ���^9  ���^�  ����^�  ����^9  ���^9      C  , ,  ����^9  ����^�  ����^�  ����^9  ����^9      C  , , ���^9 ���^� z��^� z��^9 ���^9      C  , , ���^9 ���^� ^��^� ^��^9 ���^9      C  , , ���`U ���`� z��`� z��`U ���`U      C  , , ���`U ���`� ^��`� ^��`U ���`U      C  , ,  ����\  ����\�  �x��\�  �x��\  ����\      C  , ,  ����\  ����\�  �\��\�  �\��\  ����\      C  , ,  ����\  ����\�  �@��\�  �@��\  ����\      C  , ,  �z��\  �z��\�  �$��\�  �$��\  �z��\      C  , ,  ^��\  ^��\� ��\� ��\  ^��\      C  , , B��\ B��\� ���\� ���\ B��\      C  , ,  �$��`U  �$��`�  ����`�  ����`U  �$��`U      C  , ,  ����eF  ����e�  �x��e�  �x��eF  ����eF      C  , ,  ����eF  ����e�  �\��e�  �\��eF  ����eF      C  , ,  ����eF  ����e�  �@��e�  �@��eF  ����eF      C  , ,  �z��eF  �z��e�  �$��e�  �$��eF  �z��eF      C  , ,  ^��eF  ^��e� ��e� ��eF  ^��eF      C  , , B��eF B��e� ���e� ���eF B��eF      C  , ,  �$��^9  �$��^�  ����^�  ����^9  �$��^9      C  , ,  ����f�  ����gX  �x��gX  �x��f�  ����f�      C  , ,  ����f�  ����gX  �\��gX  �\��f�  ����f�      C  , ,  ����c�  ����d�  �@��d�  �@��c�  ����c�      C  , ,  �z��c�  �z��d�  �$��d�  �$��c�  �z��c�      C  , ,  ^��c�  ^��d� ��d� ��c�  ^��c�      C  , , B��c� B��d� ���d� ���c� B��c�      C  , ,  ����f�  ����gX  �@��gX  �@��f�  ����f�      C  , ,  �z��f�  �z��gX  �$��gX  �$��f�  �z��f�      C  , ,  ^��f�  ^��gX ��gX ��f�  ^��f�      C  , , B��f� B��gX ���gX ���f� B��f�      C  , ,  ����h  ����h�  �x��h�  �x��h  ����h      C  , ,  ����h  ����h�  �\��h�  �\��h  ����h      C  , ,  ����h  ����h�  �@��h�  �@��h  ����h      C  , ,  �z��h  �z��h�  �$��h�  �$��h  �z��h      C  , ,  ����c�  ����d�  �x��d�  �x��c�  ����c�      C  , ,  ����c�  ����d�  �\��d�  �\��c�  ����c�      C  , ,  ����bv  ����c   �x��c   �x��bv  ����bv      C  , ,  ����bv  ����c   �\��c   �\��bv  ����bv      C  , ,  ����bv  ����c   �@��c   �@��bv  ����bv      C  , ,  �z��bv  �z��c   �$��c   �$��bv  �z��bv      C  , ,  ^��bv  ^��c  ��c  ��bv  ^��bv      C  , , B��bv B��c  ���c  ���bv B��bv      C  , ,  ����W�  ����X�  �@��X�  �@��W�  ����W�      C  , ,  �z��W�  �z��X�  �$��X�  �$��W�  �z��W�      C  , ,  ^��W�  ^��X� ��X� ��W�  ^��W�      C  , , B��W� B��X� ���X� ���W� B��W�      C  , ,  ����Vx  ����W"  �x��W"  �x��Vx  ����Vx      C  , ,  ����Vx  ����W"  �\��W"  �\��Vx  ����Vx      C  , ,  ����Vx  ����W"  �@��W"  �@��Vx  ����Vx      C  , ,  �z��Vx  �z��W"  �$��W"  �$��Vx  �z��Vx      C  , ,  ^��Vx  ^��W" ��W" ��Vx  ^��Vx      C  , , B��Vx B��W" ���W" ���Vx B��Vx      C  , ,  ����YH  ����Y�  �@��Y�  �@��YH  ����YH      C  , ,  ����U  ����U�  �x��U�  �x��U  ����U      C  , ,  ����U  ����U�  �\��U�  �\��U  ����U      C  , ,  ����U  ����U�  �@��U�  �@��U  ����U      C  , ,  �z��U  �z��U�  �$��U�  �$��U  �z��U      C  , ,  ^��U  ^��U� ��U� ��U  ^��U      C  , , B��U B��U� ���U� ���U B��U      C  , ,  �z��YH  �z��Y�  �$��Y�  �$��YH  �z��YH      C  , ,  ����S�  ����TR  �x��TR  �x��S�  ����S�      C  , ,  ����S�  ����TR  �\��TR  �\��S�  ����S�      C  , ,  ����S�  ����TR  �@��TR  �@��S�  ����S�      C  , ,  �z��S�  �z��TR  �$��TR  �$��S�  �z��S�      C  , ,  ^��S�  ^��TR ��TR ��S�  ^��S�      C  , , B��S� B��TR ���TR ���S� B��S�      C  , ,  ^��YH  ^��Y� ��Y� ��YH  ^��YH      C  , ,  ����R@  ����R�  �x��R�  �x��R@  ����R@      C  , ,  ����R@  ����R�  �\��R�  �\��R@  ����R@      C  , ,  ����R@  ����R�  �@��R�  �@��R@  ����R@      C  , ,  �z��R@  �z��R�  �$��R�  �$��R@  �z��R@      C  , ,  ^��R@  ^��R� ��R� ��R@  ^��R@      C  , , B��R@ B��R� ���R� ���R@ B��R@      C  , , B��YH B��Y� ���Y� ���YH B��YH      C  , ,  ����P�  ����Q�  �x��Q�  �x��P�  ����P�      C  , ,  ����P�  ����Q�  �\��Q�  �\��P�  ����P�      C  , ,  ����P�  ����Q�  �@��Q�  �@��P�  ����P�      C  , ,  �z��P�  �z��Q�  �$��Q�  �$��P�  �z��P�      C  , ,  ^��P�  ^��Q� ��Q� ��P�  ^��P�      C  , , B��P� B��Q� ���Q� ���P� B��P�      C  , ,  ����YH  ����Y�  �x��Y�  �x��YH  ����YH      C  , ,  ����Op  ����P  �x��P  �x��Op  ����Op      C  , ,  ����Op  ����P  �\��P  �\��Op  ����Op      C  , ,  ����Op  ����P  �@��P  �@��Op  ����Op      C  , ,  �z��Op  �z��P  �$��P  �$��Op  �z��Op      C  , ,  ^��Op  ^��P ��P ��Op  ^��Op      C  , , B��Op B��P ���P ���Op B��Op      C  , ,  ����YH  ����Y�  �\��Y�  �\��YH  ����YH      C  , ,  ����N  ����N�  �x��N�  �x��N  ����N      C  , ,  ����N  ����N�  �\��N�  �\��N  ����N      C  , ,  ����N  ����N�  �@��N�  �@��N  ����N      C  , ,  �z��N  �z��N�  �$��N�  �$��N  �z��N      C  , ,  ^��N  ^��N� ��N� ��N  ^��N      C  , , B��N B��N� ���N� ���N B��N      C  , ,  ����W�  ����X�  �x��X�  �x��W�  ����W�      C  , ,  ����L�  ����MJ  �x��MJ  �x��L�  ����L�      C  , ,  ����L�  ����MJ  �\��MJ  �\��L�  ����L�      C  , ,  ����L�  ����MJ  �@��MJ  �@��L�  ����L�      C  , ,  �z��L�  �z��MJ  �$��MJ  �$��L�  �z��L�      C  , ,  ^��L�  ^��MJ ��MJ ��L�  ^��L�      C  , , B��L� B��MJ ���MJ ���L� B��L�      C  , ,  ����W�  ����X�  �\��X�  �\��W�  ����W�      C  , , ���S� ���TR `��TR `��S� ���S�      C  , , ���S� ���TR D��TR D��S� ���S�      C  , , ~��S� ~��TR (��TR (��S� ~��S�      C  , , b��S� b��TR ��TR ��S� b��S�      C  , , ���YH ���Y� ���Y� ���YH ���YH      C  , , ���YH ���Y� |��Y� |��YH ���YH      C  , , &��Vx &��W" ���W" ���Vx &��Vx      C  , , 	
��Vx 	
��W" 	���W" 	���Vx 	
��Vx      C  , , ���Vx ���W" ���W" ���Vx ���Vx      C  , , ���Vx ���W" |��W" |��Vx ���Vx      C  , , ���Vx ���W" `��W" `��Vx ���Vx      C  , , &��R@ &��R� ���R� ���R@ &��R@      C  , , 	
��R@ 	
��R� 	���R� 	���R@ 	
��R@      C  , , ���R@ ���R� ���R� ���R@ ���R@      C  , , ���R@ ���R� |��R� |��R@ ���R@      C  , , ���R@ ���R� `��R� `��R@ ���R@      C  , , ���R@ ���R� D��R� D��R@ ���R@      C  , , ~��R@ ~��R� (��R� (��R@ ~��R@      C  , , b��R@ b��R� ��R� ��R@ b��R@      C  , , ���Vx ���W" D��W" D��Vx ���Vx      C  , , ~��Vx ~��W" (��W" (��Vx ~��Vx      C  , , b��Vx b��W" ��W" ��Vx b��Vx      C  , , ���YH ���Y� `��Y� `��YH ���YH      C  , , ���YH ���Y� D��Y� D��YH ���YH      C  , , ~��YH ~��Y� (��Y� (��YH ~��YH      C  , , b��YH b��Y� ��Y� ��YH b��YH      C  , , &��P� &��Q� ���Q� ���P� &��P�      C  , , 	
��P� 	
��Q� 	���Q� 	���P� 	
��P�      C  , , ���P� ���Q� ���Q� ���P� ���P�      C  , , ���P� ���Q� |��Q� |��P� ���P�      C  , , ���P� ���Q� `��Q� `��P� ���P�      C  , , ���P� ���Q� D��Q� D��P� ���P�      C  , , ~��P� ~��Q� (��Q� (��P� ~��P�      C  , , b��P� b��Q� ��Q� ��P� b��P�      C  , , &��YH &��Y� ���Y� ���YH &��YH      C  , , 	
��YH 	
��Y� 	���Y� 	���YH 	
��YH      C  , , &��W� &��X� ���X� ���W� &��W�      C  , , &��U &��U� ���U� ���U &��U      C  , , 	
��U 	
��U� 	���U� 	���U 	
��U      C  , , ���U ���U� ���U� ���U ���U      C  , , ���U ���U� |��U� |��U ���U      C  , , &��Op &��P ���P ���Op &��Op      C  , , 	
��Op 	
��P 	���P 	���Op 	
��Op      C  , , ���Op ���P ���P ���Op ���Op      C  , , ���Op ���P |��P |��Op ���Op      C  , , ���Op ���P `��P `��Op ���Op      C  , , ���Op ���P D��P D��Op ���Op      C  , , ~��Op ~��P (��P (��Op ~��Op      C  , , b��Op b��P ��P ��Op b��Op      C  , , ���U ���U� `��U� `��U ���U      C  , , ���U ���U� D��U� D��U ���U      C  , , ~��U ~��U� (��U� (��U ~��U      C  , , b��U b��U� ��U� ��U b��U      C  , , 	
��W� 	
��X� 	���X� 	���W� 	
��W�      C  , , ���W� ���X� ���X� ���W� ���W�      C  , , ���W� ���X� |��X� |��W� ���W�      C  , , &��N &��N� ���N� ���N &��N      C  , , 	
��N 	
��N� 	���N� 	���N 	
��N      C  , , ���N ���N� ���N� ���N ���N      C  , , ���N ���N� |��N� |��N ���N      C  , , ���N ���N� `��N� `��N ���N      C  , , ���N ���N� D��N� D��N ���N      C  , , ~��N ~��N� (��N� (��N ~��N      C  , , b��N b��N� ��N� ��N b��N      C  , , ���W� ���X� `��X� `��W� ���W�      C  , , ���W� ���X� D��X� D��W� ���W�      C  , , ~��W� ~��X� (��X� (��W� ~��W�      C  , , b��W� b��X� ��X� ��W� b��W�      C  , , &��S� &��TR ���TR ���S� &��S�      C  , , 	
��S� 	
��TR 	���TR 	���S� 	
��S�      C  , , ���S� ���TR ���TR ���S� ���S�      C  , , &��L� &��MJ ���MJ ���L� &��L�      C  , , 	
��L� 	
��MJ 	���MJ 	���L� 	
��L�      C  , , ���L� ���MJ ���MJ ���L� ���L�      C  , , ���L� ���MJ |��MJ |��L� ���L�      C  , , ���L� ���MJ `��MJ `��L� ���L�      C  , , ���L� ���MJ D��MJ D��L� ���L�      C  , , ~��L� ~��MJ (��MJ (��L� ~��L�      C  , , b��L� b��MJ ��MJ ��L� b��L�      C  , , ���S� ���TR |��TR |��S� ���S�      C  , , ���c� ���d� �8��d� �8��c� ���c�      C  , , ���o ���o� �8��o� �8��o ���o      C  , , ���bv ���c  �8��c  �8��bv ���bv      C  , , ���j� ���k� �8��k� �8��j� ���j�      C  , , ���p� ���q0 �8��q0 �8��p� ���p�      C  , , ���i~ ���j( �8��j( �8��i~ ���i~      C  , , ���\ ���\� �8��\� �8��\ ���\      C  , , ���m� ���n` �8��n` �8��m� ���m�      C  , , ���h ���h� �8��h� �8��h ���h      C  , , ���Z� ���[Z �8��[Z �8��Z� ���Z�      C  , , ���YH ���Y� �8��Y� �8��YH ���YH      C  , , ���f� ���gX �8��gX �8��f� ���f�      C  , , ���W� ���X� �8��X� �8��W� ���W�      C  , , ���q� ���r� �8��r� �8��q� ���q�      C  , , ���Vx ���W" �8��W" �8��Vx ���Vx      C  , , ���U ���U� �8��U� �8��U ���U      C  , , ���S� ���TR �8��TR �8��S� ���S�      C  , , ���eF ���e� �8��e� �8��eF ���eF      C  , , ���R@ ���R� �8��R� �8��R@ ���R@      C  , , ���P� ���Q� �8��Q� �8��P� ���P�      C  , , ���Op ���P �8��P �8��Op ���Op      C  , , ���N ���N� �8��N� �8��N ���N      C  , , ���lN ���l� �8��l� �8��lN ���lN      C  , , ���L� ���MJ �8��MJ �8��L� ���L�      C  , , Nj��o Nj��o� O��o� O��o Nj��o      C  , , Nj��bv Nj��c  O��c  O��bv Nj��bv      C  , , Nj��j� Nj��k� O��k� O��j� Nj��j�      C  , , Nj��p� Nj��q0 O��q0 O��p� Nj��p�      C  , ,  *��i~  *��j(  ���j(  ���i~  *��i~      C  , , #��i~ #��j( #���j( #���i~ #��i~      C  , , %���i~ %���j( &���j( &���i~ %���i~      C  , , (���i~ (���j( )���j( )���i~ (���i~      C  , , +���i~ +���j( ,d��j( ,d��i~ +���i~      C  , , .���i~ .���j( /H��j( /H��i~ .���i~      C  , , 1���i~ 1���j( 2,��j( 2,��i~ 1���i~      C  , , 4f��i~ 4f��j( 5��j( 5��i~ 4f��i~      C  , , 7J��i~ 7J��j( 7���j( 7���i~ 7J��i~      C  , , :.��i~ :.��j( :���j( :���i~ :.��i~      C  , , =��i~ =��j( =���j( =���i~ =��i~      C  , , ?���i~ ?���j( @���j( @���i~ ?���i~      C  , , B���i~ B���j( C���j( C���i~ B���i~      C  , , E���i~ E���j( Fh��j( Fh��i~ E���i~      C  , , H���i~ H���j( IL��j( IL��i~ H���i~      C  , , K���i~ K���j( L0��j( L0��i~ K���i~      C  , , Nj��i~ Nj��j( O��j( O��i~ Nj��i~      C  , , QN��i~ QN��j( Q���j( Q���i~ QN��i~      C  , , T2��i~ T2��j( T���j( T���i~ T2��i~      C  , , W��i~ W��j( W���j( W���i~ W��i~      C  , , Y���i~ Y���j( Z���j( Z���i~ Y���i~      C  , , \���i~ \���j( ]���j( ]���i~ \���i~      C  , , _���i~ _���j( `l��j( `l��i~ _���i~      C  , , b���i~ b���j( cP��j( cP��i~ b���i~      C  , , e���i~ e���j( f4��j( f4��i~ e���i~      C  , , hn��i~ hn��j( i��j( i��i~ hn��i~      C  , , kR��i~ kR��j( k���j( k���i~ kR��i~      C  , , n6��i~ n6��j( n���j( n���i~ n6��i~      C  , , q��i~ q��j( q���j( q���i~ q��i~      C  , , s���i~ s���j( t���j( t���i~ s���i~      C  , , v���i~ v���j( w���j( w���i~ v���i~      C  , , y���i~ y���j( zp��j( zp��i~ y���i~      C  , , |���i~ |���j( }T��j( }T��i~ |���i~      C  , , Nj��m� Nj��n` O��n` O��m� Nj��m�      C  , , Nj��\ Nj��\� O��\� O��\ Nj��\      C  , , Nj��h Nj��h� O��h� O��h Nj��h      C  , , Nj��Z� Nj��[Z O��[Z O��Z� Nj��Z�      C  , , Nj��q� Nj��r� O��r� O��q� Nj��q�      C  , , Nj��YH Nj��Y� O��Y� O��YH Nj��YH      C  , , Nj��f� Nj��gX O��gX O��f� Nj��f�      C  , , Nj��W� Nj��X� O��X� O��W� Nj��W�      C  , , Nj��Vx Nj��W" O��W" O��Vx Nj��Vx      C  , , Nj��U Nj��U� O��U� O��U Nj��U      C  , , Nj��eF Nj��e� O��e� O��eF Nj��eF      C  , , Nj��S� Nj��TR O��TR O��S� Nj��S�      C  , , Nj��c� Nj��d� O��d� O��c� Nj��c�      C  , , Nj��R@ Nj��R� O��R� O��R@ Nj��R@      C  , , Nj��P� Nj��Q� O��Q� O��P� Nj��P�      C  , , Nj��Op Nj��P O��P O��Op Nj��Op      C  , , Nj��lN Nj��l� O��l� O��lN Nj��lN      C  , , Nj��N Nj��N� O��N� O��N Nj��N      C  , , Nj��L� Nj��MJ O��MJ O��L� Nj��L�      C  , , e���o e���o� f4��o� f4��o e���o      C  , , hn��o hn��o� i��o� i��o hn��o      C  , , kR��o kR��o� k���o� k���o kR��o      C  , , n6��o n6��o� n���o� n���o n6��o      C  , , q��o q��o� q���o� q���o q��o      C  , , s���o s���o� t���o� t���o s���o      C  , , v���o v���o� w���o� w���o v���o      C  , , y���o y���o� zp��o� zp��o y���o      C  , , |���o |���o� }T��o� }T��o |���o      C  , , QN��o QN��o� Q���o� Q���o QN��o      C  , , T2��o T2��o� T���o� T���o T2��o      C  , , QN��j� QN��k� Q���k� Q���j� QN��j�      C  , , T2��j� T2��k� T���k� T���j� T2��j�      C  , , W��j� W��k� W���k� W���j� W��j�      C  , , Y���j� Y���k� Z���k� Z���j� Y���j�      C  , , \���j� \���k� ]���k� ]���j� \���j�      C  , , _���j� _���k� `l��k� `l��j� _���j�      C  , , b���j� b���k� cP��k� cP��j� b���j�      C  , , e���j� e���k� f4��k� f4��j� e���j�      C  , , hn��j� hn��k� i��k� i��j� hn��j�      C  , , kR��j� kR��k� k���k� k���j� kR��j�      C  , , n6��j� n6��k� n���k� n���j� n6��j�      C  , , q��j� q��k� q���k� q���j� q��j�      C  , , s���j� s���k� t���k� t���j� s���j�      C  , , v���j� v���k� w���k� w���j� v���j�      C  , , y���j� y���k� zp��k� zp��j� y���j�      C  , , |���j� |���k� }T��k� }T��j� |���j�      C  , , W��o W��o� W���o� W���o W��o      C  , , QN��p� QN��q0 Q���q0 Q���p� QN��p�      C  , , T2��p� T2��q0 T���q0 T���p� T2��p�      C  , , QN��m� QN��n` Q���n` Q���m� QN��m�      C  , , T2��m� T2��n` T���n` T���m� T2��m�      C  , , W��m� W��n` W���n` W���m� W��m�      C  , , Y���m� Y���n` Z���n` Z���m� Y���m�      C  , , \���m� \���n` ]���n` ]���m� \���m�      C  , , _���m� _���n` `l��n` `l��m� _���m�      C  , , b���m� b���n` cP��n` cP��m� b���m�      C  , , e���m� e���n` f4��n` f4��m� e���m�      C  , , hn��m� hn��n` i��n` i��m� hn��m�      C  , , kR��m� kR��n` k���n` k���m� kR��m�      C  , , n6��m� n6��n` n���n` n���m� n6��m�      C  , , q��m� q��n` q���n` q���m� q��m�      C  , , s���m� s���n` t���n` t���m� s���m�      C  , , v���m� v���n` w���n` w���m� v���m�      C  , , y���m� y���n` zp��n` zp��m� y���m�      C  , , |���m� |���n` }T��n` }T��m� |���m�      C  , , W��p� W��q0 W���q0 W���p� W��p�      C  , , Y���p� Y���q0 Z���q0 Z���p� Y���p�      C  , , \���p� \���q0 ]���q0 ]���p� \���p�      C  , , _���p� _���q0 `l��q0 `l��p� _���p�      C  , , b���p� b���q0 cP��q0 cP��p� b���p�      C  , , QN��q� QN��r� Q���r� Q���q� QN��q�      C  , , T2��q� T2��r� T���r� T���q� T2��q�      C  , , W��q� W��r� W���r� W���q� W��q�      C  , , Y���q� Y���r� Z���r� Z���q� Y���q�      C  , , \���q� \���r� ]���r� ]���q� \���q�      C  , , _���q� _���r� `l��r� `l��q� _���q�      C  , , b���q� b���r� cP��r� cP��q� b���q�      C  , , e���q� e���r� f4��r� f4��q� e���q�      C  , , hn��q� hn��r� i��r� i��q� hn��q�      C  , , kR��q� kR��r� k���r� k���q� kR��q�      C  , , n6��q� n6��r� n���r� n���q� n6��q�      C  , , e���p� e���q0 f4��q0 f4��p� e���p�      C  , , hn��p� hn��q0 i��q0 i��p� hn��p�      C  , , q��q� q��r� q���r� q���q� q��q�      C  , , s���q� s���r� t���r� t���q� s���q�      C  , , v���q� v���r� w���r� w���q� v���q�      C  , , y���q� y���r� zp��r� zp��q� y���q�      C  , , |���q� |���r� }T��r� }T��q� |���q�      C  , , kR��p� kR��q0 k���q0 k���p� kR��p�      C  , , n6��p� n6��q0 n���q0 n���p� n6��p�      C  , , q��p� q��q0 q���q0 q���p� q��p�      C  , , s���p� s���q0 t���q0 t���p� s���p�      C  , , v���p� v���q0 w���q0 w���p� v���p�      C  , , y���p� y���q0 zp��q0 zp��p� y���p�      C  , , |���p� |���q0 }T��q0 }T��p� |���p�      C  , , Y���o Y���o� Z���o� Z���o Y���o      C  , , \���o \���o� ]���o� ]���o \���o      C  , , QN��lN QN��l� Q���l� Q���lN QN��lN      C  , , T2��lN T2��l� T���l� T���lN T2��lN      C  , , W��lN W��l� W���l� W���lN W��lN      C  , , Y���lN Y���l� Z���l� Z���lN Y���lN      C  , , \���lN \���l� ]���l� ]���lN \���lN      C  , , _���lN _���l� `l��l� `l��lN _���lN      C  , , b���lN b���l� cP��l� cP��lN b���lN      C  , , e���lN e���l� f4��l� f4��lN e���lN      C  , , hn��lN hn��l� i��l� i��lN hn��lN      C  , , kR��lN kR��l� k���l� k���lN kR��lN      C  , , _���o _���o� `l��o� `l��o _���o      C  , , n6��lN n6��l� n���l� n���lN n6��lN      C  , , q��lN q��l� q���l� q���lN q��lN      C  , , s���lN s���l� t���l� t���lN s���lN      C  , , v���lN v���l� w���l� w���lN v���lN      C  , , y���lN y���l� zp��l� zp��lN y���lN      C  , , |���lN |���l� }T��l� }T��lN |���lN      C  , , b���o b���o� cP��o� cP��o b���o      C  , , 1���j� 1���k� 2,��k� 2,��j� 1���j�      C  , , 4f��j� 4f��k� 5��k� 5��j� 4f��j�      C  , , 7J��j� 7J��k� 7���k� 7���j� 7J��j�      C  , , :.��j� :.��k� :���k� :���j� :.��j�      C  , , =��j� =��k� =���k� =���j� =��j�      C  , , ?���j� ?���k� @���k� @���j� ?���j�      C  , , B���j� B���k� C���k� C���j� B���j�      C  , , E���j� E���k� Fh��k� Fh��j� E���j�      C  , , H���j� H���k� IL��k� IL��j� H���j�      C  , , K���j� K���k� L0��k� L0��j� K���j�      C  , , %���o %���o� &���o� &���o %���o      C  , , (���o (���o� )���o� )���o (���o      C  , , +���o +���o� ,d��o� ,d��o +���o      C  , , .���o .���o� /H��o� /H��o .���o      C  , , 1���o 1���o� 2,��o� 2,��o 1���o      C  , , 4f��o 4f��o� 5��o� 5��o 4f��o      C  , , 7J��o 7J��o� 7���o� 7���o 7J��o      C  , ,  *��q�  *��r�  ���r�  ���q�  *��q�      C  , , #��q� #��r� #���r� #���q� #��q�      C  , , %���q� %���r� &���r� &���q� %���q�      C  , , (���q� (���r� )���r� )���q� (���q�      C  , , +���q� +���r� ,d��r� ,d��q� +���q�      C  , , .���q� .���r� /H��r� /H��q� .���q�      C  , , 1���q� 1���r� 2,��r� 2,��q� 1���q�      C  , , 4f��q� 4f��r� 5��r� 5��q� 4f��q�      C  , , 7J��q� 7J��r� 7���r� 7���q� 7J��q�      C  , , :.��q� :.��r� :���r� :���q� :.��q�      C  , , =��q� =��r� =���r� =���q� =��q�      C  , , ?���q� ?���r� @���r� @���q� ?���q�      C  , , B���q� B���r� C���r� C���q� B���q�      C  , , E���q� E���r� Fh��r� Fh��q� E���q�      C  , , H���q� H���r� IL��r� IL��q� H���q�      C  , , K���q� K���r� L0��r� L0��q� K���q�      C  , , :.��o :.��o� :���o� :���o :.��o      C  , , =��o =��o� =���o� =���o =��o      C  , , ?���o ?���o� @���o� @���o ?���o      C  , , B���o B���o� C���o� C���o B���o      C  , , E���o E���o� Fh��o� Fh��o E���o      C  , , H���o H���o� IL��o� IL��o H���o      C  , , K���o K���o� L0��o� L0��o K���o      C  , ,  *��o  *��o�  ���o�  ���o  *��o      C  , , #��o #��o� #���o� #���o #��o      C  , ,  *��j�  *��k�  ���k�  ���j�  *��j�      C  , ,  *��p�  *��q0  ���q0  ���p�  *��p�      C  , , #��p� #��q0 #���q0 #���p� #��p�      C  , , %���p� %���q0 &���q0 &���p� %���p�      C  , , (���p� (���q0 )���q0 )���p� (���p�      C  , , +���p� +���q0 ,d��q0 ,d��p� +���p�      C  , , .���p� .���q0 /H��q0 /H��p� .���p�      C  , , 1���p� 1���q0 2,��q0 2,��p� 1���p�      C  , , 4f��p� 4f��q0 5��q0 5��p� 4f��p�      C  , , 7J��p� 7J��q0 7���q0 7���p� 7J��p�      C  , , :.��p� :.��q0 :���q0 :���p� :.��p�      C  , , =��p� =��q0 =���q0 =���p� =��p�      C  , , ?���p� ?���q0 @���q0 @���p� ?���p�      C  , , B���p� B���q0 C���q0 C���p� B���p�      C  , , E���p� E���q0 Fh��q0 Fh��p� E���p�      C  , , H���p� H���q0 IL��q0 IL��p� H���p�      C  , , K���p� K���q0 L0��q0 L0��p� K���p�      C  , , #��j� #��k� #���k� #���j� #��j�      C  , ,  *��lN  *��l�  ���l�  ���lN  *��lN      C  , , #��lN #��l� #���l� #���lN #��lN      C  , , %���lN %���l� &���l� &���lN %���lN      C  , , (���lN (���l� )���l� )���lN (���lN      C  , , +���lN +���l� ,d��l� ,d��lN +���lN      C  , , .���lN .���l� /H��l� /H��lN .���lN      C  , , 1���lN 1���l� 2,��l� 2,��lN 1���lN      C  , , 4f��lN 4f��l� 5��l� 5��lN 4f��lN      C  , , 7J��lN 7J��l� 7���l� 7���lN 7J��lN      C  , , :.��lN :.��l� :���l� :���lN :.��lN      C  , , =��lN =��l� =���l� =���lN =��lN      C  , , ?���lN ?���l� @���l� @���lN ?���lN      C  , , %���j� %���k� &���k� &���j� %���j�      C  , , B���lN B���l� C���l� C���lN B���lN      C  , , E���lN E���l� Fh��l� Fh��lN E���lN      C  , , H���lN H���l� IL��l� IL��lN H���lN      C  , , K���lN K���l� L0��l� L0��lN K���lN      C  , ,  *��m�  *��n`  ���n`  ���m�  *��m�      C  , , #��m� #��n` #���n` #���m� #��m�      C  , , %���m� %���n` &���n` &���m� %���m�      C  , , (���m� (���n` )���n` )���m� (���m�      C  , , +���m� +���n` ,d��n` ,d��m� +���m�      C  , , .���m� .���n` /H��n` /H��m� .���m�      C  , , 1���m� 1���n` 2,��n` 2,��m� 1���m�      C  , , 4f��m� 4f��n` 5��n` 5��m� 4f��m�      C  , , 7J��m� 7J��n` 7���n` 7���m� 7J��m�      C  , , :.��m� :.��n` :���n` :���m� :.��m�      C  , , =��m� =��n` =���n` =���m� =��m�      C  , , ?���m� ?���n` @���n` @���m� ?���m�      C  , , B���m� B���n` C���n` C���m� B���m�      C  , , E���m� E���n` Fh��n` Fh��m� E���m�      C  , , H���m� H���n` IL��n` IL��m� H���m�      C  , , K���m� K���n` L0��n` L0��m� K���m�      C  , , (���j� (���k� )���k� )���j� (���j�      C  , , +���j� +���k� ,d��k� ,d��j� +���j�      C  , , .���j� .���k� /H��k� /H��j� .���j�      C  , ,  *��Z�  *��[Z  ���[Z  ���Z�  *��Z�      C  , , #��Z� #��[Z #���[Z #���Z� #��Z�      C  , , %���Z� %���[Z &���[Z &���Z� %���Z�      C  , , (���Z� (���[Z )���[Z )���Z� (���Z�      C  , , +���Z� +���[Z ,d��[Z ,d��Z� +���Z�      C  , , .���Z� .���[Z /H��[Z /H��Z� .���Z�      C  , , 1���Z� 1���[Z 2,��[Z 2,��Z� 1���Z�      C  , , 4f��Z� 4f��[Z 5��[Z 5��Z� 4f��Z�      C  , , 7J��Z� 7J��[Z 7���[Z 7���Z� 7J��Z�      C  , , :.��Z� :.��[Z :���[Z :���Z� :.��Z�      C  , , =��Z� =��[Z =���[Z =���Z� =��Z�      C  , , ?���Z� ?���[Z @���[Z @���Z� ?���Z�      C  , , B���Z� B���[Z C���[Z C���Z� B���Z�      C  , , E���Z� E���[Z Fh��[Z Fh��Z� E���Z�      C  , , H���Z� H���[Z IL��[Z IL��Z� H���Z�      C  , , K���Z� K���[Z L0��[Z L0��Z� K���Z�      C  , , 5���`U 5���`� 6���`� 6���`U 5���`U      C  , , 5���^9 5���^� 6���^� 6���^9 5���^9      C  , , 7J��h 7J��h� 7���h� 7���h 7J��h      C  , , :.��h :.��h� :���h� :���h :.��h      C  , , =��h =��h� =���h� =���h =��h      C  , , ?���h ?���h� @���h� @���h ?���h      C  , , B���h B���h� C���h� C���h B���h      C  , , E���h E���h� Fh��h� Fh��h E���h      C  , , H���h H���h� IL��h� IL��h H���h      C  , , :.��c� :.��d� :���d� :���c� :.��c�      C  , , K���h K���h� L0��h� L0��h K���h      C  , , 7J��c� 7J��d� 7���d� 7���c� 7J��c�      C  , , 8���^9 8���^� 9f��^� 9f��^9 8���^9      C  , , ;���^9 ;���^� <J��^� <J��^9 ;���^9      C  , , >���^9 >���^� ?.��^� ?.��^9 >���^9      C  , , Ah��^9 Ah��^� B��^� B��^9 Ah��^9      C  , , DL��^9 DL��^� D���^� D���^9 DL��^9      C  , , G0��^9 G0��^� G���^� G���^9 G0��^9      C  , , =��c� =��d� =���d� =���c� =��c�      C  , , J��^9 J��^� J���^� J���^9 J��^9      C  , , L���^9 L���^� M���^� M���^9 L���^9      C  , , 8���`U 8���`� 9f��`� 9f��`U 8���`U      C  , , ;���`U ;���`� <J��`� <J��`U ;���`U      C  , , >���`U >���`� ?.��`� ?.��`U >���`U      C  , , Ah��`U Ah��`� B��`� B��`U Ah��`U      C  , , DL��`U DL��`� D���`� D���`U DL��`U      C  , , G0��`U G0��`� G���`� G���`U G0��`U      C  , , J��`U J��`� J���`� J���`U J��`U      C  , , L���`U L���`� M���`� M���`U L���`U      C  , , 7J��f� 7J��gX 7���gX 7���f� 7J��f�      C  , , :.��f� :.��gX :���gX :���f� :.��f�      C  , , =��f� =��gX =���gX =���f� =��f�      C  , , ?���f� ?���gX @���gX @���f� ?���f�      C  , , B���f� B���gX C���gX C���f� B���f�      C  , , E���f� E���gX Fh��gX Fh��f� E���f�      C  , , H���f� H���gX IL��gX IL��f� H���f�      C  , , K���f� K���gX L0��gX L0��f� K���f�      C  , , E���bv E���c  Fh��c  Fh��bv E���bv      C  , , ?���c� ?���d� @���d� @���c� ?���c�      C  , , H���bv H���c  IL��c  IL��bv H���bv      C  , , B���c� B���d� C���d� C���c� B���c�      C  , , K���bv K���c  L0��c  L0��bv K���bv      C  , , E���c� E���d� Fh��d� Fh��c� E���c�      C  , , H���c� H���d� IL��d� IL��c� H���c�      C  , , 7J��eF 7J��e� 7���e� 7���eF 7J��eF      C  , , :.��eF :.��e� :���e� :���eF :.��eF      C  , , =��eF =��e� =���e� =���eF =��eF      C  , , ?���eF ?���e� @���e� @���eF ?���eF      C  , , B���eF B���e� C���e� C���eF B���eF      C  , , K���c� K���d� L0��d� L0��c� K���c�      C  , , E���eF E���e� Fh��e� Fh��eF E���eF      C  , , H���eF H���e� IL��e� IL��eF H���eF      C  , , K���eF K���e� L0��e� L0��eF K���eF      C  , , 7J��bv 7J��c  7���c  7���bv 7J��bv      C  , , :.��bv :.��c  :���c  :���bv :.��bv      C  , , =��bv =��c  =���c  =���bv =��bv      C  , , ?���bv ?���c  @���c  @���bv ?���bv      C  , , B���bv B���c  C���c  C���bv B���bv      C  , , 7J��\ 7J��\� 7���\� 7���\ 7J��\      C  , , :.��\ :.��\� :���\� :���\ :.��\      C  , , =��\ =��\� =���\� =���\ =��\      C  , , ?���\ ?���\� @���\� @���\ ?���\      C  , , B���\ B���\� C���\� C���\ B���\      C  , , E���\ E���\� Fh��\� Fh��\ E���\      C  , , H���\ H���\� IL��\� IL��\ H���\      C  , , K���\ K���\� L0��\� L0��\ K���\      C  , , #��c� #��d� #���d� #���c� #��c�      C  , ,  *��bv  *��c   ���c   ���bv  *��bv      C  , , .���c� .���d� /H��d� /H��c� .���c�      C  , , #��bv #��c  #���c  #���bv #��bv      C  , ,  *��f�  *��gX  ���gX  ���f�  *��f�      C  , ,  *��eF  *��e�  ���e�  ���eF  *��eF      C  , , #��eF #��e� #���e� #���eF #��eF      C  , , %���eF %���e� &���e� &���eF %���eF      C  , , (���eF (���e� )���e� )���eF (���eF      C  , , +���eF +���e� ,d��e� ,d��eF +���eF      C  , , .���eF .���e� /H��e� /H��eF .���eF      C  , , 1���eF 1���e� 2,��e� 2,��eF 1���eF      C  , , 4f��eF 4f��e� 5��e� 5��eF 4f��eF      C  , , #��f� #��gX #���gX #���f� #��f�      C  , , %���f� %���gX &���gX &���f� %���f�      C  , , (���f� (���gX )���gX )���f� (���f�      C  , , +���f� +���gX ,d��gX ,d��f� +���f�      C  , , .���f� .���gX /H��gX /H��f� .���f�      C  , , %���bv %���c  &���c  &���bv %���bv      C  , , 1���f� 1���gX 2,��gX 2,��f� 1���f�      C  , , 4f��f� 4f��gX 5��gX 5��f� 4f��f�      C  , , ���^9 ���^� b��^� b��^9 ���^9      C  , , !���^9 !���^� "F��^� "F��^9 !���^9      C  , , (���bv (���c  )���c  )���bv (���bv      C  , , +���bv +���c  ,d��c  ,d��bv +���bv      C  , , .���bv .���c  /H��c  /H��bv .���bv      C  , , 1���bv 1���c  2,��c  2,��bv 1���bv      C  , , 4f��bv 4f��c  5��c  5��bv 4f��bv      C  , , $���^9 $���^� %*��^� %*��^9 $���^9      C  , , 'd��^9 'd��^� (��^� (��^9 'd��^9      C  , , *H��^9 *H��^� *���^� *���^9 *H��^9      C  , , -,��^9 -,��^� -���^� -���^9 -,��^9      C  , , 0��^9 0��^� 0���^� 0���^9 0��^9      C  , , (���c� (���d� )���d� )���c� (���c�      C  , , ���`U ���`� b��`� b��`U ���`U      C  , , !���`U !���`� "F��`� "F��`U !���`U      C  , , $���`U $���`� %*��`� %*��`U $���`U      C  , , 'd��`U 'd��`� (��`� (��`U 'd��`U      C  , ,  *��\  *��\�  ���\�  ���\  *��\      C  , , #��\ #��\� #���\� #���\ #��\      C  , , %���\ %���\� &���\� &���\ %���\      C  , , (���\ (���\� )���\� )���\ (���\      C  , , +���\ +���\� ,d��\� ,d��\ +���\      C  , , .���\ .���\� /H��\� /H��\ .���\      C  , , 1���\ 1���\� 2,��\� 2,��\ 1���\      C  , , 4f��\ 4f��\� 5��\� 5��\ 4f��\      C  , , 2���^9 2���^� 3���^� 3���^9 2���^9      C  , , 0��`U 0��`� 0���`� 0���`U 0��`U      C  , , +���c� +���d� ,d��d� ,d��c� +���c�      C  , , -,��`U -,��`� -���`� -���`U -,��`U      C  , , 2���`U 2���`� 3���`� 3���`U 2���`U      C  , , 4f��h 4f��h� 5��h� 5��h 4f��h      C  , ,  *��c�  *��d�  ���d�  ���c�  *��c�      C  , , %���c� %���d� &���d� &���c� %���c�      C  , , *H��`U *H��`� *���`� *���`U *H��`U      C  , , 1���c� 1���d� 2,��d� 2,��c� 1���c�      C  , , 4f��c� 4f��d� 5��d� 5��c� 4f��c�      C  , ,  *��h  *��h�  ���h�  ���h  *��h      C  , , #��h #��h� #���h� #���h #��h      C  , , %���h %���h� &���h� &���h %���h      C  , , (���h (���h� )���h� )���h (���h      C  , , +���h +���h� ,d��h� ,d��h +���h      C  , , .���h .���h� /H��h� /H��h .���h      C  , , 1���h 1���h� 2,��h� 2,��h 1���h      C  , , .���Vx .���W" /H��W" /H��Vx .���Vx      C  , , 1���Vx 1���W" 2,��W" 2,��Vx 1���Vx      C  , ,  *��R@  *��R�  ���R�  ���R@  *��R@      C  , , #��R@ #��R� #���R� #���R@ #��R@      C  , , %���R@ %���R� &���R� &���R@ %���R@      C  , , (���R@ (���R� )���R� )���R@ (���R@      C  , , +���R@ +���R� ,d��R� ,d��R@ +���R@      C  , , .���R@ .���R� /H��R� /H��R@ .���R@      C  , , 1���R@ 1���R� 2,��R� 2,��R@ 1���R@      C  , , 4f��R@ 4f��R� 5��R� 5��R@ 4f��R@      C  , , 4f��Vx 4f��W" 5��W" 5��Vx 4f��Vx      C  , ,  *��P�  *��Q�  ���Q�  ���P�  *��P�      C  , , #��P� #��Q� #���Q� #���P� #��P�      C  , , %���P� %���Q� &���Q� &���P� %���P�      C  , , (���P� (���Q� )���Q� )���P� (���P�      C  , , +���P� +���Q� ,d��Q� ,d��P� +���P�      C  , , .���P� .���Q� /H��Q� /H��P� .���P�      C  , , 1���P� 1���Q� 2,��Q� 2,��P� 1���P�      C  , , 4f��P� 4f��Q� 5��Q� 5��P� 4f��P�      C  , ,  *��W�  *��X�  ���X�  ���W�  *��W�      C  , , #��W� #��X� #���X� #���W� #��W�      C  , , %���W� %���X� &���X� &���W� %���W�      C  , , (���W� (���X� )���X� )���W� (���W�      C  , , +���W� +���X� ,d��X� ,d��W� +���W�      C  , , .���W� .���X� /H��X� /H��W� .���W�      C  , , 1���W� 1���X� 2,��X� 2,��W� 1���W�      C  , , 4f��W� 4f��X� 5��X� 5��W� 4f��W�      C  , , 4f��YH 4f��Y� 5��Y� 5��YH 4f��YH      C  , ,  *��YH  *��Y�  ���Y�  ���YH  *��YH      C  , , #��YH #��Y� #���Y� #���YH #��YH      C  , , %���YH %���Y� &���Y� &���YH %���YH      C  , , (���YH (���Y� )���Y� )���YH (���YH      C  , ,  *��Op  *��P  ���P  ���Op  *��Op      C  , , #��Op #��P #���P #���Op #��Op      C  , , %���Op %���P &���P &���Op %���Op      C  , , (���Op (���P )���P )���Op (���Op      C  , , +���Op +���P ,d��P ,d��Op +���Op      C  , , .���Op .���P /H��P /H��Op .���Op      C  , , 1���Op 1���P 2,��P 2,��Op 1���Op      C  , , 4f��Op 4f��P 5��P 5��Op 4f��Op      C  , , +���YH +���Y� ,d��Y� ,d��YH +���YH      C  , , .���YH .���Y� /H��Y� /H��YH .���YH      C  , ,  *��U  *��U�  ���U�  ���U  *��U      C  , , #��U #��U� #���U� #���U #��U      C  , , %���U %���U� &���U� &���U %���U      C  , , (���U (���U� )���U� )���U (���U      C  , , +���U +���U� ,d��U� ,d��U +���U      C  , , .���U .���U� /H��U� /H��U .���U      C  , , 1���U 1���U� 2,��U� 2,��U 1���U      C  , , 4f��U 4f��U� 5��U� 5��U 4f��U      C  , , 1���YH 1���Y� 2,��Y� 2,��YH 1���YH      C  , ,  *��Vx  *��W"  ���W"  ���Vx  *��Vx      C  , , #��Vx #��W" #���W" #���Vx #��Vx      C  , , %���Vx %���W" &���W" &���Vx %���Vx      C  , , (���Vx (���W" )���W" )���Vx (���Vx      C  , , +���Vx +���W" ,d��W" ,d��Vx +���Vx      C  , ,  *��N  *��N�  ���N�  ���N  *��N      C  , , #��N #��N� #���N� #���N #��N      C  , , %���N %���N� &���N� &���N %���N      C  , , (���N (���N� )���N� )���N (���N      C  , , +���N +���N� ,d��N� ,d��N +���N      C  , , .���N .���N� /H��N� /H��N .���N      C  , , 1���N 1���N� 2,��N� 2,��N 1���N      C  , , 4f��N 4f��N� 5��N� 5��N 4f��N      C  , ,  *��S�  *��TR  ���TR  ���S�  *��S�      C  , , #��S� #��TR #���TR #���S� #��S�      C  , , %���S� %���TR &���TR &���S� %���S�      C  , , (���S� (���TR )���TR )���S� (���S�      C  , , +���S� +���TR ,d��TR ,d��S� +���S�      C  , , .���S� .���TR /H��TR /H��S� .���S�      C  , , 1���S� 1���TR 2,��TR 2,��S� 1���S�      C  , ,  *��L�  *��MJ  ���MJ  ���L�  *��L�      C  , , #��L� #��MJ #���MJ #���L� #��L�      C  , , %���L� %���MJ &���MJ &���L� %���L�      C  , , (���L� (���MJ )���MJ )���L� (���L�      C  , , +���L� +���MJ ,d��MJ ,d��L� +���L�      C  , , .���L� .���MJ /H��MJ /H��L� .���L�      C  , , 1���L� 1���MJ 2,��MJ 2,��L� 1���L�      C  , , 4f��L� 4f��MJ 5��MJ 5��L� 4f��L�      C  , , 4f��S� 4f��TR 5��TR 5��S� 4f��S�      C  , , B���YH B���Y� C���Y� C���YH B���YH      C  , , E���YH E���Y� Fh��Y� Fh��YH E���YH      C  , , H���YH H���Y� IL��Y� IL��YH H���YH      C  , , 7J��W� 7J��X� 7���X� 7���W� 7J��W�      C  , , :.��W� :.��X� :���X� :���W� :.��W�      C  , , =��W� =��X� =���X� =���W� =��W�      C  , , ?���W� ?���X� @���X� @���W� ?���W�      C  , , B���W� B���X� C���X� C���W� B���W�      C  , , 7J��S� 7J��TR 7���TR 7���S� 7J��S�      C  , , :.��S� :.��TR :���TR :���S� :.��S�      C  , , =��S� =��TR =���TR =���S� =��S�      C  , , ?���S� ?���TR @���TR @���S� ?���S�      C  , , B���S� B���TR C���TR C���S� B���S�      C  , , E���S� E���TR Fh��TR Fh��S� E���S�      C  , , H���S� H���TR IL��TR IL��S� H���S�      C  , , K���S� K���TR L0��TR L0��S� K���S�      C  , , 7J��Op 7J��P 7���P 7���Op 7J��Op      C  , , :.��Op :.��P :���P :���Op :.��Op      C  , , =��Op =��P =���P =���Op =��Op      C  , , ?���Op ?���P @���P @���Op ?���Op      C  , , B���Op B���P C���P C���Op B���Op      C  , , E���Op E���P Fh��P Fh��Op E���Op      C  , , H���Op H���P IL��P IL��Op H���Op      C  , , K���Op K���P L0��P L0��Op K���Op      C  , , E���W� E���X� Fh��X� Fh��W� E���W�      C  , , H���W� H���X� IL��X� IL��W� H���W�      C  , , K���W� K���X� L0��X� L0��W� K���W�      C  , , 7J��Vx 7J��W" 7���W" 7���Vx 7J��Vx      C  , , :.��Vx :.��W" :���W" :���Vx :.��Vx      C  , , =��Vx =��W" =���W" =���Vx =��Vx      C  , , ?���Vx ?���W" @���W" @���Vx ?���Vx      C  , , B���Vx B���W" C���W" C���Vx B���Vx      C  , , E���Vx E���W" Fh��W" Fh��Vx E���Vx      C  , , H���Vx H���W" IL��W" IL��Vx H���Vx      C  , , 7J��R@ 7J��R� 7���R� 7���R@ 7J��R@      C  , , :.��R@ :.��R� :���R� :���R@ :.��R@      C  , , =��R@ =��R� =���R� =���R@ =��R@      C  , , ?���R@ ?���R� @���R� @���R@ ?���R@      C  , , B���R@ B���R� C���R� C���R@ B���R@      C  , , E���R@ E���R� Fh��R� Fh��R@ E���R@      C  , , H���R@ H���R� IL��R� IL��R@ H���R@      C  , , K���R@ K���R� L0��R� L0��R@ K���R@      C  , , 7J��U 7J��U� 7���U� 7���U 7J��U      C  , , :.��U :.��U� :���U� :���U :.��U      C  , , =��U =��U� =���U� =���U =��U      C  , , ?���U ?���U� @���U� @���U ?���U      C  , , B���U B���U� C���U� C���U B���U      C  , , E���U E���U� Fh��U� Fh��U E���U      C  , , 7J��N 7J��N� 7���N� 7���N 7J��N      C  , , :.��N :.��N� :���N� :���N :.��N      C  , , =��N =��N� =���N� =���N =��N      C  , , ?���N ?���N� @���N� @���N ?���N      C  , , B���N B���N� C���N� C���N B���N      C  , , E���N E���N� Fh��N� Fh��N E���N      C  , , H���N H���N� IL��N� IL��N H���N      C  , , K���N K���N� L0��N� L0��N K���N      C  , , H���U H���U� IL��U� IL��U H���U      C  , , K���U K���U� L0��U� L0��U K���U      C  , , K���Vx K���W" L0��W" L0��Vx K���Vx      C  , , 7J��P� 7J��Q� 7���Q� 7���P� 7J��P�      C  , , :.��P� :.��Q� :���Q� :���P� :.��P�      C  , , =��P� =��Q� =���Q� =���P� =��P�      C  , , ?���P� ?���Q� @���Q� @���P� ?���P�      C  , , B���P� B���Q� C���Q� C���P� B���P�      C  , , E���P� E���Q� Fh��Q� Fh��P� E���P�      C  , , H���P� H���Q� IL��Q� IL��P� H���P�      C  , , K���P� K���Q� L0��Q� L0��P� K���P�      C  , , K���YH K���Y� L0��Y� L0��YH K���YH      C  , , 7J��YH 7J��Y� 7���Y� 7���YH 7J��YH      C  , , :.��YH :.��Y� :���Y� :���YH :.��YH      C  , , =��YH =��Y� =���Y� =���YH =��YH      C  , , 7J��L� 7J��MJ 7���MJ 7���L� 7J��L�      C  , , :.��L� :.��MJ :���MJ :���L� :.��L�      C  , , =��L� =��MJ =���MJ =���L� =��L�      C  , , ?���L� ?���MJ @���MJ @���L� ?���L�      C  , , B���L� B���MJ C���MJ C���L� B���L�      C  , , E���L� E���MJ Fh��MJ Fh��L� E���L�      C  , , H���L� H���MJ IL��MJ IL��L� H���L�      C  , , K���L� K���MJ L0��MJ L0��L� K���L�      C  , , ?���YH ?���Y� @���Y� @���YH ?���YH      C  , , f���`U f���`� g���`� g���`U f���`U      C  , , f���^9 f���^� g���^� g���^9 f���^9      C  , , QN��Z� QN��[Z Q���[Z Q���Z� QN��Z�      C  , , T2��Z� T2��[Z T���[Z T���Z� T2��Z�      C  , , W��Z� W��[Z W���[Z W���Z� W��Z�      C  , , Y���Z� Y���[Z Z���[Z Z���Z� Y���Z�      C  , , \���Z� \���[Z ]���[Z ]���Z� \���Z�      C  , , _���Z� _���[Z `l��[Z `l��Z� _���Z�      C  , , b���Z� b���[Z cP��[Z cP��Z� b���Z�      C  , , e���Z� e���[Z f4��[Z f4��Z� e���Z�      C  , , hn��Z� hn��[Z i��[Z i��Z� hn��Z�      C  , , kR��Z� kR��[Z k���[Z k���Z� kR��Z�      C  , , n6��Z� n6��[Z n���[Z n���Z� n6��Z�      C  , , q��Z� q��[Z q���[Z q���Z� q��Z�      C  , , s���Z� s���[Z t���[Z t���Z� s���Z�      C  , , v���Z� v���[Z w���[Z w���Z� v���Z�      C  , , y���Z� y���[Z zp��[Z zp��Z� y���Z�      C  , , |���Z� |���[Z }T��[Z }T��Z� |���Z�      C  , , y���\ y���\� zp��\� zp��\ y���\      C  , , q��eF q��e� q���e� q���eF q��eF      C  , , s���eF s���e� t���e� t���eF s���eF      C  , , v���eF v���e� w���e� w���eF v���eF      C  , , y���eF y���e� zp��e� zp��eF y���eF      C  , , |���eF |���e� }T��e� }T��eF |���eF      C  , , |���\ |���\� }T��\� }T��\ |���\      C  , , i���`U i���`� j���`� j���`U i���`U      C  , , i���^9 i���^� j���^� j���^9 i���^9      C  , , l���^9 l���^� mn��^� mn��^9 l���^9      C  , , o���^9 o���^� pR��^� pR��^9 o���^9      C  , , r���^9 r���^� s6��^� s6��^9 r���^9      C  , , up��^9 up��^� v��^� v��^9 up��^9      C  , , xT��^9 xT��^� x���^� x���^9 xT��^9      C  , , {8��^9 {8��^� {���^� {���^9 {8��^9      C  , , ~��^9 ~��^� ~���^� ~���^9 ~��^9      C  , , hn��c� hn��d� i��d� i��c� hn��c�      C  , , kR��c� kR��d� k���d� k���c� kR��c�      C  , , n6��c� n6��d� n���d� n���c� n6��c�      C  , , q��c� q��d� q���d� q���c� q��c�      C  , , s���c� s���d� t���d� t���c� s���c�      C  , , v���c� v���d� w���d� w���c� v���c�      C  , , hn��f� hn��gX i��gX i��f� hn��f�      C  , , kR��f� kR��gX k���gX k���f� kR��f�      C  , , n6��f� n6��gX n���gX n���f� n6��f�      C  , , q��f� q��gX q���gX q���f� q��f�      C  , , s���f� s���gX t���gX t���f� s���f�      C  , , v���f� v���gX w���gX w���f� v���f�      C  , , y���f� y���gX zp��gX zp��f� y���f�      C  , , |���f� |���gX }T��gX }T��f� |���f�      C  , , hn��h hn��h� i��h� i��h hn��h      C  , , kR��h kR��h� k���h� k���h kR��h      C  , , n6��h n6��h� n���h� n���h n6��h      C  , , q��h q��h� q���h� q���h q��h      C  , , s���h s���h� t���h� t���h s���h      C  , , v���h v���h� w���h� w���h v���h      C  , , y���h y���h� zp��h� zp��h y���h      C  , , |���h |���h� }T��h� }T��h |���h      C  , , hn��bv hn��c  i��c  i��bv hn��bv      C  , , kR��bv kR��c  k���c  k���bv kR��bv      C  , , n6��bv n6��c  n���c  n���bv n6��bv      C  , , q��bv q��c  q���c  q���bv q��bv      C  , , s���bv s���c  t���c  t���bv s���bv      C  , , v���bv v���c  w���c  w���bv v���bv      C  , , y���bv y���c  zp��c  zp��bv y���bv      C  , , |���bv |���c  }T��c  }T��bv |���bv      C  , , y���c� y���d� zp��d� zp��c� y���c�      C  , , |���c� |���d� }T��d� }T��c� |���c�      C  , , l���`U l���`� mn��`� mn��`U l���`U      C  , , o���`U o���`� pR��`� pR��`U o���`U      C  , , r���`U r���`� s6��`� s6��`U r���`U      C  , , up��`U up��`� v��`� v��`U up��`U      C  , , xT��`U xT��`� x���`� x���`U xT��`U      C  , , {8��`U {8��`� {���`� {���`U {8��`U      C  , , ~��`U ~��`� ~���`� ~���`U ~��`U      C  , , hn��\ hn��\� i��\� i��\ hn��\      C  , , kR��\ kR��\� k���\� k���\ kR��\      C  , , n6��\ n6��\� n���\� n���\ n6��\      C  , , q��\ q��\� q���\� q���\ q��\      C  , , s���\ s���\� t���\� t���\ s���\      C  , , hn��eF hn��e� i��e� i��eF hn��eF      C  , , kR��eF kR��e� k���e� k���eF kR��eF      C  , , n6��eF n6��e� n���e� n���eF n6��eF      C  , , v���\ v���\� w���\� w���\ v���\      C  , , QN��f� QN��gX Q���gX Q���f� QN��f�      C  , , T2��f� T2��gX T���gX T���f� T2��f�      C  , , W��f� W��gX W���gX W���f� W��f�      C  , , Y���f� Y���gX Z���gX Z���f� Y���f�      C  , , \���f� \���gX ]���gX ]���f� \���f�      C  , , _���f� _���gX `l��gX `l��f� _���f�      C  , , b���f� b���gX cP��gX cP��f� b���f�      C  , , W��c� W��d� W���d� W���c� W��c�      C  , , e���f� e���gX f4��gX f4��f� e���f�      C  , , _���eF _���e� `l��e� `l��eF _���eF      C  , , b���eF b���e� cP��e� cP��eF b���eF      C  , , e���eF e���e� f4��e� f4��eF e���eF      C  , , O���^9 O���^� P���^� P���^9 O���^9      C  , , R���^9 R���^� Sj��^� Sj��^9 R���^9      C  , , U���^9 U���^� VN��^� VN��^9 U���^9      C  , , X���^9 X���^� Y2��^� Y2��^9 X���^9      C  , , [l��^9 [l��^� \��^� \��^9 [l��^9      C  , , e���h e���h� f4��h� f4��h e���h      C  , , ^P��^9 ^P��^� ^���^� ^���^9 ^P��^9      C  , , a4��^9 a4��^� a���^� a���^9 a4��^9      C  , , d��^9 d��^� d���^� d���^9 d��^9      C  , , QN��\ QN��\� Q���\� Q���\ QN��\      C  , , T2��\ T2��\� T���\� T���\ T2��\      C  , , QN��c� QN��d� Q���d� Q���c� QN��c�      C  , , W��\ W��\� W���\� W���\ W��\      C  , , Y���\ Y���\� Z���\� Z���\ Y���\      C  , , \���bv \���c  ]���c  ]���bv \���bv      C  , , _���bv _���c  `l��c  `l��bv _���bv      C  , , b���bv b���c  cP��c  cP��bv b���bv      C  , , e���bv e���c  f4��c  f4��bv e���bv      C  , , \���\ \���\� ]���\� ]���\ \���\      C  , , _���\ _���\� `l��\� `l��\ _���\      C  , , b���\ b���\� cP��\� cP��\ b���\      C  , , e���\ e���\� f4��\� f4��\ e���\      C  , , ^P��`U ^P��`� ^���`� ^���`U ^P��`U      C  , , Y���c� Y���d� Z���d� Z���c� Y���c�      C  , , a4��`U a4��`� a���`� a���`U a4��`U      C  , , d��`U d��`� d���`� d���`U d��`U      C  , , [l��`U [l��`� \��`� \��`U [l��`U      C  , , e���c� e���d� f4��d� f4��c� e���c�      C  , , QN��eF QN��e� Q���e� Q���eF QN��eF      C  , , O���`U O���`� P���`� P���`U O���`U      C  , , R���`U R���`� Sj��`� Sj��`U R���`U      C  , , U���`U U���`� VN��`� VN��`U U���`U      C  , , X���`U X���`� Y2��`� Y2��`U X���`U      C  , , T2��eF T2��e� T���e� T���eF T2��eF      C  , , W��eF W��e� W���e� W���eF W��eF      C  , , Y���eF Y���e� Z���e� Z���eF Y���eF      C  , , \���eF \���e� ]���e� ]���eF \���eF      C  , , QN��bv QN��c  Q���c  Q���bv QN��bv      C  , , T2��c� T2��d� T���d� T���c� T2��c�      C  , , T2��bv T2��c  T���c  T���bv T2��bv      C  , , W��bv W��c  W���c  W���bv W��bv      C  , , Y���bv Y���c  Z���c  Z���bv Y���bv      C  , , \���c� \���d� ]���d� ]���c� \���c�      C  , , QN��h QN��h� Q���h� Q���h QN��h      C  , , T2��h T2��h� T���h� T���h T2��h      C  , , W��h W��h� W���h� W���h W��h      C  , , Y���h Y���h� Z���h� Z���h Y���h      C  , , \���h \���h� ]���h� ]���h \���h      C  , , _���h _���h� `l��h� `l��h _���h      C  , , _���c� _���d� `l��d� `l��c� _���c�      C  , , b���h b���h� cP��h� cP��h b���h      C  , , b���c� b���d� cP��d� cP��c� b���c�      C  , , \���U \���U� ]���U� ]���U \���U      C  , , _���U _���U� `l��U� `l��U _���U      C  , , b���U b���U� cP��U� cP��U b���U      C  , , e���U e���U� f4��U� f4��U e���U      C  , , QN��YH QN��Y� Q���Y� Q���YH QN��YH      C  , , T2��YH T2��Y� T���Y� T���YH T2��YH      C  , , W��YH W��Y� W���Y� W���YH W��YH      C  , , Y���YH Y���Y� Z���Y� Z���YH Y���YH      C  , , \���YH \���Y� ]���Y� ]���YH \���YH      C  , , _���YH _���Y� `l��Y� `l��YH _���YH      C  , , b���YH b���Y� cP��Y� cP��YH b���YH      C  , , QN��W� QN��X� Q���X� Q���W� QN��W�      C  , , T2��W� T2��X� T���X� T���W� T2��W�      C  , , QN��Op QN��P Q���P Q���Op QN��Op      C  , , T2��Op T2��P T���P T���Op T2��Op      C  , , W��Op W��P W���P W���Op W��Op      C  , , Y���Op Y���P Z���P Z���Op Y���Op      C  , , \���Op \���P ]���P ]���Op \���Op      C  , , _���Op _���P `l��P `l��Op _���Op      C  , , b���Op b���P cP��P cP��Op b���Op      C  , , e���Op e���P f4��P f4��Op e���Op      C  , , e���YH e���Y� f4��Y� f4��YH e���YH      C  , , W��W� W��X� W���X� W���W� W��W�      C  , , Y���W� Y���X� Z���X� Z���W� Y���W�      C  , , \���W� \���X� ]���X� ]���W� \���W�      C  , , _���W� _���X� `l��X� `l��W� _���W�      C  , , b���W� b���X� cP��X� cP��W� b���W�      C  , , e���W� e���X� f4��X� f4��W� e���W�      C  , , QN��U QN��U� Q���U� Q���U QN��U      C  , , QN��S� QN��TR Q���TR Q���S� QN��S�      C  , , T2��S� T2��TR T���TR T���S� T2��S�      C  , , QN��P� QN��Q� Q���Q� Q���P� QN��P�      C  , , T2��P� T2��Q� T���Q� T���P� T2��P�      C  , , W��P� W��Q� W���Q� W���P� W��P�      C  , , Y���P� Y���Q� Z���Q� Z���P� Y���P�      C  , , \���P� \���Q� ]���Q� ]���P� \���P�      C  , , _���P� _���Q� `l��Q� `l��P� _���P�      C  , , b���P� b���Q� cP��Q� cP��P� b���P�      C  , , e���P� e���Q� f4��Q� f4��P� e���P�      C  , , W��S� W��TR W���TR W���S� W��S�      C  , , Y���S� Y���TR Z���TR Z���S� Y���S�      C  , , \���S� \���TR ]���TR ]���S� \���S�      C  , , _���S� _���TR `l��TR `l��S� _���S�      C  , , b���S� b���TR cP��TR cP��S� b���S�      C  , , e���S� e���TR f4��TR f4��S� e���S�      C  , , QN��R@ QN��R� Q���R� Q���R@ QN��R@      C  , , QN��N QN��N� Q���N� Q���N QN��N      C  , , T2��N T2��N� T���N� T���N T2��N      C  , , W��N W��N� W���N� W���N W��N      C  , , Y���N Y���N� Z���N� Z���N Y���N      C  , , \���N \���N� ]���N� ]���N \���N      C  , , _���N _���N� `l��N� `l��N _���N      C  , , b���N b���N� cP��N� cP��N b���N      C  , , e���N e���N� f4��N� f4��N e���N      C  , , T2��R@ T2��R� T���R� T���R@ T2��R@      C  , , W��R@ W��R� W���R� W���R@ W��R@      C  , , Y���R@ Y���R� Z���R� Z���R@ Y���R@      C  , , \���R@ \���R� ]���R� ]���R@ \���R@      C  , , _���R@ _���R� `l��R� `l��R@ _���R@      C  , , b���R@ b���R� cP��R� cP��R@ b���R@      C  , , e���R@ e���R� f4��R� f4��R@ e���R@      C  , , T2��U T2��U� T���U� T���U T2��U      C  , , QN��Vx QN��W" Q���W" Q���Vx QN��Vx      C  , , T2��Vx T2��W" T���W" T���Vx T2��Vx      C  , , W��Vx W��W" W���W" W���Vx W��Vx      C  , , Y���Vx Y���W" Z���W" Z���Vx Y���Vx      C  , , \���Vx \���W" ]���W" ]���Vx \���Vx      C  , , _���Vx _���W" `l��W" `l��Vx _���Vx      C  , , b���Vx b���W" cP��W" cP��Vx b���Vx      C  , , e���Vx e���W" f4��W" f4��Vx e���Vx      C  , , W��U W��U� W���U� W���U W��U      C  , , QN��L� QN��MJ Q���MJ Q���L� QN��L�      C  , , T2��L� T2��MJ T���MJ T���L� T2��L�      C  , , W��L� W��MJ W���MJ W���L� W��L�      C  , , Y���L� Y���MJ Z���MJ Z���L� Y���L�      C  , , \���L� \���MJ ]���MJ ]���L� \���L�      C  , , _���L� _���MJ `l��MJ `l��L� _���L�      C  , , b���L� b���MJ cP��MJ cP��L� b���L�      C  , , e���L� e���MJ f4��MJ f4��L� e���L�      C  , , Y���U Y���U� Z���U� Z���U Y���U      C  , , s���W� s���X� t���X� t���W� s���W�      C  , , v���W� v���X� w���X� w���W� v���W�      C  , , y���W� y���X� zp��X� zp��W� y���W�      C  , , |���W� |���X� }T��X� }T��W� |���W�      C  , , |���R@ |���R� }T��R� }T��R@ |���R@      C  , , kR��U kR��U� k���U� k���U kR��U      C  , , n6��U n6��U� n���U� n���U n6��U      C  , , q��U q��U� q���U� q���U q��U      C  , , s���U s���U� t���U� t���U s���U      C  , , v���U v���U� w���U� w���U v���U      C  , , y���U y���U� zp��U� zp��U y���U      C  , , |���U |���U� }T��U� }T��U |���U      C  , , hn��YH hn��Y� i��Y� i��YH hn��YH      C  , , hn��S� hn��TR i��TR i��S� hn��S�      C  , , kR��S� kR��TR k���TR k���S� kR��S�      C  , , n6��S� n6��TR n���TR n���S� n6��S�      C  , , q��S� q��TR q���TR q���S� q��S�      C  , , s���S� s���TR t���TR t���S� s���S�      C  , , v���S� v���TR w���TR w���S� v���S�      C  , , y���S� y���TR zp��TR zp��S� y���S�      C  , , |���S� |���TR }T��TR }T��S� |���S�      C  , , kR��YH kR��Y� k���Y� k���YH kR��YH      C  , , n6��YH n6��Y� n���Y� n���YH n6��YH      C  , , q��YH q��Y� q���Y� q���YH q��YH      C  , , s���YH s���Y� t���Y� t���YH s���YH      C  , , v���YH v���Y� w���Y� w���YH v���YH      C  , , y���YH y���Y� zp��Y� zp��YH y���YH      C  , , |���YH |���Y� }T��Y� }T��YH |���YH      C  , , hn��U hn��U� i��U� i��U hn��U      C  , , hn��R@ hn��R� i��R� i��R@ hn��R@      C  , , hn��N hn��N� i��N� i��N hn��N      C  , , kR��N kR��N� k���N� k���N kR��N      C  , , n6��N n6��N� n���N� n���N n6��N      C  , , q��N q��N� q���N� q���N q��N      C  , , s���N s���N� t���N� t���N s���N      C  , , v���N v���N� w���N� w���N v���N      C  , , y���N y���N� zp��N� zp��N y���N      C  , , |���N |���N� }T��N� }T��N |���N      C  , , kR��R@ kR��R� k���R� k���R@ kR��R@      C  , , hn��P� hn��Q� i��Q� i��P� hn��P�      C  , , kR��P� kR��Q� k���Q� k���P� kR��P�      C  , , n6��P� n6��Q� n���Q� n���P� n6��P�      C  , , q��P� q��Q� q���Q� q���P� q��P�      C  , , s���P� s���Q� t���Q� t���P� s���P�      C  , , v���P� v���Q� w���Q� w���P� v���P�      C  , , hn��Op hn��P i��P i��Op hn��Op      C  , , kR��Op kR��P k���P k���Op kR��Op      C  , , n6��Op n6��P n���P n���Op n6��Op      C  , , q��Op q��P q���P q���Op q��Op      C  , , s���Op s���P t���P t���Op s���Op      C  , , v���Op v���P w���P w���Op v���Op      C  , , y���Op y���P zp��P zp��Op y���Op      C  , , |���Op |���P }T��P }T��Op |���Op      C  , , y���P� y���Q� zp��Q� zp��P� y���P�      C  , , hn��Vx hn��W" i��W" i��Vx hn��Vx      C  , , kR��Vx kR��W" k���W" k���Vx kR��Vx      C  , , n6��Vx n6��W" n���W" n���Vx n6��Vx      C  , , q��Vx q��W" q���W" q���Vx q��Vx      C  , , s���Vx s���W" t���W" t���Vx s���Vx      C  , , v���Vx v���W" w���W" w���Vx v���Vx      C  , , y���Vx y���W" zp��W" zp��Vx y���Vx      C  , , |���Vx |���W" }T��W" }T��Vx |���Vx      C  , , |���P� |���Q� }T��Q� }T��P� |���P�      C  , , n6��R@ n6��R� n���R� n���R@ n6��R@      C  , , q��R@ q��R� q���R� q���R@ q��R@      C  , , s���R@ s���R� t���R� t���R@ s���R@      C  , , v���R@ v���R� w���R� w���R@ v���R@      C  , , y���R@ y���R� zp��R� zp��R@ y���R@      C  , , hn��W� hn��X� i��X� i��W� hn��W�      C  , , kR��W� kR��X� k���X� k���W� kR��W�      C  , , n6��W� n6��X� n���X� n���W� n6��W�      C  , , hn��L� hn��MJ i��MJ i��L� hn��L�      C  , , kR��L� kR��MJ k���MJ k���L� kR��L�      C  , , n6��L� n6��MJ n���MJ n���L� n6��L�      C  , , q��L� q��MJ q���MJ q���L� q��L�      C  , , s���L� s���MJ t���MJ t���L� s���L�      C  , , v���L� v���MJ w���MJ w���L� v���L�      C  , , y���L� y���MJ zp��MJ zp��L� y���L�      C  , , |���L� |���MJ }T��MJ }T��L� |���L�      C  , , q��W� q��X� q���X� q���W� q��W�      C  , , �r��i~ �r��j( ���j( ���i~ �r��i~      C  , , �V��i~ �V��j( � ��j( � ��i~ �V��i~      C  , , �:��i~ �:��j( ����j( ����i~ �:��i~      C  , , ���i~ ���j( ����j( ����i~ ���i~      C  , , ���i~ ���j( ����j( ����i~ ���i~      C  , , ����i~ ����j( ����j( ����i~ ����i~      C  , , ����i~ ����j( �t��j( �t��i~ ����i~      C  , , ����i~ ����j( �X��j( �X��i~ ����i~      C  , , ����i~ ����j( �<��j( �<��i~ ����i~      C  , , �v��i~ �v��j( � ��j( � ��i~ �v��i~      C  , , �Z��i~ �Z��j( ���j( ���i~ �Z��i~      C  , , �>��i~ �>��j( ����j( ����i~ �>��i~      C  , , �"��i~ �"��j( ����j( ����i~ �"��i~      C  , , ���i~ ���j( ����j( ����i~ ���i~      C  , , ����i~ ����j( ����j( ����i~ ����i~      C  , , ����i~ ����j( �x��j( �x��i~ ����i~      C  , , ����i~ ����j( �\��j( �\��i~ ����i~      C  , , ����i~ ����j( �@��j( �@��i~ ����i~      C  , , �z��i~ �z��j( �$��j( �$��i~ �z��i~      C  , , �^��i~ �^��j( ���j( ���i~ �^��i~      C  , , �B��i~ �B��j( ����j( ����i~ �B��i~      C  , , �&��i~ �&��j( ����j( ����i~ �&��i~      C  , , �
��i~ �
��j( ´��j( ´��i~ �
��i~      C  , , ����i~ ����j( Ř��j( Ř��i~ ����i~      C  , , ����i~ ����j( �|��j( �|��i~ ����i~      C  , , ͚��i~ ͚��j( �D��j( �D��i~ ͚��i~      C  , , ����m� ����n` �|��n` �|��m� ����m�      C  , , ͚��m� ͚��n` �D��n` �D��m� ͚��m�      C  , , �z��p� �z��q0 �$��q0 �$��p� �z��p�      C  , , �^��p� �^��q0 ���q0 ���p� �^��p�      C  , , �B��p� �B��q0 ����q0 ����p� �B��p�      C  , , �&��p� �&��q0 ����q0 ����p� �&��p�      C  , , �
��p� �
��q0 ´��q0 ´��p� �
��p�      C  , , ����p� ����q0 Ř��q0 Ř��p� ����p�      C  , , ����p� ����q0 �|��q0 �|��p� ����p�      C  , , ͚��p� ͚��q0 �D��q0 �D��p� ͚��p�      C  , , �
��q� �
��r� ´��r� ´��q� �
��q�      C  , , ����q� ����r� Ř��r� Ř��q� ����q�      C  , , ����q� ����r� �|��r� �|��q� ����q�      C  , , ͚��q� ͚��r� �D��r� �D��q� ͚��q�      C  , , ����j� ����k� �\��k� �\��j� ����j�      C  , , ����j� ����k� �@��k� �@��j� ����j�      C  , , �z��j� �z��k� �$��k� �$��j� �z��j�      C  , , �^��j� �^��k� ���k� ���j� �^��j�      C  , , �B��j� �B��k� ����k� ����j� �B��j�      C  , , �&��j� �&��k� ����k� ����j� �&��j�      C  , , �
��j� �
��k� ´��k� ´��j� �
��j�      C  , , ����j� ����k� Ř��k� Ř��j� ����j�      C  , , ����j� ����k� �|��k� �|��j� ����j�      C  , , ͚��j� ͚��k� �D��k� �D��j� ͚��j�      C  , , ����o ����o� �\��o� �\��o ����o      C  , , ����o ����o� �@��o� �@��o ����o      C  , , �&��lN �&��l� ����l� ����lN �&��lN      C  , , �
��lN �
��l� ´��l� ´��lN �
��lN      C  , , ����lN ����l� Ř��l� Ř��lN ����lN      C  , , ����lN ����l� �|��l� �|��lN ����lN      C  , , ͚��lN ͚��l� �D��l� �D��lN ͚��lN      C  , , ����q� ����r� �\��r� �\��q� ����q�      C  , , ����q� ����r� �@��r� �@��q� ����q�      C  , , ����lN ����l� �\��l� �\��lN ����lN      C  , , �^��lN �^��l� ���l� ���lN �^��lN      C  , , �B��lN �B��l� ����l� ����lN �B��lN      C  , , �z��o �z��o� �$��o� �$��o �z��o      C  , , �^��o �^��o� ���o� ���o �^��o      C  , , �B��o �B��o� ����o� ����o �B��o      C  , , �&��o �&��o� ����o� ����o �&��o      C  , , �
��o �
��o� ´��o� ´��o �
��o      C  , , ����o ����o� Ř��o� Ř��o ����o      C  , , ����o ����o� �|��o� �|��o ����o      C  , , ͚��o ͚��o� �D��o� �D��o ͚��o      C  , , �z��q� �z��r� �$��r� �$��q� �z��q�      C  , , �^��q� �^��r� ���r� ���q� �^��q�      C  , , �B��q� �B��r� ����r� ����q� �B��q�      C  , , �&��q� �&��r� ����r� ����q� �&��q�      C  , , ����lN ����l� �@��l� �@��lN ����lN      C  , , �z��lN �z��l� �$��l� �$��lN �z��lN      C  , , ����m� ����n` �\��n` �\��m� ����m�      C  , , ����m� ����n` �@��n` �@��m� ����m�      C  , , �z��m� �z��n` �$��n` �$��m� �z��m�      C  , , �^��m� �^��n` ���n` ���m� �^��m�      C  , , �B��m� �B��n` ����n` ����m� �B��m�      C  , , �&��m� �&��n` ����n` ����m� �&��m�      C  , , �
��m� �
��n` ´��n` ´��m� �
��m�      C  , , ����m� ����n` Ř��n` Ř��m� ����m�      C  , , ����p� ����q0 �\��q0 �\��p� ����p�      C  , , ����p� ����q0 �@��q0 �@��p� ����p�      C  , , �>��lN �>��l� ����l� ����lN �>��lN      C  , , �"��lN �"��l� ����l� ����lN �"��lN      C  , , ���lN ���l� ����l� ����lN ���lN      C  , , ����lN ����l� ����l� ����lN ����lN      C  , , ����lN ����l� �x��l� �x��lN ����lN      C  , , �r��q� �r��r� ���r� ���q� �r��q�      C  , , �V��q� �V��r� � ��r� � ��q� �V��q�      C  , , �:��q� �:��r� ����r� ����q� �:��q�      C  , , ���q� ���r� ����r� ����q� ���q�      C  , , ����q� ����r� �X��r� �X��q� ����q�      C  , , ����q� ����r� �<��r� �<��q� ����q�      C  , , �r��m� �r��n` ���n` ���m� �r��m�      C  , , �v��q� �v��r� � ��r� � ��q� �v��q�      C  , , �V��m� �V��n` � ��n` � ��m� �V��m�      C  , , �:��m� �:��n` ����n` ����m� �:��m�      C  , , ���m� ���n` ����n` ����m� ���m�      C  , , ���m� ���n` ����n` ����m� ���m�      C  , , ����m� ����n` ����n` ����m� ����m�      C  , , ����m� ����n` �t��n` �t��m� ����m�      C  , , �>��j� �>��k� ����k� ����j� �>��j�      C  , , �"��j� �"��k� ����k� ����j� �"��j�      C  , , ���j� ���k� ����k� ����j� ���j�      C  , , ����j� ����k� ����k� ����j� ����j�      C  , , ����j� ����k� �x��k� �x��j� ����j�      C  , , ����m� ����n` �X��n` �X��m� ����m�      C  , , ����m� ����n` �<��n` �<��m� ����m�      C  , , �v��m� �v��n` � ��n` � ��m� �v��m�      C  , , �>��o �>��o� ����o� ����o �>��o      C  , , �"��o �"��o� ����o� ����o �"��o      C  , , ���o ���o� ����o� ����o ���o      C  , , �r��p� �r��q0 ���q0 ���p� �r��p�      C  , , �V��p� �V��q0 � ��q0 � ��p� �V��p�      C  , , �:��p� �:��q0 ����q0 ����p� �:��p�      C  , , ���p� ���q0 ����q0 ����p� ���p�      C  , , ����o ����o� ����o� ����o ����o      C  , , ����o ����o� �x��o� �x��o ����o      C  , , ���p� ���q0 ����q0 ����p� ���p�      C  , , ����p� ����q0 ����q0 ����p� ����p�      C  , , �r��o �r��o� ���o� ���o �r��o      C  , , �V��o �V��o� � ��o� � ��o �V��o      C  , , �:��o �:��o� ����o� ����o �:��o      C  , , ���o ���o� ����o� ����o ���o      C  , , ���o ���o� ����o� ����o ���o      C  , , �Z��q� �Z��r� ���r� ���q� �Z��q�      C  , , �>��q� �>��r� ����r� ����q� �>��q�      C  , , �"��q� �"��r� ����r� ����q� �"��q�      C  , , ���q� ���r� ����r� ����q� ���q�      C  , , ����q� ����r� ����r� ����q� ����q�      C  , , ����q� ����r� �x��r� �x��q� ����q�      C  , , ����o ����o� ����o� ����o ����o      C  , , ����o ����o� �t��o� �t��o ����o      C  , , ����o ����o� �X��o� �X��o ����o      C  , , ����o ����o� �<��o� �<��o ����o      C  , , �v��o �v��o� � ��o� � ��o �v��o      C  , , �Z��o �Z��o� ���o� ���o �Z��o      C  , , �r��j� �r��k� ���k� ���j� �r��j�      C  , , �V��j� �V��k� � ��k� � ��j� �V��j�      C  , , �:��j� �:��k� ����k� ����j� �:��j�      C  , , ���j� ���k� ����k� ����j� ���j�      C  , , ���j� ���k� ����k� ����j� ���j�      C  , , ����j� ����k� ����k� ����j� ����j�      C  , , ����j� ����k� �t��k� �t��j� ����j�      C  , , ����j� ����k� �X��k� �X��j� ����j�      C  , , �r��lN �r��l� ���l� ���lN �r��lN      C  , , �V��lN �V��l� � ��l� � ��lN �V��lN      C  , , �:��lN �:��l� ����l� ����lN �:��lN      C  , , ���lN ���l� ����l� ����lN ���lN      C  , , ���lN ���l� ����l� ����lN ���lN      C  , , ����lN ����l� ����l� ����lN ����lN      C  , , ����lN ����l� �t��l� �t��lN ����lN      C  , , ����lN ����l� �X��l� �X��lN ����lN      C  , , ����j� ����k� �<��k� �<��j� ����j�      C  , , �v��j� �v��k� � ��k� � ��j� �v��j�      C  , , ���q� ���r� ����r� ����q� ���q�      C  , , ����q� ����r� ����r� ����q� ����q�      C  , , �Z��j� �Z��k� ���k� ���j� �Z��j�      C  , , �Z��m� �Z��n` ���n` ���m� �Z��m�      C  , , �>��m� �>��n` ����n` ����m� �>��m�      C  , , �"��m� �"��n` ����n` ����m� �"��m�      C  , , ���m� ���n` ����n` ����m� ���m�      C  , , ����m� ����n` ����n` ����m� ����m�      C  , , ����m� ����n` �x��n` �x��m� ����m�      C  , , ����q� ����r� �t��r� �t��q� ����q�      C  , , ����lN ����l� �<��l� �<��lN ����lN      C  , , ����p� ����q0 �t��q0 �t��p� ����p�      C  , , ����p� ����q0 �X��q0 �X��p� ����p�      C  , , ����p� ����q0 �<��q0 �<��p� ����p�      C  , , �v��p� �v��q0 � ��q0 � ��p� �v��p�      C  , , �Z��p� �Z��q0 ���q0 ���p� �Z��p�      C  , , �>��p� �>��q0 ����q0 ����p� �>��p�      C  , , �"��p� �"��q0 ����q0 ����p� �"��p�      C  , , ���p� ���q0 ����q0 ����p� ���p�      C  , , ����p� ����q0 ����q0 ����p� ����p�      C  , , ����p� ����q0 �x��q0 �x��p� ����p�      C  , , �v��lN �v��l� � ��l� � ��lN �v��lN      C  , , �Z��lN �Z��l� ���l� ���lN �Z��lN      C  , , �r��Z� �r��[Z ���[Z ���Z� �r��Z�      C  , , �V��Z� �V��[Z � ��[Z � ��Z� �V��Z�      C  , , �:��Z� �:��[Z ����[Z ����Z� �:��Z�      C  , , ���Z� ���[Z ����[Z ����Z� ���Z�      C  , , ���Z� ���[Z ����[Z ����Z� ���Z�      C  , , ����Z� ����[Z ����[Z ����Z� ����Z�      C  , , ����Z� ����[Z �t��[Z �t��Z� ����Z�      C  , , ����Z� ����[Z �X��[Z �X��Z� ����Z�      C  , , ����Z� ����[Z �<��[Z �<��Z� ����Z�      C  , , �v��Z� �v��[Z � ��[Z � ��Z� �v��Z�      C  , , �Z��Z� �Z��[Z ���[Z ���Z� �Z��Z�      C  , , �>��Z� �>��[Z ����[Z ����Z� �>��Z�      C  , , �"��Z� �"��[Z ����[Z ����Z� �"��Z�      C  , , ���Z� ���[Z ����[Z ����Z� ���Z�      C  , , ����Z� ����[Z ����[Z ����Z� ����Z�      C  , , ����Z� ����[Z �x��[Z �x��Z� ����Z�      C  , , � ��`U � ��`� ����`� ����`U � ��`U      C  , , � ��^9 � ��^� ����^� ����^9 � ��^9      C  , , ����f� ����gX ����gX ����f� ����f�      C  , , ����f� ����gX �x��gX �x��f� ����f�      C  , , �x��`U �x��`� �"��`� �"��`U �x��`U      C  , , �\��`U �\��`� ���`� ���`U �\��`U      C  , , �@��`U �@��`� ����`� ����`U �@��`U      C  , , �v��f� �v��gX � ��gX � ��f� �v��f�      C  , , �Z��f� �Z��gX ���gX ���f� �Z��f�      C  , , �>��f� �>��gX ����gX ����f� �>��f�      C  , , �"��f� �"��gX ����gX ����f� �"��f�      C  , , ����eF ����e� �<��e� �<��eF ����eF      C  , , �Z��h �Z��h� ���h� ���h �Z��h      C  , , �>��h �>��h� ����h� ����h �>��h      C  , , ���h ���h� ����h� ����h ���h      C  , , �v��eF �v��e� � ��e� � ��eF �v��eF      C  , , �Z��eF �Z��e� ���e� ���eF �Z��eF      C  , , �>��eF �>��e� ����e� ����eF �>��eF      C  , , �"��eF �"��e� ����e� ����eF �"��eF      C  , , ���eF ���e� ����e� ����eF ���eF      C  , , ����eF ����e� ����e� ����eF ����eF      C  , , ����eF ����e� �x��e� �x��eF ����eF      C  , , ����h ����h� ����h� ����h ����h      C  , , ����h ����h� �x��h� �x��h ����h      C  , , ����bv ����c  �<��c  �<��bv ����bv      C  , , �v��bv �v��c  � ��c  � ��bv �v��bv      C  , , �Z��bv �Z��c  ���c  ���bv �Z��bv      C  , , �>��bv �>��c  ����c  ����bv �>��bv      C  , , �"��bv �"��c  ����c  ����bv �"��bv      C  , , �"��h �"��h� ����h� ����h �"��h      C  , , ����\ ����\� �<��\� �<��\ ����\      C  , , �v��\ �v��\� � ��\� � ��\ �v��\      C  , , �Z��\ �Z��\� ���\� ���\ �Z��\      C  , , �>��\ �>��\� ����\� ����\ �>��\      C  , , �"��\ �"��\� ����\� ����\ �"��\      C  , , ���\ ���\� ����\� ����\ ���\      C  , , ����\ ����\� ����\� ����\ ����\      C  , , ����\ ����\� �x��\� �x��\ ����\      C  , , ���bv ���c  ����c  ����bv ���bv      C  , , ���`U ���`� ����`� ����`U ���`U      C  , , ����`U ����`� ����`� ����`U ����`U      C  , , ����`U ����`� �v��`� �v��`U ����`U      C  , , ����`U ����`� �Z��`� �Z��`U ����`U      C  , , ����`U ����`� �>��`� �>��`U ����`U      C  , , ����bv ����c  ����c  ����bv ����bv      C  , , ����bv ����c  �x��c  �x��bv ����bv      C  , , ���f� ���gX ����gX ����f� ���f�      C  , , ���^9 ���^� ����^� ����^9 ���^9      C  , , ����^9 ����^� ����^� ����^9 ����^9      C  , , ����^9 ����^� �v��^� �v��^9 ����^9      C  , , ����^9 ����^� �Z��^� �Z��^9 ����^9      C  , , ����^9 ����^� �>��^� �>��^9 ����^9      C  , , �x��^9 �x��^� �"��^� �"��^9 �x��^9      C  , , �\��^9 �\��^� ���^� ���^9 �\��^9      C  , , �@��^9 �@��^� ����^� ����^9 �@��^9      C  , , ����c� ����d� �<��d� �<��c� ����c�      C  , , �v��c� �v��d� � ��d� � ��c� �v��c�      C  , , �Z��c� �Z��d� ���d� ���c� �Z��c�      C  , , �>��c� �>��d� ����d� ����c� �>��c�      C  , , �"��c� �"��d� ����d� ����c� �"��c�      C  , , ���c� ���d� ����d� ����c� ���c�      C  , , ����c� ����d� ����d� ����c� ����c�      C  , , ����c� ����d� �x��d� �x��c� ����c�      C  , , ����h ����h� �<��h� �<��h ����h      C  , , �v��h �v��h� � ��h� � ��h �v��h      C  , , ����f� ����gX �<��gX �<��f� ����f�      C  , , �:��bv �:��c  ����c  ����bv �:��bv      C  , , ���bv ���c  ����c  ����bv ���bv      C  , , ���bv ���c  ����c  ����bv ���bv      C  , , � ��`U � ��`� ����`� ����`U � ��`U      C  , , ����`U ����`� ����`� ����`U ����`U      C  , , ����`U ����`� �r��`� �r��`U ����`U      C  , , ����`U ����`� �V��`� �V��`U ����`U      C  , , �V��c� �V��d� � ��d� � ��c� �V��c�      C  , , �:��c� �:��d� ����d� ����c� �:��c�      C  , , �r��bv �r��c  ���c  ���bv �r��bv      C  , , �r��eF �r��e� ���e� ���eF �r��eF      C  , , �V��eF �V��e� � ��e� � ��eF �V��eF      C  , , �:��eF �:��e� ����e� ����eF �:��eF      C  , , ����`U ����`� �:��`� �:��`U ����`U      C  , , �t��`U �t��`� ���`� ���`U �t��`U      C  , , ���c� ���d� ����d� ����c� ���c�      C  , , � ��^9 � ��^� ����^� ����^9 � ��^9      C  , , ����^9 ����^� ����^� ����^9 ����^9      C  , , ����^9 ����^� �r��^� �r��^9 ����^9      C  , , ����^9 ����^� �V��^� �V��^9 ����^9      C  , , ����^9 ����^� �:��^� �:��^9 ����^9      C  , , �t��^9 �t��^� ���^� ���^9 �t��^9      C  , , �X��^9 �X��^� ���^� ���^9 �X��^9      C  , , �<��^9 �<��^� ����^� ����^9 �<��^9      C  , , �X��`U �X��`� ���`� ���`U �X��`U      C  , , ����bv ����c  ����c  ����bv ����bv      C  , , ����bv ����c  �t��c  �t��bv ����bv      C  , , ����bv ����c  �X��c  �X��bv ����bv      C  , , ���eF ���e� ����e� ����eF ���eF      C  , , ���eF ���e� ����e� ����eF ���eF      C  , , ����eF ����e� ����e� ����eF ����eF      C  , , ����eF ����e� �t��e� �t��eF ����eF      C  , , ����eF ����e� �X��e� �X��eF ����eF      C  , , ���c� ���d� ����d� ����c� ���c�      C  , , ����c� ����d� ����d� ����c� ����c�      C  , , ����c� ����d� �t��d� �t��c� ����c�      C  , , ����c� ����d� �X��d� �X��c� ����c�      C  , , �r��\ �r��\� ���\� ���\ �r��\      C  , , �V��\ �V��\� � ��\� � ��\ �V��\      C  , , �:��\ �:��\� ����\� ����\ �:��\      C  , , ���\ ���\� ����\� ����\ ���\      C  , , ���\ ���\� ����\� ����\ ���\      C  , , ����\ ����\� ����\� ����\ ����\      C  , , ����\ ����\� �t��\� �t��\ ����\      C  , , �<��`U �<��`� ����`� ����`U �<��`U      C  , , �r��h �r��h� ���h� ���h �r��h      C  , , �V��h �V��h� � ��h� � ��h �V��h      C  , , �:��h �:��h� ����h� ����h �:��h      C  , , ���h ���h� ����h� ����h ���h      C  , , ���h ���h� ����h� ����h ���h      C  , , ����h ����h� ����h� ����h ����h      C  , , ����h ����h� �t��h� �t��h ����h      C  , , ����h ����h� �X��h� �X��h ����h      C  , , �r��c� �r��d� ���d� ���c� �r��c�      C  , , ����\ ����\� �X��\� �X��\ ����\      C  , , �r��f� �r��gX ���gX ���f� �r��f�      C  , , �V��f� �V��gX � ��gX � ��f� �V��f�      C  , , �:��f� �:��gX ����gX ����f� �:��f�      C  , , ���f� ���gX ����gX ����f� ���f�      C  , , ���f� ���gX ����gX ����f� ���f�      C  , , ����f� ����gX ����gX ����f� ����f�      C  , , ����f� ����gX �t��gX �t��f� ����f�      C  , , ����f� ����gX �X��gX �X��f� ����f�      C  , , �V��bv �V��c  � ��c  � ��bv �V��bv      C  , , �V��Op �V��P � ��P � ��Op �V��Op      C  , , �:��Op �:��P ����P ����Op �:��Op      C  , , ���Op ���P ����P ����Op ���Op      C  , , ���Op ���P ����P ����Op ���Op      C  , , ����Op ����P ����P ����Op ����Op      C  , , ����Op ����P �t��P �t��Op ����Op      C  , , ����Op ����P �X��P �X��Op ����Op      C  , , ����P� ����Q� �X��Q� �X��P� ����P�      C  , , ���Vx ���W" ����W" ����Vx ���Vx      C  , , ����Vx ����W" ����W" ����Vx ����Vx      C  , , ����Vx ����W" �t��W" �t��Vx ����Vx      C  , , ����Vx ����W" �X��W" �X��Vx ����Vx      C  , , ���R@ ���R� ����R� ����R@ ���R@      C  , , ���R@ ���R� ����R� ����R@ ���R@      C  , , ����R@ ����R� ����R� ����R@ ����R@      C  , , ����R@ ����R� �t��R� �t��R@ ����R@      C  , , ����R@ ����R� �X��R� �X��R@ ����R@      C  , , �r��YH �r��Y� ���Y� ���YH �r��YH      C  , , �V��YH �V��Y� � ��Y� � ��YH �V��YH      C  , , �:��YH �:��Y� ����Y� ����YH �:��YH      C  , , ���YH ���Y� ����Y� ����YH ���YH      C  , , ���YH ���Y� ����Y� ����YH ���YH      C  , , ����YH ����Y� ����Y� ����YH ����YH      C  , , ����YH ����Y� �t��Y� �t��YH ����YH      C  , , ����YH ����Y� �X��Y� �X��YH ����YH      C  , , ����S� ����TR �X��TR �X��S� ����S�      C  , , �r��S� �r��TR ���TR ���S� �r��S�      C  , , �r��U �r��U� ���U� ���U �r��U      C  , , �V��U �V��U� � ��U� � ��U �V��U      C  , , �r��N �r��N� ���N� ���N �r��N      C  , , �V��N �V��N� � ��N� � ��N �V��N      C  , , �:��N �:��N� ����N� ����N �:��N      C  , , ���N ���N� ����N� ����N ���N      C  , , ���N ���N� ����N� ����N ���N      C  , , ����N ����N� ����N� ����N ����N      C  , , ����N ����N� �t��N� �t��N ����N      C  , , ����N ����N� �X��N� �X��N ����N      C  , , �:��U �:��U� ����U� ����U �:��U      C  , , ���U ���U� ����U� ����U ���U      C  , , ���U ���U� ����U� ����U ���U      C  , , ����U ����U� ����U� ����U ����U      C  , , ����U ����U� �t��U� �t��U ����U      C  , , ����U ����U� �X��U� �X��U ����U      C  , , �V��S� �V��TR � ��TR � ��S� �V��S�      C  , , �:��S� �:��TR ����TR ����S� �:��S�      C  , , ���S� ���TR ����TR ����S� ���S�      C  , , ���S� ���TR ����TR ����S� ���S�      C  , , ����S� ����TR ����TR ����S� ����S�      C  , , ����S� ����TR �t��TR �t��S� ����S�      C  , , �r��R@ �r��R� ���R� ���R@ �r��R@      C  , , �V��R@ �V��R� � ��R� � ��R@ �V��R@      C  , , �:��R@ �:��R� ����R� ����R@ �:��R@      C  , , �r��Vx �r��W" ���W" ���Vx �r��Vx      C  , , �r��W� �r��X� ���X� ���W� �r��W�      C  , , �V��W� �V��X� � ��X� � ��W� �V��W�      C  , , �:��W� �:��X� ����X� ����W� �:��W�      C  , , ���W� ���X� ����X� ����W� ���W�      C  , , ���W� ���X� ����X� ����W� ���W�      C  , , �V��Vx �V��W" � ��W" � ��Vx �V��Vx      C  , , �:��Vx �:��W" ����W" ����Vx �:��Vx      C  , , ����W� ����X� ����X� ����W� ����W�      C  , , ����W� ����X� �t��X� �t��W� ����W�      C  , , ����W� ����X� �X��X� �X��W� ����W�      C  , , ���Vx ���W" ����W" ����Vx ���Vx      C  , , �r��P� �r��Q� ���Q� ���P� �r��P�      C  , , �V��P� �V��Q� � ��Q� � ��P� �V��P�      C  , , �:��P� �:��Q� ����Q� ����P� �:��P�      C  , , ���P� ���Q� ����Q� ����P� ���P�      C  , , ���P� ���Q� ����Q� ����P� ���P�      C  , , ����P� ����Q� ����Q� ����P� ����P�      C  , , ����P� ����Q� �t��Q� �t��P� ����P�      C  , , �r��Op �r��P ���P ���Op �r��Op      C  , , �r��L� �r��MJ ���MJ ���L� �r��L�      C  , , �V��L� �V��MJ � ��MJ � ��L� �V��L�      C  , , �:��L� �:��MJ ����MJ ����L� �:��L�      C  , , ���L� ���MJ ����MJ ����L� ���L�      C  , , ���L� ���MJ ����MJ ����L� ���L�      C  , , ����L� ����MJ ����MJ ����L� ����L�      C  , , ����L� ����MJ �t��MJ �t��L� ����L�      C  , , ����L� ����MJ �X��MJ �X��L� ����L�      C  , , ����Vx ����W" ����W" ����Vx ����Vx      C  , , ����Vx ����W" �x��W" �x��Vx ����Vx      C  , , �Z��S� �Z��TR ���TR ���S� �Z��S�      C  , , �>��S� �>��TR ����TR ����S� �>��S�      C  , , �"��S� �"��TR ����TR ����S� �"��S�      C  , , ����R@ ����R� �<��R� �<��R@ ����R@      C  , , �v��R@ �v��R� � ��R� � ��R@ �v��R@      C  , , ����N ����N� �<��N� �<��N ����N      C  , , �v��N �v��N� � ��N� � ��N �v��N      C  , , �Z��N �Z��N� ���N� ���N �Z��N      C  , , �>��N �>��N� ����N� ����N �>��N      C  , , �"��N �"��N� ����N� ����N �"��N      C  , , ���N ���N� ����N� ����N ���N      C  , , ����N ����N� ����N� ����N ����N      C  , , ����N ����N� �x��N� �x��N ����N      C  , , �Z��R@ �Z��R� ���R� ���R@ �Z��R@      C  , , �>��R@ �>��R� ����R� ����R@ �>��R@      C  , , �"��R@ �"��R� ����R� ����R@ �"��R@      C  , , ���R@ ���R� ����R� ����R@ ���R@      C  , , ����Op ����P �<��P �<��Op ����Op      C  , , �v��Op �v��P � ��P � ��Op �v��Op      C  , , ����U ����U� �<��U� �<��U ����U      C  , , �v��U �v��U� � ��U� � ��U �v��U      C  , , �Z��U �Z��U� ���U� ���U �Z��U      C  , , �>��U �>��U� ����U� ����U �>��U      C  , , �"��U �"��U� ����U� ����U �"��U      C  , , ���U ���U� ����U� ����U ���U      C  , , ����U ����U� ����U� ����U ����U      C  , , ����U ����U� �x��U� �x��U ����U      C  , , �Z��Op �Z��P ���P ���Op �Z��Op      C  , , �>��Op �>��P ����P ����Op �>��Op      C  , , �"��Op �"��P ����P ����Op �"��Op      C  , , ���Op ���P ����P ����Op ���Op      C  , , ����Op ����P ����P ����Op ����Op      C  , , ����Op ����P �x��P �x��Op ����Op      C  , , ����R@ ����R� ����R� ����R@ ����R@      C  , , ����W� ����X� �<��X� �<��W� ����W�      C  , , �v��W� �v��X� � ��X� � ��W� �v��W�      C  , , �Z��W� �Z��X� ���X� ���W� �Z��W�      C  , , �>��W� �>��X� ����X� ����W� �>��W�      C  , , �"��W� �"��X� ����X� ����W� �"��W�      C  , , ���W� ���X� ����X� ����W� ���W�      C  , , ����R@ ����R� �x��R� �x��R@ ����R@      C  , , ���S� ���TR ����TR ����S� ���S�      C  , , ����S� ����TR ����TR ����S� ����S�      C  , , ����S� ����TR �x��TR �x��S� ����S�      C  , , ����P� ����Q� �<��Q� �<��P� ����P�      C  , , �v��P� �v��Q� � ��Q� � ��P� �v��P�      C  , , �Z��P� �Z��Q� ���Q� ���P� �Z��P�      C  , , �>��P� �>��Q� ����Q� ����P� �>��P�      C  , , �"��P� �"��Q� ����Q� ����P� �"��P�      C  , , ���P� ���Q� ����Q� ����P� ���P�      C  , , ����P� ����Q� ����Q� ����P� ����P�      C  , , ����P� ����Q� �x��Q� �x��P� ����P�      C  , , ����W� ����X� �x��X� �x��W� ����W�      C  , , ����W� ����X� ����X� ����W� ����W�      C  , , ����S� ����TR �<��TR �<��S� ����S�      C  , , �v��S� �v��TR � ��TR � ��S� �v��S�      C  , , ����Vx ����W" �<��W" �<��Vx ����Vx      C  , , ����YH ����Y� �<��Y� �<��YH ����YH      C  , , �v��YH �v��Y� � ��Y� � ��YH �v��YH      C  , , �Z��YH �Z��Y� ���Y� ���YH �Z��YH      C  , , �>��YH �>��Y� ����Y� ����YH �>��YH      C  , , �"��YH �"��Y� ����Y� ����YH �"��YH      C  , , ���YH ���Y� ����Y� ����YH ���YH      C  , , ����YH ����Y� ����Y� ����YH ����YH      C  , , ����YH ����Y� �x��Y� �x��YH ����YH      C  , , �v��Vx �v��W" � ��W" � ��Vx �v��Vx      C  , , �Z��Vx �Z��W" ���W" ���Vx �Z��Vx      C  , , �>��Vx �>��W" ����W" ����Vx �>��Vx      C  , , �"��Vx �"��W" ����W" ����Vx �"��Vx      C  , , ���Vx ���W" ����W" ����Vx ���Vx      C  , , ����L� ����MJ �<��MJ �<��L� ����L�      C  , , �v��L� �v��MJ � ��MJ � ��L� �v��L�      C  , , �Z��L� �Z��MJ ���MJ ���L� �Z��L�      C  , , �>��L� �>��MJ ����MJ ����L� �>��L�      C  , , �"��L� �"��MJ ����MJ ����L� �"��L�      C  , , ���L� ���MJ ����MJ ����L� ���L�      C  , , ����L� ����MJ ����MJ ����L� ����L�      C  , , ����L� ����MJ �x��MJ �x��L� ����L�      C  , , ����Z� ����[Z �\��[Z �\��Z� ����Z�      C  , , ����Z� ����[Z �@��[Z �@��Z� ����Z�      C  , , �z��Z� �z��[Z �$��[Z �$��Z� �z��Z�      C  , , �^��Z� �^��[Z ���[Z ���Z� �^��Z�      C  , , �B��Z� �B��[Z ����[Z ����Z� �B��Z�      C  , , �&��Z� �&��[Z ����[Z ����Z� �&��Z�      C  , , �
��Z� �
��[Z ´��[Z ´��Z� �
��Z�      C  , , ����Z� ����[Z Ř��[Z Ř��Z� ����Z�      C  , , ����Z� ����[Z �|��[Z �|��Z� ����Z�      C  , , �D��^9 �D��^� ����^� ����^9 �D��^9      C  , , �(��^9 �(��^� ����^� ����^9 �(��^9      C  , , ͚��c� ͚��d� �D��d� �D��c� ͚��c�      C  , , ͚��eF ͚��e� �D��e� �D��eF ͚��eF      C  , , �D��`U �D��`� ����`� ����`U �D��`U      C  , , �(��`U �(��`� ����`� ����`U �(��`U      C  , , ͚��f� ͚��gX �D��gX �D��f� ͚��f�      C  , , ͚��h ͚��h� �D��h� �D��h ͚��h      C  , , ͚��bv ͚��c  �D��c  �D��bv ͚��bv      C  , , �^��h �^��h� ���h� ���h �^��h      C  , , �B��h �B��h� ����h� ����h �B��h      C  , , �&��h �&��h� ����h� ����h �&��h      C  , , �
��h �
��h� ´��h� ´��h �
��h      C  , , ����h ����h� Ř��h� Ř��h ����h      C  , , ����h ����h� �|��h� �|��h ����h      C  , , �$��`U �$��`� ����`� ����`U �$��`U      C  , , ����`U ����`� ����`� ����`U ����`U      C  , , ���^9 ���^� ����^� ����^9 ���^9      C  , , ����^9 ����^� ����^� ����^9 ����^9      C  , , ����^9 ����^� �z��^� �z��^9 ����^9      C  , , ����^9 ����^� �^��^� �^��^9 ����^9      C  , , ����^9 ����^� �B��^� �B��^9 ����^9      C  , , �|��^9 �|��^� �&��^� �&��^9 �|��^9      C  , , �`��^9 �`��^� �
��^� �
��^9 �`��^9      C  , , ���`U ���`� ����`� ����`U ���`U      C  , , �&��c� �&��d� ����d� ����c� �&��c�      C  , , �
��c� �
��d� ´��d� ´��c� �
��c�      C  , , ����f� ����gX �\��gX �\��f� ����f�      C  , , ����`U ����`� �z��`� �z��`U ����`U      C  , , ����`U ����`� �^��`� �^��`U ����`U      C  , , ����`U ����`� �B��`� �B��`U ����`U      C  , , ����\ ����\� �\��\� �\��\ ����\      C  , , ����\ ����\� �@��\� �@��\ ����\      C  , , �z��\ �z��\� �$��\� �$��\ �z��\      C  , , �^��\ �^��\� ���\� ���\ �^��\      C  , , ����eF ����e� �|��e� �|��eF ����eF      C  , , ����c� ����d� Ř��d� Ř��c� ����c�      C  , , �B��\ �B��\� ����\� ����\ �B��\      C  , , �&��\ �&��\� ����\� ����\ �&��\      C  , , �
��\ �
��\� ´��\� ´��\ �
��\      C  , , ����\ ����\� Ř��\� Ř��\ ����\      C  , , ����\ ����\� �|��\� �|��\ ����\      C  , , �|��`U �|��`� �&��`� �&��`U �|��`U      C  , , �`��`U �`��`� �
��`� �
��`U �`��`U      C  , , ����c� ����d� �|��d� �|��c� ����c�      C  , , ����eF ����e� �\��e� �\��eF ����eF      C  , , ����f� ����gX �@��gX �@��f� ����f�      C  , , �z��f� �z��gX �$��gX �$��f� �z��f�      C  , , �^��f� �^��gX ���gX ���f� �^��f�      C  , , �B��f� �B��gX ����gX ����f� �B��f�      C  , , �&��f� �&��gX ����gX ����f� �&��f�      C  , , �
��f� �
��gX ´��gX ´��f� �
��f�      C  , , ����f� ����gX Ř��gX Ř��f� ����f�      C  , , ����f� ����gX �|��gX �|��f� ����f�      C  , , ����eF ����e� �@��e� �@��eF ����eF      C  , , ����bv ����c  �\��c  �\��bv ����bv      C  , , ����bv ����c  �@��c  �@��bv ����bv      C  , , �z��bv �z��c  �$��c  �$��bv �z��bv      C  , , �z��eF �z��e� �$��e� �$��eF �z��eF      C  , , �^��eF �^��e� ���e� ���eF �^��eF      C  , , �B��eF �B��e� ����e� ����eF �B��eF      C  , , �&��eF �&��e� ����e� ����eF �&��eF      C  , , �
��eF �
��e� ´��e� ´��eF �
��eF      C  , , ����eF ����e� Ř��e� Ř��eF ����eF      C  , , �$��^9 �$��^� ����^� ����^9 �$��^9      C  , , ����h ����h� �\��h� �\��h ����h      C  , , ����h ����h� �@��h� �@��h ����h      C  , , �^��bv �^��c  ���c  ���bv �^��bv      C  , , ����c� ����d� �\��d� �\��c� ����c�      C  , , ����c� ����d� �@��d� �@��c� ����c�      C  , , �z��c� �z��d� �$��d� �$��c� �z��c�      C  , , �^��c� �^��d� ���d� ���c� �^��c�      C  , , �B��c� �B��d� ����d� ����c� �B��c�      C  , , �B��bv �B��c  ����c  ����bv �B��bv      C  , , �&��bv �&��c  ����c  ����bv �&��bv      C  , , �
��bv �
��c  ´��c  ´��bv �
��bv      C  , , ����bv ����c  Ř��c  Ř��bv ����bv      C  , , ����bv ����c  �|��c  �|��bv ����bv      C  , , �z��h �z��h� �$��h� �$��h �z��h      C  , , ����S� ����TR �|��TR �|��S� ����S�      C  , , �
��R@ �
��R� ´��R� ´��R@ �
��R@      C  , , ����R@ ����R� Ř��R� Ř��R@ ����R@      C  , , ����U ����U� �\��U� �\��U ����U      C  , , ����U ����U� �@��U� �@��U ����U      C  , , �z��U �z��U� �$��U� �$��U �z��U      C  , , �^��U �^��U� ���U� ���U �^��U      C  , , ����N ����N� �\��N� �\��N ����N      C  , , ����N ����N� �@��N� �@��N ����N      C  , , �z��N �z��N� �$��N� �$��N �z��N      C  , , �^��N �^��N� ���N� ���N �^��N      C  , , �B��N �B��N� ����N� ����N �B��N      C  , , �&��N �&��N� ����N� ����N �&��N      C  , , �
��N �
��N� ´��N� ´��N �
��N      C  , , ����N ����N� Ř��N� Ř��N ����N      C  , , ����N ����N� �|��N� �|��N ����N      C  , , �B��U �B��U� ����U� ����U �B��U      C  , , �&��U �&��U� ����U� ����U �&��U      C  , , �
��U �
��U� ´��U� ´��U �
��U      C  , , ����U ����U� Ř��U� Ř��U ����U      C  , , ����U ����U� �|��U� �|��U ����U      C  , , ����R@ ����R� �|��R� �|��R@ ����R@      C  , , �^��Vx �^��W" ���W" ���Vx �^��Vx      C  , , �B��Vx �B��W" ����W" ����Vx �B��Vx      C  , , �&��W� �&��X� ����X� ����W� �&��W�      C  , , �^��W� �^��X� ���X� ���W� �^��W�      C  , , �B��W� �B��X� ����X� ����W� �B��W�      C  , , ����R@ ����R� �\��R� �\��R@ ����R@      C  , , ����P� ����Q� �\��Q� �\��P� ����P�      C  , , ����P� ����Q� �@��Q� �@��P� ����P�      C  , , �z��P� �z��Q� �$��Q� �$��P� �z��P�      C  , , �^��P� �^��Q� ���Q� ���P� �^��P�      C  , , �B��P� �B��Q� ����Q� ����P� �B��P�      C  , , �&��P� �&��Q� ����Q� ����P� �&��P�      C  , , �
��P� �
��Q� ´��Q� ´��P� �
��P�      C  , , ����P� ����Q� Ř��Q� Ř��P� ����P�      C  , , ����P� ����Q� �|��Q� �|��P� ����P�      C  , , ����Vx ����W" �\��W" �\��Vx ����Vx      C  , , ����Vx ����W" �@��W" �@��Vx ����Vx      C  , , �z��Vx �z��W" �$��W" �$��Vx �z��Vx      C  , , ����Op ����P �\��P �\��Op ����Op      C  , , ����Op ����P �@��P �@��Op ����Op      C  , , �z��Op �z��P �$��P �$��Op �z��Op      C  , , �^��Op �^��P ���P ���Op �^��Op      C  , , �&��Vx �&��W" ����W" ����Vx �&��Vx      C  , , �
��Vx �
��W" ´��W" ´��Vx �
��Vx      C  , , ����Vx ����W" Ř��W" Ř��Vx ����Vx      C  , , ����Vx ����W" �|��W" �|��Vx ����Vx      C  , , �B��Op �B��P ����P ����Op �B��Op      C  , , �
��W� �
��X� ´��X� ´��W� �
��W�      C  , , ����YH ����Y� �\��Y� �\��YH ����YH      C  , , ����YH ����Y� �@��Y� �@��YH ����YH      C  , , �z��YH �z��Y� �$��Y� �$��YH �z��YH      C  , , �^��YH �^��Y� ���Y� ���YH �^��YH      C  , , �B��YH �B��Y� ����Y� ����YH �B��YH      C  , , �&��YH �&��Y� ����Y� ����YH �&��YH      C  , , �
��YH �
��Y� ´��Y� ´��YH �
��YH      C  , , ����YH ����Y� Ř��Y� Ř��YH ����YH      C  , , ����YH ����Y� �|��Y� �|��YH ����YH      C  , , �&��Op �&��P ����P ����Op �&��Op      C  , , �
��Op �
��P ´��P ´��Op �
��Op      C  , , ����Op ����P Ř��P Ř��Op ����Op      C  , , ����Op ����P �|��P �|��Op ����Op      C  , , ����R@ ����R� �@��R� �@��R@ ����R@      C  , , �z��R@ �z��R� �$��R� �$��R@ �z��R@      C  , , �^��R@ �^��R� ���R� ���R@ �^��R@      C  , , �B��R@ �B��R� ����R� ����R@ �B��R@      C  , , �&��R@ �&��R� ����R� ����R@ �&��R@      C  , , ����W� ����X� Ř��X� Ř��W� ����W�      C  , , ����W� ����X� �|��X� �|��W� ����W�      C  , , ����W� ����X� �\��X� �\��W� ����W�      C  , , ����W� ����X� �@��X� �@��W� ����W�      C  , , �z��W� �z��X� �$��X� �$��W� �z��W�      C  , , ����S� ����TR �\��TR �\��S� ����S�      C  , , ����S� ����TR �@��TR �@��S� ����S�      C  , , �z��S� �z��TR �$��TR �$��S� �z��S�      C  , , �^��S� �^��TR ���TR ���S� �^��S�      C  , , �B��S� �B��TR ����TR ����S� �B��S�      C  , , �&��S� �&��TR ����TR ����S� �&��S�      C  , , �
��S� �
��TR ´��TR ´��S� �
��S�      C  , , ����S� ����TR Ř��TR Ř��S� ����S�      C  , , ����L� ����MJ �\��MJ �\��L� ����L�      C  , , ����L� ����MJ �@��MJ �@��L� ����L�      C  , , �z��L� �z��MJ �$��MJ �$��L� �z��L�      C  , , �^��L� �^��MJ ���MJ ���L� �^��L�      C  , , �B��L� �B��MJ ����MJ ����L� �B��L�      C  , , �&��L� �&��MJ ����MJ ����L� �&��L�      C  , , �
��L� �
��MJ ´��MJ ´��L� �
��L�      C  , , ����L� ����MJ Ř��MJ Ř��L� ����L�      C  , , ����L� ����MJ �|��MJ �|��L� ����L�      D   , W  )" W  4 �  4 �  )" W  )"      D   , !  $� !  '� �  '� �  $� !  $�      D   , W  � W  #� �  #� �  � W  �      D   ,  ]�����  ]�����  ^�����  ^�����  ]�����      D   ,  _�����  _�����  aS����  aS����  _�����      D   ,  b/����  b/����  c�����  c�����  b/����      D   ,  d�����  d�����  e�����  e�����  d�����      D   ,  f�����  f�����  h3����  h3����  f�����      D   ,  i#����  i#����  j�����  j�����  i#����      D   ,  kg����  kg����  l�����  l�����  kg����      D   ,  m�����  m�����  o'����  o'����  m�����      D   ,  p����  p����  qk����  qk����  p����      D   ,  r[����  r[����  s�����  s�����  r[����      D   ,  t�����  t�����  v����  v����  t�����      D   ,  v�����  v�����  x_����  x_����  v�����      D   ,  y;����  y;����  z�����  z�����  y;����      D   ,  {�����  {�����  |�����  |�����  {�����      D   ,  }�����  }�����  ?����  ?����  }�����      D   ,  �/����  �/����  ������  ������  �/����      D   ,  �s����  �s����  ������  ������  �s����      D   ,  ������  ������  �3����  �3����  ������      D   ,  �����  �����  �w����  �w����  �����      D   ,  �g����  �g����  ������  ������  �g����      D   ,  ������  ������  �����  �����  ������      D   ,  �����  �����  �k����  �k����  �����      D   ,  �G����  �G����  ������  ������  �G����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �K����  �K����  ������      D   ,  �;����  �;����  ������  ������  �;����      D   ,  �����  �����  ������  ������  �����      D   ,  ������  ������  �?����  �?����  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �s����  �s����  ������  ������  �s����      D   ,  ������  ������  �����  �����  ������      D   ,  �����  �����  �w����  �w����  �����      D   ,  �S����  �S����  ������  ������  �S����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �W����  �W����  ������      D   ,  �G����  �G����  ������  ������  �G����      D   ,  ������  ������  ������  ������  ������      D   ,  ������  ������  �K����  �K����  ������      D   ,  �'����  �'����  ������  ������  �'����      D   ,  �����  �����  ������  ������  �����      D   ,  ������  ������  �+����  �+����  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �_����  �_����  ������  ������  �_����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �c����  �c����  ������      D   ,  �S����  �S����  ƻ����  ƻ����  �S����      D   ,  Ǘ����  Ǘ����  ������  ������  Ǘ����      D   ,  ������  ������  �W����  �W����  ������      D   ,  �3����  �3����  ͛����  ͛����  �3����      D   ,  ΋����  ΋����  ������  ������  ΋����      D   ,  ������  ������  �7����  �7����  ������      D   , N��^ N��a t��a t��^ N��^      D   , {�  4 {�  4v |�  4v |�  4 {�  4      D   , {�  )" {�  4 }  4 }  )" {�  )"      D   , {�  (� {�  )" |�  )" |�  (� {�  (�      D   , {�  #� {�  $" |�  $" |�  #� {�  #�      D   , {�  � {�  #� }  #� }  � {�  �      D   , {�  j {�  � |�  � |�  j {�  j      D   , �-  )" �-  4 ��  4 ��  )" �-  )"      D   , �E  $� �E  '� ��  '� ��  $� �E  $�      D   , �-  � �-  #� ��  #� ��  � �-  �      D   , ��  4 ��  4v ��  4v ��  4 ��  4      D   , ��  4 ��  4v ��  4v ��  4 ��  4      D   , �B  4 �B  4v �(  4v �(  4 �B  4      D   , ��  4 ��  4v �v  4v �v  4 ��  4      D   , ��  4 ��  4v ��  4v ��  4 ��  4      D   , �,  4 �,  4v �  4v �  4 �,  4      D   , �z  4 �z  4v �`  4v �`  4 �z  4      D   , ��  4 ��  4v Ȯ  4v Ȯ  4 ��  4      D   , �  4 �  4v ��  4v ��  4 �  4      D   , �d  4 �d  4v �J  4v �J  4 �d  4      D   , β  4 β  4v Ϙ  4v Ϙ  4 β  4      D   , ��  4 ��  4v ��  4v ��  4 ��  4      D   , �{  )" �{  4 ��  4 ��  )" �{  )"      D   , ��  )" ��  4 �1  4 �1  )" ��  )"      D   , �  )" �  4 �  4 �  )" �  )"      D   , �e  )" �e  4 ��  4 ��  )" �e  )"      D   , ��  )" ��  4 �  4 �  )" ��  )"      D   , �  )" �  4 �i  4 �i  )" �  )"      D   , �O  )" �O  4 ��  4 ��  )" �O  )"      D   , ��  )" ��  4 �  4 �  )" ��  )"      D   , ��  )" ��  4 �S  4 �S  )" ��  )"      D   , �9  )" �9  4 ơ  4 ơ  )" �9  )"      D   , Ǉ  )" Ǉ  4 ��  4 ��  )" Ǉ  )"      D   , ��  )" ��  4 �=  4 �=  )" ��  )"      D   , �#  )" �#  4 ͋  4 ͋  )" �#  )"      D   , �q  )" �q  4 ��  4 ��  )" �q  )"      D   , ��  (� ��  )" ��  )" ��  (� ��  (�      D   , �
  (� �
  )" ��  )" ��  (� �
  (�      D   , �X  (� �X  )" �>  )" �>  (� �X  (�      D   , ��  (� ��  )" ��  )" ��  (� ��  (�      D   , ��  (� ��  )" ��  )" ��  (� ��  (�      D   , �B  (� �B  )" �(  )" �(  (� �B  (�      D   , ��  (� ��  )" �v  )" �v  (� ��  (�      D   , ��  (� ��  )" ��  )" ��  (� ��  (�      D   , �,  (� �,  )" �  )" �  (� �,  (�      D   , �z  (� �z  )" �`  )" �`  (� �z  (�      D   , ��  (� ��  )" Ȯ  )" Ȯ  (� ��  (�      D   , �  (� �  )" ��  )" ��  (� �  (�      D   , �d  (� �d  )" �J  )" �J  (� �d  (�      D   , β  (� β  )" Ϙ  )" Ϙ  (� β  (�      D   , �
  4 �
  4v ��  4v ��  4 �
  4      D   , ��  $� ��  '� �  '� �  $� ��  $�      D   , ��  $� ��  '� �g  '� �g  $� ��  $�      D   , �/  $� �/  '� ��  '� ��  $� �/  $�      D   , �}  $� �}  '� �  '� �  $� �}  $�      D   , ��  $� ��  '� �Q  '� �Q  $� ��  $�      D   , �  $� �  '� ��  '� ��  $� �  $�      D   , �g  $� �g  '� ��  '� ��  $� �g  $�      D   , ��  $� ��  '� �;  '� �;  $� ��  $�      D   , �  $� �  '� ŉ  '� ŉ  $� �  $�      D   , �Q  $� �Q  '� ��  '� ��  $� �Q  $�      D   , ȟ  $� ȟ  '� �%  '� �%  $� ȟ  $�      D   , ��  $� ��  '� �s  '� �s  $� ��  $�      D   , �;  $� �;  '� ��  '� ��  $� �;  $�      D   , ��  #� ��  $" ��  $" ��  #� ��  #�      D   , �
  #� �
  $" ��  $" ��  #� �
  #�      D   , �X  #� �X  $" �>  $" �>  #� �X  #�      D   , ��  #� ��  $" ��  $" ��  #� ��  #�      D   , ��  #� ��  $" ��  $" ��  #� ��  #�      D   , �B  #� �B  $" �(  $" �(  #� �B  #�      D   , ��  #� ��  $" �v  $" �v  #� ��  #�      D   , ��  #� ��  $" ��  $" ��  #� ��  #�      D   , �,  #� �,  $" �  $" �  #� �,  #�      D   , �z  #� �z  $" �`  $" �`  #� �z  #�      D   , ��  #� ��  $" Ȯ  $" Ȯ  #� ��  #�      D   , �  #� �  $" ��  $" ��  #� �  #�      D   , �d  #� �d  $" �J  $" �J  #� �d  #�      D   , β  #� β  $" Ϙ  $" Ϙ  #� β  #�      D   , �X  4 �X  4v �>  4v �>  4 �X  4      D   , �{  � �{  #� ��  #� ��  � �{  �      D   , ��  � ��  #� �1  #� �1  � ��  �      D   , �  � �  #� �  #� �  � �  �      D   , �e  � �e  #� ��  #� ��  � �e  �      D   , ��  � ��  #� �  #� �  � ��  �      D   , �  � �  #� �i  #� �i  � �  �      D   , �O  � �O  #� ��  #� ��  � �O  �      D   , ��  � ��  #� �  #� �  � ��  �      D   , ��  � ��  #� �S  #� �S  � ��  �      D   , �9  � �9  #� ơ  #� ơ  � �9  �      D   , Ǉ  � Ǉ  #� ��  #� ��  � Ǉ  �      D   , ��  � ��  #� �=  #� �=  � ��  �      D   , �#  � �#  #� ͋  #� ͋  � �#  �      D   , �q  � �q  #� ��  #� ��  � �q  �      D   , ��  j ��  � ��  � ��  j ��  j      D   , �
  j �
  � ��  � ��  j �
  j      D   , �X  j �X  � �>  � �>  j �X  j      D   , ��  j ��  � ��  � ��  j ��  j      D   , ��  j ��  � ��  � ��  j ��  j      D   , �B  j �B  � �(  � �(  j �B  j      D   , ��  j ��  � �v  � �v  j ��  j      D   , ��  j ��  � ��  � ��  j ��  j      D   , �,  j �,  � �  � �  j �,  j      D   , �z  j �z  � �`  � �`  j �z  j      D   , ��  j ��  � Ȯ  � Ȯ  j ��  j      D   , �  j �  � ��  � ��  j �  j      D   , �d  j �d  � �J  � �J  j �d  j      D   , β  j β  � Ϙ  � Ϙ  j β  j      D   , �'  � �'  4� �]  4� �]  � �'  �      D   , }�  � }�  #� R  #� R  � }�  �      D   , ~+  (� ~+  )"   )"   (� ~+  (�      D   , ~+  j ~+  �   �   j ~+  j      D   , ��  � ��  4� ��  4� ��  � ��  �      D   , ��  4 ��  4v ��  4v ��  4 ��  4      D   , ��  4 ��  4v ��  4v ��  4 ��  4      D   , �  #� �  $" ��  $" ��  #� �  #�      D   , �b  #� �b  $" �H  $" �H  #� �b  #�      D   , ��  #� ��  $" ��  $" ��  #� ��  #�      D   , ��  #� ��  $" ��  $" ��  #� ��  #�      D   , �L  #� �L  $" �2  $" �2  #� �L  #�      D   , ��  #� ��  $" ��  $" ��  #� ��  #�      D   , ��  #� ��  $" ��  $" ��  #� ��  #�      D   , �6  #� �6  $" �  $" �  #� �6  #�      D   , ��  #� ��  $" �j  $" �j  #� ��  #�      D   , ��  #� ��  $" ��  $" ��  #� ��  #�      D   , �   #� �   $" �  $" �  #� �   #�      D   , �n  #� �n  $" �T  $" �T  #� �n  #�      D   , �L  4 �L  4v �2  4v �2  4 �L  4      D   , ��  (� ��  )" ��  )" ��  (� ��  (�      D   , ��  (� ��  )" ��  )" ��  (� ��  (�      D   , �L  (� �L  )" �2  )" �2  (� �L  (�      D   , ��  (� ��  )" ��  )" ��  (� ��  (�      D   , ��  (� ��  )" ��  )" ��  (� ��  (�      D   , �6  (� �6  )" �  )" �  (� �6  (�      D   , ��  (� ��  )" �j  )" �j  (� ��  (�      D   , ��  (� ��  )" ��  )" ��  (� ��  (�      D   , �   (� �   )" �  )" �  (� �   (�      D   , �n  (� �n  )" �T  )" �T  (� �n  (�      D   , ��  4 ��  4v ��  4v ��  4 ��  4      D   , ��  4 ��  4v ��  4v ��  4 ��  4      D   , �6  4 �6  4v �  4v �  4 �6  4      D   , ��  � ��  #� �;  #� �;  � ��  �      D   , �!  � �!  #� ��  #� ��  � �!  �      D   , �o  � �o  #� ��  #� ��  � �o  �      D   , ��  � ��  #� �%  #� �%  � ��  �      D   , �  � �  #� �s  #� �s  � �  �      D   , �Y  � �Y  #� ��  #� ��  � �Y  �      D   , ��  � ��  #� �  #� �  � ��  �      D   , ��  � ��  #� �]  #� �]  � ��  �      D   , �C  � �C  #� ��  #� ��  � �C  �      D   , ��  � ��  #� ��  #� ��  � ��  �      D   , ��  � ��  #� �G  #� �G  � ��  �      D   , ��  )" ��  4 �;  4 �;  )" ��  )"      D   , �!  )" �!  4 ��  4 ��  )" �!  )"      D   , �o  )" �o  4 ��  4 ��  )" �o  )"      D   , ��  )" ��  4 �%  4 �%  )" ��  )"      D   , �  )" �  4 �s  4 �s  )" �  )"      D   , �Y  )" �Y  4 ��  4 ��  )" �Y  )"      D   , ��  )" ��  4 �  4 �  )" ��  )"      D   , ��  )" ��  4 �]  4 �]  )" ��  )"      D   , �C  )" �C  4 ��  4 ��  )" �C  )"      D   , ��  )" ��  4 ��  4 ��  )" ��  )"      D   , ��  )" ��  4 �G  4 �G  )" ��  )"      D   , ��  $� ��  '� �q  '� �q  $� ��  $�      D   , �9  $� �9  '� ��  '� ��  $� �9  $�      D   , ��  $� ��  '� �  '� �  $� ��  $�      D   , ��  $� ��  '� �[  '� �[  $� ��  $�      D   , �  j �  � ��  � ��  j �  j      D   , �b  j �b  � �H  � �H  j �b  j      D   , ��  j ��  � ��  � ��  j ��  j      D   , ��  j ��  � ��  � ��  j ��  j      D   , �L  j �L  � �2  � �2  j �L  j      D   , ��  j ��  � ��  � ��  j ��  j      D   , ��  j ��  � ��  � ��  j ��  j      D   , �6  j �6  � �  � �  j �6  j      D   , ��  j ��  � �j  � �j  j ��  j      D   , ��  j ��  � ��  � ��  j ��  j      D   , �   j �   � �  � �  j �   j      D   , �n  j �n  � �T  � �T  j �n  j      D   , �#  $� �#  '� ��  '� ��  $� �#  $�      D   , �q  $� �q  '� ��  '� ��  $� �q  $�      D   , ��  $� ��  '� �E  '� �E  $� ��  $�      D   , �  $� �  '� ��  '� ��  $� �  $�      D   , �[  $� �[  '� ��  '� ��  $� �[  $�      D   , ��  $� ��  '� �/  '� �/  $� ��  $�      D   , ��  $� ��  '� �}  '� �}  $� ��  $�      D   , ��  4 ��  4v �j  4v �j  4 ��  4      D   , ��  4 ��  4v ��  4v ��  4 ��  4      D   , �   4 �   4v �  4v �  4 �   4      D   , �n  4 �n  4v �T  4v �T  4 �n  4      D   , |�  $� |�  '� ~:  '� ~:  $� |�  $�      D   , }�  )" }�  4 R  4 R  )" }�  )"      D   , ~+  #� ~+  $"   $"   #� ~+  #�      D   , ~+  4 ~+  4v   4v   4 ~+  4      D   , I)  4 I)  4v J  4v J  4 I)  4      D   , H�  )" H�  4 JP  4 JP  )" H�  )"      D   , I)  (� I)  )" J  )" J  (� I)  (�      D   , I)  #� I)  $" J  $" J  #� I)  #�      D   , H�  � H�  #� JP  #� JP  � H�  �      D   , I)  j I)  � J  � J  j I)  j      D   , b�  4 b�  4v ci  4v ci  4 b�  4      D   , bB  )" bB  4 c�  4 c�  )" bB  )"      D   , b�  (� b�  )" ci  )" ci  (� b�  (�      D   , J   $� J   '� K�  '� K�  $� J   $�      D   , LN  $� LN  '� M�  '� M�  $� LN  $�      D   , N�  $� N�  '� P"  '� P"  $� N�  $�      D   , P�  $� P�  '� Rp  '� Rp  $� P�  $�      D   , S8  $� S8  '� T�  '� T�  $� S8  $�      D   , U�  $� U�  '� W  '� W  $� U�  $�      D   , W�  $� W�  '� YZ  '� YZ  $� W�  $�      D   , Z"  $� Z"  '� [�  '� [�  $� Z"  $�      D   , \p  $� \p  '� ]�  '� ]�  $� \p  $�      D   , ^�  $� ^�  '� `D  '� `D  $� ^�  $�      D   , a  $� a  '� b�  '� b�  $� a  $�      D   , cZ  $� cZ  '� d�  '� d�  $� cZ  $�      D   , e�  $� e�  '� g.  '� g.  $� e�  $�      D   , g�  $� g�  '� i|  '� i|  $� g�  $�      D   , jD  $� jD  '� k�  '� k�  $� jD  $�      D   , l�  $� l�  '� n  '� n  $� l�  $�      D   , n�  $� n�  '� pf  '� pf  $� n�  $�      D   , q.  $� q.  '� r�  '� r�  $� q.  $�      D   , s|  $� s|  '� u  '� u  $� s|  $�      D   , u�  $� u�  '� wP  '� wP  $� u�  $�      D   , x  $� x  '� y�  '� y�  $� x  $�      D   , zf  $� zf  '� {�  '� {�  $� zf  $�      D   , b�  #� b�  $" ci  $" ci  #� b�  #�      D   , bB  � bB  #� c�  #� c�  � bB  �      D   , b�  j b�  � ci  � ci  j b�  j      D   , pW  (� pW  )" q=  )" q=  (� pW  (�      D   , r�  (� r�  )" s�  )" s�  (� r�  (�      D   , t�  (� t�  )" u�  )" u�  (� t�  (�      D   , wA  (� wA  )" x'  )" x'  (� wA  (�      D   , y�  (� y�  )" zu  )" zu  (� y�  (�      D   , im  4 im  4v jS  4v jS  4 im  4      D   , k�  4 k�  4v l�  4v l�  4 k�  4      D   , n	  4 n	  4v n�  4v n�  4 n	  4      D   , pW  4 pW  4v q=  4v q=  4 pW  4      D   , r�  4 r�  4v s�  4v s�  4 r�  4      D   , t�  4 t�  4v u�  4v u�  4 t�  4      D   , wA  4 wA  4v x'  4v x'  4 wA  4      D   , y�  4 y�  4v zu  4v zu  4 y�  4      D   , d�  4 d�  4v e�  4v e�  4 d�  4      D   , d�  )" d�  4 e�  4 e�  )" d�  )"      D   , f�  )" f�  4 hF  4 hF  )" f�  )"      D   , i,  )" i,  4 j�  4 j�  )" i,  )"      D   , kz  )" kz  4 l�  4 l�  )" kz  )"      D   , m�  )" m�  4 o0  4 o0  )" m�  )"      D   , p  )" p  4 q~  4 q~  )" p  )"      D   , rd  )" rd  4 s�  4 s�  )" rd  )"      D   , t�  )" t�  4 v  4 v  )" t�  )"      D   , w   )" w   4 xh  4 xh  )" w   )"      D   , yN  )" yN  4 z�  4 z�  )" yN  )"      D   , g  4 g  4v h  4v h  4 g  4      D   , d�  (� d�  )" e�  )" e�  (� d�  (�      D   , g  (� g  )" h  )" h  (� g  (�      D   , im  (� im  )" jS  )" jS  (� im  (�      D   , k�  (� k�  )" l�  )" l�  (� k�  (�      D   , n	  (� n	  )" n�  )" n�  (� n	  (�      D   , [X  )" [X  4 \�  4 \�  )" [X  )"      D   , ]�  )" ]�  4 _  4 _  )" ]�  )"      D   , _�  )" _�  4 a\  4 a\  )" _�  )"      D   , M�  4 M�  4v N�  4v N�  4 M�  4      D   , P  4 P  4v P�  4v P�  4 P  4      D   , Ra  4 Ra  4v SG  4v SG  4 Ra  4      D   , T�  4 T�  4v U�  4v U�  4 T�  4      D   , V�  4 V�  4v W�  4v W�  4 V�  4      D   , YK  4 YK  4v Z1  4v Z1  4 YK  4      D   , [�  4 [�  4v \  4v \  4 [�  4      D   , ]�  4 ]�  4v ^�  4v ^�  4 ]�  4      D   , `5  4 `5  4v a  4v a  4 `5  4      D   , Kw  4 Kw  4v L]  4v L]  4 Kw  4      D   , K6  )" K6  4 L�  4 L�  )" K6  )"      D   , Kw  (� Kw  )" L]  )" L]  (� Kw  (�      D   , M�  (� M�  )" N�  )" N�  (� M�  (�      D   , P  (� P  )" P�  )" P�  (� P  (�      D   , Ra  (� Ra  )" SG  )" SG  (� Ra  (�      D   , T�  (� T�  )" U�  )" U�  (� T�  (�      D   , V�  (� V�  )" W�  )" W�  (� V�  (�      D   , YK  (� YK  )" Z1  )" Z1  (� YK  (�      D   , [�  (� [�  )" \  )" \  (� [�  (�      D   , ]�  (� ]�  )" ^�  )" ^�  (� ]�  (�      D   , `5  (� `5  )" a  )" a  (� `5  (�      D   , M�  )" M�  4 N�  4 N�  )" M�  )"      D   , O�  )" O�  4 Q:  4 Q:  )" O�  )"      D   , R   )" R   4 S�  4 S�  )" R   )"      D   , Tn  )" Tn  4 U�  4 U�  )" Tn  )"      D   , V�  )" V�  4 X$  4 X$  )" V�  )"      D   , Y
  )" Y
  4 Zr  4 Zr  )" Y
  )"      D   , Ra  #� Ra  $" SG  $" SG  #� Ra  #�      D   , T�  #� T�  $" U�  $" U�  #� T�  #�      D   , V�  #� V�  $" W�  $" W�  #� V�  #�      D   , YK  #� YK  $" Z1  $" Z1  #� YK  #�      D   , [�  #� [�  $" \  $" \  #� [�  #�      D   , ]�  #� ]�  $" ^�  $" ^�  #� ]�  #�      D   , `5  #� `5  $" a  $" a  #� `5  #�      D   , Kw  #� Kw  $" L]  $" L]  #� Kw  #�      D   , K6  � K6  #� L�  #� L�  � K6  �      D   , M�  � M�  #� N�  #� N�  � M�  �      D   , O�  � O�  #� Q:  #� Q:  � O�  �      D   , R   � R   #� S�  #� S�  � R   �      D   , Tn  � Tn  #� U�  #� U�  � Tn  �      D   , V�  � V�  #� X$  #� X$  � V�  �      D   , Y
  � Y
  #� Zr  #� Zr  � Y
  �      D   , [X  � [X  #� \�  #� \�  � [X  �      D   , ]�  � ]�  #� _  #� _  � ]�  �      D   , _�  � _�  #� a\  #� a\  � _�  �      D   , M�  #� M�  $" N�  $" N�  #� M�  #�      D   , Kw  j Kw  � L]  � L]  j Kw  j      D   , M�  j M�  � N�  � N�  j M�  j      D   , P  j P  � P�  � P�  j P  j      D   , Ra  j Ra  � SG  � SG  j Ra  j      D   , T�  j T�  � U�  � U�  j T�  j      D   , V�  j V�  � W�  � W�  j V�  j      D   , YK  j YK  � Z1  � Z1  j YK  j      D   , [�  j [�  � \  � \  j [�  j      D   , ]�  j ]�  � ^�  � ^�  j ]�  j      D   , `5  j `5  � a  � a  j `5  j      D   , P  #� P  $" P�  $" P�  #� P  #�      D   , k�  #� k�  $" l�  $" l�  #� k�  #�      D   , n	  #� n	  $" n�  $" n�  #� n	  #�      D   , pW  #� pW  $" q=  $" q=  #� pW  #�      D   , r�  #� r�  $" s�  $" s�  #� r�  #�      D   , d�  � d�  #� e�  #� e�  � d�  �      D   , f�  � f�  #� hF  #� hF  � f�  �      D   , i,  � i,  #� j�  #� j�  � i,  �      D   , kz  � kz  #� l�  #� l�  � kz  �      D   , m�  � m�  #� o0  #� o0  � m�  �      D   , p  � p  #� q~  #� q~  � p  �      D   , rd  � rd  #� s�  #� s�  � rd  �      D   , t�  � t�  #� v  #� v  � t�  �      D   , w   � w   #� xh  #� xh  � w   �      D   , yN  � yN  #� z�  #� z�  � yN  �      D   , y�  j y�  � zu  � zu  j y�  j      D   , t�  #� t�  $" u�  $" u�  #� t�  #�      D   , wA  #� wA  $" x'  $" x'  #� wA  #�      D   , y�  #� y�  $" zu  $" zu  #� y�  #�      D   , wA  j wA  � x'  � x'  j wA  j      D   , t�  j t�  � u�  � u�  j t�  j      D   , n	  j n	  � n�  � n�  j n	  j      D   , r�  j r�  � s�  � s�  j r�  j      D   , pW  j pW  � q=  � q=  j pW  j      D   , d�  #� d�  $" e�  $" e�  #� d�  #�      D   , g  #� g  $" h  $" h  #� g  #�      D   , im  #� im  $" jS  $" jS  #� im  #�      D   , d�  j d�  � e�  � e�  j d�  j      D   , g  j g  � h  � h  j g  j      D   , im  j im  � jS  � jS  j im  j      D   , k�  j k�  � l�  � l�  j k�  j      D   , -�  j -�  � .�  � .�  j -�  j      D   , 1  � 1  4� AO  4� AO  � 1  �      D   , �  j �  � ~  � ~  j �  j      D   , �  j �  � �  � �  j �  j      D   , 4  j 4  �   �   j 4  j      D   , �  j �  � h  � h  j �  j      D   , �  � �  #� [  #� [  � �  �      D   , A  � A  #� �  #� �  � A  �      D   , �  j �  �  �  �  �  j �  j      D   , "  j "  � #  � #  j "  j      D   , $l  j $l  � %R  � %R  j $l  j      D   , &�  j &�  � '�  � '�  j &�  j      D   , �  � �  #�  �  #�  �  � �  �      D   , +  � +  #� ,}  #� ,}  � +  �      D   , -c  � -c  #� .�  #� .�  � -c  �      D   , D�  j D�  � Es  � Es  j D�  j      D   , F�  j F�  � G�  � G�  j F�  j      D   , !�  � !�  #� #E  #� #E  � !�  �      D   , Ed  $� Ed  '� F�  '� F�  $� Ed  $�      D   , G�  $� G�  '� I8  '� I8  $� G�  $�      D   , &y  � &y  #� '�  #� '�  � &y  �      D   , (�  � (�  #� */  #� */  � (�  �      D   , DL  � DL  #� E�  #� E�  � DL  �      D   , F�  � F�  #� H  #� H  � F�  �      D   , $+  � $+  #� %�  #� %�  � $+  �      D   , D�  #� D�  $" Es  $" Es  #� D�  #�      D   , F�  #� F�  $" G�  $" G�  #� F�  #�      D   , )  j )  � )�  � )�  j )  j      D   , +V  j +V  � ,<  � ,<  j +V  j      D   , 4  4 4  4v   4v   4 4  4      D   , �  � �  #�   #�   � �  �      D   , DL  )" DL  4 E�  4 E�  )" DL  )"      D   , F�  )" F�  4 H  4 H  )" F�  )"      D   , �  4 �  4v h  4v h  4 �  4      D   , �  4 �  4v  �  4v  �  4 �  4      D   , "  4 "  4v #  4v #  4 "  4      D   , $l  4 $l  4v %R  4v %R  4 $l  4      D   , &�  4 &�  4v '�  4v '�  4 &�  4      D   , )  4 )  4v )�  4v )�  4 )  4      D   , +V  4 +V  4v ,<  4v ,<  4 +V  4      D   , -�  4 -�  4v .�  4v .�  4 -�  4      D   , �  4 �  4v ~  4v ~  4 �  4      D   , �  )" �  4   4   )" �  )"      D   , �  )" �  4 [  4 [  )" �  )"      D   , A  )" A  4 �  4 �  )" A  )"      D   , �  )" �  4  �  4  �  )" �  )"      D   , !�  )" !�  4 #E  4 #E  )" !�  )"      D   , $+  )" $+  4 %�  4 %�  )" $+  )"      D   , &y  )" &y  4 '�  4 '�  )" &y  )"      D   , (�  )" (�  4 */  4 */  )" (�  )"      D   , +  )" +  4 ,}  4 ,}  )" +  )"      D   , -c  )" -c  4 .�  4 .�  )" -c  )"      D   , �  (� �  )" ~  )" ~  (� �  (�      D   , �  (� �  )" �  )" �  (� �  (�      D   , 4  (� 4  )"   )"   (� 4  (�      D   , �  (� �  )" h  )" h  (� �  (�      D   , �  (� �  )"  �  )"  �  (� �  (�      D   , "  (� "  )" #  )" #  (� "  (�      D   , $l  (� $l  )" %R  )" %R  (� $l  (�      D   , &�  (� &�  )" '�  )" '�  (� &�  (�      D   , )  (� )  )" )�  )" )�  (� )  (�      D   , +V  (� +V  )" ,<  )" ,<  (� +V  (�      D   , -�  (� -�  )" .�  )" .�  (� -�  (�      D   , �  4 �  4v �  4v �  4 �  4      D   , o  $� o  '� �  '� �  $� o  $�      D   , �  $� �  '� C  '� C  $� �  $�      D   ,   $�   '� �  '� �  $�   $�      D   , Y  $� Y  '� �  '� �  $� Y  $�      D   ,  �  $�  �  '� "-  '� "-  $�  �  $�      D   , "�  $� "�  '� ${  '� ${  $� "�  $�      D   , %C  $� %C  '� &�  '� &�  $� %C  $�      D   , '�  $� '�  '� )  '� )  $� '�  $�      D   , )�  $� )�  '� +e  '� +e  $� )�  $�      D   , ,-  $� ,-  '� -�  '� -�  $� ,-  $�      D   , �  #� �  $" ~  $" ~  #� �  #�      D   , �  #� �  $" �  $" �  #� �  #�      D   , 4  #� 4  $"   $"   #� 4  #�      D   , �  #� �  $" h  $" h  #� �  #�      D   , �  #� �  $"  �  $"  �  #� �  #�      D   , "  #� "  $" #  $" #  #� "  #�      D   , $l  #� $l  $" %R  $" %R  #� $l  #�      D   , &�  #� &�  $" '�  $" '�  #� &�  #�      D   , )  #� )  $" )�  $" )�  #� )  #�      D   , +V  #� +V  $" ,<  $" ,<  #� +V  #�      D   , -�  #� -�  $" .�  $" .�  #� -�  #�      D   ,  �!  L  �!  `  �1  `  �1  L  �!  L      D   ,  ��  3  ��  L  �1  L  �1  3  ��  3      D   ,  \�  5  \�  3  �  3  �  5  \�  5      D   ,  �U  �  �U  
�  ��  
�  ��  �  �U  �      D   ,  \�����  \�����  ������  ������  \�����      D   ,  �U��߭  �U���  �����  ����߭  �U��߭      D   ,  \�����  \���У  ����У  ������  \�����      D   ,  ��  �  ��  #�  �-  #�  �-  �  ��  �      D   ,  �  �  �  #�  �{  #�  �{  �  �  �      D   ,  �a  �  �a  #�  ��  #�  ��  �  �a  �      D   ,  ��  �  ��  #�  �  #�  �  �  ��  �      D   ,  ��  �  ��  #�  �e  #�  �e  �  ��  �      D   ,  �K  �  �K  #�  �  #�  �  �  �K  �      D   , �  � �  #�   #�   � �  �      D   , �  � �  #� O  #� O  � �  �      D   , 5  � 5  #� �  #� �  � 5  �      D   , �  � �  #� 	�  #� 	�  � �  �      D   , 
�  � 
�  #� 9  #� 9  � 
�  �      D   ,   �   #� �  #� �  �   �      D   , m  � m  #� �  #� �  � m  �      D   , �  � �  #� #  #� #  � �  �      D   , 	  � 	  #� q  #� q  � 	  �      D   , �  (� �  )" �  )" �  (� �  (�      D   , (  (� (  )"   )"   (� (  (�      D   , v  (� v  )" \  )" \  (� v  (�      D   , �  (� �  )" 	�  )" 	�  (� �  (�      D   ,   (�   )" �  )" �  (�   (�      D   , `  (� `  )" F  )" F  (� `  (�      D   , �  (� �  )" �  )" �  (� �  (�      D   , �  (� �  )" �  )" �  (� �  (�      D   , J  (� J  )" 0  )" 0  (� J  (�      D   , �  4 �  4v 	�  4v 	�  4 �  4      D   ,   4   4v �  4v �  4   4      D   ,  �  j  �  �  ��  �  ��  j  �  j      D   ,  �T  j  �T  �  �:  �  �:  j  �T  j      D   ,  ��  j  ��  �  ��  �  ��  j  ��  j      D   ,  ��  j  ��  �  ��  �  ��  j  ��  j      D   ,  �>  j  �>  �  �$  �  �$  j  �>  j      D   ,  ��  j  ��  �  r  �  r  j  ��  j      D   , �  j �  � �  � �  j �  j      D   , (  j (  �   �   j (  j      D   , v  j v  � \  � \  j v  j      D   , �  j �  � 	�  � 	�  j �  j      D   ,   j   � �  � �  j   j      D   , `  j `  � F  � F  j `  j      D   , �  j �  � �  � �  j �  j      D   , �  j �  � �  � �  j �  j      D   , J  j J  � 0  � 0  j J  j      D   , `  4 `  4v F  4v F  4 `  4      D   ,  ��  )"  ��  4  �-  4  �-  )"  ��  )"      D   ,  �  )"  �  4  �{  4  �{  )"  �  )"      D   ,  �a  )"  �a  4  ��  4  ��  )"  �a  )"      D   ,  ��  )"  ��  4  �  4  �  )"  ��  )"      D   ,  ��  )"  ��  4  �e  4  �e  )"  ��  )"      D   ,  �K  )"  �K  4  �  4  �  )"  �K  )"      D   , �  )" �  4   4   )" �  )"      D   , �  )" �  4 O  4 O  )" �  )"      D   ,  ��  $�  ��  '�  �c  '�  �c  $�  ��  $�      D   ,  �+  $�  �+  '�  ��  '�  ��  $�  �+  $�      D   ,  �y  $�  �y  '�  ��  '�  ��  $�  �y  $�      D   ,  ��  $�  ��  '�  �M  '�  �M  $�  ��  $�      D   ,  �  $�  �  '�  ��  '�  ��  $�  �  $�      D   ,  c  $�  c  '� �  '� �  $�  c  $�      D   , �  $� �  '� 7  '� 7  $� �  $�      D   , �  $� �  '� �  '� �  $� �  $�      D   , M  $� M  '� �  '� �  $� M  $�      D   , 	�  $� 	�  '� !  '� !  $� 	�  $�      D   , �  $� �  '� o  '� o  $� �  $�      D   , 7  $� 7  '� �  '� �  $� 7  $�      D   , �  $� �  '�   '�   $� �  $�      D   , �  $� �  '� Y  '� Y  $� �  $�      D   , 5  )" 5  4 �  4 �  )" 5  )"      D   , �  )" �  4 	�  4 	�  )" �  )"      D   , 
�  )" 
�  4 9  4 9  )" 
�  )"      D   ,   )"   4 �  4 �  )"   )"      D   , m  )" m  4 �  4 �  )" m  )"      D   , �  )" �  4 #  4 #  )" �  )"      D   , 	  )" 	  4 q  4 q  )" 	  )"      D   , �  4 �  4v �  4v �  4 �  4      D   , �  4 �  4v �  4v �  4 �  4      D   , J  4 J  4v 0  4v 0  4 J  4      D   ,  �  #�  �  $"  ��  $"  ��  #�  �  #�      D   ,  �T  #�  �T  $"  �:  $"  �:  #�  �T  #�      D   ,  ��  #�  ��  $"  ��  $"  ��  #�  ��  #�      D   ,  ��  #�  ��  $"  ��  $"  ��  #�  ��  #�      D   ,  �>  #�  �>  $"  �$  $"  �$  #�  �>  #�      D   ,  ��  #�  ��  $"  r  $"  r  #�  ��  #�      D   , �  #� �  $" �  $" �  #� �  #�      D   , (  #� (  $"   $"   #� (  #�      D   , v  #� v  $" \  $" \  #� v  #�      D   , �  #� �  $" 	�  $" 	�  #� �  #�      D   ,   #�   $" �  $" �  #�   #�      D   , `  #� `  $" F  $" F  #� `  #�      D   , �  #� �  $" �  $" �  #� �  #�      D   , �  #� �  $" �  $" �  #� �  #�      D   , J  #� J  $" 0  $" 0  #� J  #�      D   ,  ��  4  ��  4v  ��  4v  ��  4  ��  4      D   ,  ��  4  ��  4v  ��  4v  ��  4  ��  4      D   ,  �>  4  �>  4v  �$  4v  �$  4  �>  4      D   ,  ��  4  ��  4v  r  4v  r  4  ��  4      D   , �  4 �  4v �  4v �  4 �  4      D   , (  4 (  4v   4v   4 (  4      D   , v  4 v  4v \  4v \  4 v  4      D   ,  ��  (�  ��  )"  ��  )"  ��  (�  ��  (�      D   ,  ��  (�  ��  )"  ��  )"  ��  (�  ��  (�      D   ,  �>  (�  �>  )"  �$  )"  �$  (�  �>  (�      D   ,  ��  (�  ��  )"  r  )"  r  (�  ��  (�      D   ,  �=  &   �=  '�  ��  '�  ��  &   �=  &       D   ,  ��  &   ��  '�  �  '�  �  &   ��  &       D   ,  ��  &   ��  '�  �_  '�  �_  &   ��  &       D   ,  �'  &   �'  '�  ��  '�  ��  &   �'  &       D   ,  ��  3  ��  �  ��  �  ��  3  ��  3      D   ,  �e  3  �e  �  �i  �  �i  3  �e  3      D   ,  �  3  �  �  �  �  �  3  �  3      D   ,  �-  `  �-  �  �1  �  �1  `  �-  `      D   ,  �u  &   �u  '�  ��  '�  ��  &   �u  &       D   ,  ��  &   ��  '�  �I  '�  �I  &   ��  &       D   ,  �  &   �  '�    '�    &   �  &       D   ,  �_  &   �_  '�  ��  '�  ��  &   �_  &       D   ,  ŭ  &   ŭ  '�  �3  '�  �3  &   ŭ  &       D   ,  ��  &   ��  '�  Ɂ  '�  Ɂ  &   ��  &       D   ,  ��  �  ��  5  ��  5  ��  �  ��  �      D   ,  ��  �  ��  5  ��  5  ��  �  ��  �      D   ,  �-  �  �-  5  �1  5  �1  �  �-  �      D   ,  ��  �  ��  5  ��  5  ��  �  ��  �      D   ,  �e  �  �e  5  �i  5  �i  �  �e  �      D   ,  �  �  �  5  �  5  �  �  �  �      D   ,  ��  �  ��  5  ��  5  ��  �  ��  �      D   ,  �Y  �  �Y  5  �]  5  �]  �  �Y  �      D   ,  �!  '�  �!  '�  �C  '�  �C  '�  �!  '�      D   ,  �o  '�  �o  '�  ��  '�  ��  '�  �o  '�      D   ,  ��  '�  ��  '�  ��  '�  ��  '�  ��  '�      D   ,  �  '�  �  '�  �-  '�  �-  '�  �  '�      D   ,  �Y  '�  �Y  '�  �{  '�  �{  '�  �Y  '�      D   ,  ��  '�  ��  '�  ��  '�  ��  '�  ��  '�      D   ,  ��  '�  ��  '�  �  '�  �  '�  ��  '�      D   ,  �C  '�  �C  '�  �e  '�  �e  '�  �C  '�      D   ,  Ñ  '�  Ñ  '�  ĳ  '�  ĳ  '�  Ñ  '�      D   ,  ��  '�  ��  '�  �  '�  �  '�  ��  '�      D   ,  �-  '�  �-  '�  �O  '�  �O  '�  �-  '�      D   ,  ��  &   ��  '�  �u  '�  �u  &   ��  &       D   ,  ��  e  ��  �  ��  �  ��  e  ��  e      D   ,  �Y  e  �Y  �  �]  �  �]  e  �Y  e      D   ,  ��  `  ��  e  �]  e  �]  `  ��  `      D   ,  ��  e  ��  �  ��  �  ��  e  ��  e      D   ,  ��  e  ��  �  ��  �  ��  e  ��  e      D   ,  ��  `  ��  e  ��  e  ��  `  ��  `      D   ,  ��  �  ��  
�  �)  
�  �)  �  ��  �      D   ,  ��  �  ��  
�  �w  
�  �w  �  ��  �      D   ,  �?  �  �?  
�  ��  
�  ��  �  �?  �      D   ,  ��  �  ��  
�  �  
�  �  �  ��  �      D   ,  ��  �  ��  
�  �a  
�  �a  �  ��  �      D   ,  �)  �  �)  
�  ��  
�  ��  �  �)  �      D   ,  �w  �  �w  
�  ��  
�  ��  �  �w  �      D   ,  ��  �  ��  
�  �K  
�  �K  �  ��  �      D   ,  �  �  �  
�  ř  
�  ř  �  �  �      D   ,  �a  �  �a  
�  ��  
�  ��  �  �a  �      D   ,  ȯ  �  ȯ  
�  �5  
�  �5  �  ȯ  �      D   ,  ��  �  ��  
�  ̃  
�  ̃  �  ��  �      D   ,  �K  �  �K  
�  ��  
�  ��  �  �K  �      D   ,  ϙ  �  ϙ  
�  �  
�  �  �  ϙ  �      D   ,  ������  ��  �  �C  �  �C����  ������      D   ,  ��  �  ��  �  �C  �  �C  �  ��  �      D   ,  �&  �  �&  �  �  �  �  �  �&  �      D   ,  �t  �  �t  �  �Z  �  �Z  �  �t  �      D   ,  ��  �  ��  �  Ϩ  �  Ϩ  �  ��  �      D   ,  �&  �  �&  >  �  >  �  �  �&  �      D   ,  �t  �  �t  >  �Z  >  �Z  �  �t  �      D   ,  ��  �  ��  >  Ϩ  >  Ϩ  �  ��  �      D   ,  �  �  �  >  ��  >  ��  �  �  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  �3  �  �3  �  ͛  �  ͛  �  �3  �      D   ,  �w  �  �w  �  ��  �  ��  �  �w  �      D   ,  ��  �  ��  �  �7  �  �7  �  ��  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  �  �  �  >  ��  >  ��  �  �  �      D   ,  �R  �  �R  >  �8  >  �8  �  �R  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  �<  �  �<  >  �"  >  �"  �  �<  �      D   ,  Ŋ  �  Ŋ  >  �p  >  �p  �  Ŋ  �      D   ,  ��  �  ��  >  Ⱦ  >  Ⱦ  �  ��  �      D   ,  �<  �  �<  �  �"  �  �"  �  �<  �      D   ,  Ŋ  �  Ŋ  �  �p  �  �p  �  Ŋ  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  ��  �  ��  �  Ⱦ  �  Ⱦ  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  ��  �  ��  �  �7  �  �7  �  ��  �      D   ,  �'  �  �'  �  ��  �  ��  �  �'  �      D   ,  �k  �  �k  �  ��  �  ��  �  �k  �      D   ,  ��  �  ��  �  �+  �  �+  �  ��  �      D   ,  �  �  �  �  �o  �  �o  �  �  �      D   ,  �_  �  �_  �  ��  �  ��  �  �_  �      D   ,  ��  �  ��  �  �  �  �  �  ��  �      D   ,  ��  �  ��  �  �c  �  �c  �  ��  �      D   ,  �?  �  �?  �  Ƨ  �  Ƨ  �  �?  �      D   ,  Ǘ  �  Ǘ  �  ��  �  ��  �  Ǘ  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �  �  �  >  �   >  �   �  �  �      D   ,  �h  �  �h  >  �N  >  �N  �  �h  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �  �  �  �  �   �  �   �  �  �      D   ,  �h  �  �h  �  �N  �  �N  �  �h  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  �R  �  �R  �  �8  �  �8  �  �R  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  �R  �  �R  �  �8  �  �8  �  �R  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �<  �  �<  �  �"  �  �"  �  �<  �      D   ,  Ŋ  �  Ŋ  �  �p  �  �p  �  Ŋ  �      D   ,  ��  �  ��  �  Ⱦ  �  Ⱦ  �  ��  �      D   ,  ������  ��  �  ��  �  ������  ������      D   ,  ������  ��  �  �7  �  �7����  ������      D   ,  �'����  �'  �  ��  �  ������  �'����      D   ,  �k����  �k  �  ��  �  ������  �k����      D   ,  ������  ��  �  �+  �  �+����  ������      D   ,  �����  �  �  �o  �  �o����  �����      D   ,  �_����  �_  �  ��  �  ������  �_����      D   ,  ������  ��  �  �  �  �����  ������      D   ,  ������  ��  �  �c  �  �c����  ������      D   ,  �?����  �?  �  Ƨ  �  Ƨ����  �?����      D   ,  Ǘ����  Ǘ  �  ��  �  ������  Ǘ����      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �����2  ������  ������  �����2  �����2      D   ,  ����2  �����  � ����  � ���2  ����2      D   ,  �h���2  �h����  �N����  �N���2  �h���2      D   ,  �����2  ������  ������  �����2  �����2      D   ,  ����2  �����  ������  �����2  ����2      D   ,  �R���2  �R����  �8����  �8���2  �R���2      D   ,  �����2  ������  ������  �����2  �����2      D   ,  �����2  ������  ������  �����2  �����2      D   ,  �<���2  �<����  �"����  �"���2  �<���2      D   ,  Ŋ���2  Ŋ����  �p����  �p���2  Ŋ���2      D   ,  �����2  ������  Ⱦ����  Ⱦ���2  �����2      D   ,  �  �  �  �  �   �  �   �  �  �      D   ,  �h  �  �h  �  �N  �  �N  �  �h  �      D   ,  ������  ��  �  �7  �  �7����  ������      D   ,  �&  �  �&  �  �  �  �  �  �&  �      D   ,  �t  �  �t  �  �Z  �  �Z  �  �t  �      D   ,  ��  �  ��  �  Ϩ  �  Ϩ  �  ��  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  �&���2  �&����  �����  ����2  �&���2      D   ,  �t���2  �t����  �Z����  �Z���2  �t���2      D   ,  �����2  ������  Ϩ����  Ϩ���2  �����2      D   ,  ����2  �����  ������  �����2  ����2      D   ,  �3����  �3  �  ͛  �  ͛����  �3����      D   ,  �w����  �w  �  ��  �  ������  �w����      D   ,  |�  �  |�  
�  ~'  
�  ~'  �  |�  �      D   ,  ��  &   ��  '�  ��  '�  ��  &   ��  &       D   ,  �M  &   �M  '�  ��  '�  ��  &   �M  &       D   ,  ��  &   ��  '�  �!  '�  �!  &   ��  &       D   ,  ��  &   ��  '�  �o  '�  �o  &   ��  &       D   ,  �7  &   �7  '�  ��  '�  ��  &   �7  &       D   ,  ��  &   ��  '�  �  '�  �  &   ��  &       D   ,  ��  &   ��  '�  �Y  '�  �Y  &   ��  &       D   ,  �!  &   �!  '�  ��  '�  ��  &   �!  &       D   ,  �o  &   �o  '�  ��  '�  ��  &   �o  &       D   ,  ��  &   ��  '�  �C  '�  �C  &   ��  &       D   ,  �  &   �  '�  ��  '�  ��  &   �  &       D   ,  �Y  &   �Y  '�  ��  '�  ��  &   �Y  &       D   ,  ��  &   ��  '�  �-  '�  �-  &   ��  &       D   ,  ��  &   ��  '�  �{  '�  �{  &   ��  &       D   ,  ��  &   ��  '�  �7  '�  �7  &   ��  &       D   ,  ��  &   ��  '�  �=  '�  �=  &   ��  &       D   ,  �  &   �  '�  ��  '�  ��  &   �  &       D   ,  �S  &   �S  '�  ��  '�  ��  &   �S  &       D   ,  ��  &   ��  '�  �'  '�  �'  &   ��  &       D   ,  ��  �  ��  5  ��  5  ��  �  ��  �      D   ,  ��  �  ��  5  ��  5  ��  �  ��  �      D   ,  �!  �  �!  5  �%  5  �%  �  �!  �      D   ,  �  '�  �  '�  ��  '�  ��  '�  �  '�      D   ,  ��  '�  ��  '�  ��  '�  ��  '�  ��  '�      D   ,  �  '�  �  '�  �=  '�  �=  '�  �  '�      D   ,  �i  '�  �i  '�  ��  '�  ��  '�  �i  '�      D   ,  ��  '�  ��  '�  ��  '�  ��  '�  ��  '�      D   ,  �  '�  �  '�  �'  '�  �'  '�  �  '�      D   ,  �S  '�  �S  '�  �u  '�  �u  '�  �S  '�      D   ,  ��  '�  ��  '�  ��  '�  ��  '�  ��  '�      D   ,  ��  '�  ��  '�  �  '�  �  '�  ��  '�      D   ,  �=  '�  �=  '�  �_  '�  �_  '�  �=  '�      D   ,  ��  '�  ��  '�  ��  '�  ��  '�  ��  '�      D   ,  ��  '�  ��  '�  ��  '�  ��  '�  ��  '�      D   ,  �'  '�  �'  '�  �I  '�  �I  '�  �'  '�      D   ,  ��  (�  ��  4?  �>  4?  �>  (�  ��  (�      D   ,  ��  '�  ��  '�  �  '�  �  '�  ��  '�      D   ,  �7  '�  �7  '�  �Y  '�  �Y  '�  �7  '�      D   ,  ��  '�  ��  '�  ��  '�  ��  '�  ��  '�      D   ,  ��  '�  ��  '�  ��  '�  ��  '�  ��  '�      D   ,  ~	  �  ~	  5    5    �  ~	  �      D   ,  ��  �  ��  5  ��  5  ��  �  ��  �      D   ,  �A  �  �A  5  �E  5  �E  �  �A  �      D   ,  ��  �  ��  5  ��  5  ��  �  ��  �      D   ,  �y  �  �y  5  �}  5  �}  �  �y  �      D   ,  �  �  �  5  �  5  �  �  �  �      D   ,  ��  �  ��  5  ��  5  ��  �  ��  �      D   ,  ~	  3  ~	  �    �    3  ~	  3      D   ,  ��  3  ��  �  ��  �  ��  3  ��  3      D   ,  �A  3  �A  �  �E  �  �E  3  �A  3      D   ,  ��  3  ��  �  ��  �  ��  3  ��  3      D   ,  �y  3  �y  �  �}  �  �}  3  �y  3      D   ,  �  3  �  �  �  �  �  3  �  3      D   ,  ��  3  ��  �  ��  �  ��  3  ��  3      D   ,  �M  3  �M  �  �Q  �  �Q  3  �M  3      D   ,  ��  3  ��  �  ��  �  ��  3  ��  3      D   ,  ��  L  ��  �  ��  �  ��  L  ��  L      D   ,  �!  `  �!  �  �%  �  �%  `  �!  `      D   ,  �M  �  �M  5  �Q  5  �Q  �  �M  �      D   ,  s  &   s  '�  t�  '�  t�  &   s  &       D   ,  uS  &   uS  '�  v�  '�  v�  &   uS  &       D   ,  w�  &   w�  '�  y'  '�  y'  &   w�  &       D   ,  y�  &   y�  '�  {u  '�  {u  &   y�  &       D   ,  Y�  &   Y�  '�  [1  '�  [1  &   Y�  &       D   ,  [�  &   [�  '�  ]  '�  ]  &   [�  &       D   ,  ^G  &   ^G  '�  _�  '�  _�  &   ^G  &       D   ,  `�  &   `�  '�  b  '�  b  &   `�  &       D   ,  b�  &   b�  '�  di  '�  di  &   b�  &       D   ,  e1  &   e1  '�  f�  '�  f�  &   e1  &       D   ,  g  &   g  '�  i  '�  i  &   g  &       D   ,  i�  &   i�  '�  kS  '�  kS  &   i�  &       D   ,  ]�  �  ]�  5  ^�  5  ^�  �  ]�  �      D   ,  ba  �  ba  5  ce  5  ce  �  ba  �      D   ,  f�  �  f�  5  h  5  h  �  f�  �      D   ,  p5  �  p5  5  q9  5  q9  �  p5  �      D   ,  t�  �  t�  5  u�  5  u�  �  t�  �      D   ,  ym  �  ym  5  zq  5  zq  �  ym  �      D   ,  k�  �  k�  5  l�  5  l�  �  k�  �      D   ,  Y�  '�  Y�  '�  Z�  '�  Z�  '�  Y�  '�      D   ,  \+  '�  \+  '�  ]M  '�  ]M  '�  \+  '�      D   ,  ^y  '�  ^y  '�  _�  '�  _�  '�  ^y  '�      D   ,  `�  '�  `�  '�  a�  '�  a�  '�  `�  '�      D   ,  c  '�  c  '�  d7  '�  d7  '�  c  '�      D   ,  ec  '�  ec  '�  f�  '�  f�  '�  ec  '�      D   ,  ]�  G  ]�  �  ^�  �  ^�  G  ]�  G      D   ,  ba  G  ba  �  ce  �  ce  G  ba  G      D   ,  ]�  3  ]�  G  ce  G  ce  3  ]�  3      D   ,  f�  3  f�  �  h  �  h  3  f�  3      D   ,  k�  3  k�  �  l�  �  l�  3  k�  3      D   ,  p5  3  p5  �  q9  �  q9  3  p5  3      D   ,  t�  3  t�  �  u�  �  u�  3  t�  3      D   ,  ym  3  ym  �  zq  �  zq  3  ym  3      D   ,  g�  '�  g�  '�  h�  '�  h�  '�  g�  '�      D   ,  i�  '�  i�  '�  k!  '�  k!  '�  i�  '�      D   ,  lM  '�  lM  '�  mo  '�  mo  '�  lM  '�      D   ,  n�  '�  n�  '�  o�  '�  o�  '�  n�  '�      D   ,  p�  '�  p�  '�  r  '�  r  '�  p�  '�      D   ,  s7  '�  s7  '�  tY  '�  tY  '�  s7  '�      D   ,  u�  '�  u�  '�  v�  '�  v�  '�  u�  '�      D   ,  w�  '�  w�  '�  x�  '�  x�  '�  w�  '�      D   ,  z!  '�  z!  '�  {C  '�  {C  '�  z!  '�      D   ,  l  &   l  '�  m�  '�  m�  &   l  &       D   ,  ni  &   ni  '�  o�  '�  o�  &   ni  &       D   ,  p�  &   p�  '�  r=  '�  r=  &   p�  &       D   ,  cG  �  cG  
�  d�  
�  d�  �  cG  �      D   ,  e�  �  e�  
�  g  
�  g  �  e�  �      D   ,  g�  �  g�  
�  ii  
�  ii  �  g�  �      D   ,  j1  �  j1  
�  k�  
�  k�  �  j1  �      D   ,  l  �  l  
�  n  
�  n  �  l  �      D   ,  n�  �  n�  
�  pS  
�  pS  �  n�  �      D   ,  ]�����  ]�  �  ^�  �  ^�����  ]�����      D   ,  _�����  _�  �  a?  �  a?����  _�����      D   ,  b/����  b/  �  c�  �  c�����  b/����      D   ,  ds����  ds  �  e�  �  e�����  ds����      D   ,  f�����  f�  �  h3  �  h3����  f�����      D   ,  i����  i  �  jw  �  jw����  i����      D   ,  kg����  kg  �  l�  �  l�����  kg����      D   ,  m�����  m�  �  o  �  o����  m�����      D   ,  p����  p  �  qk  �  qk����  p����      D   ,  rG����  rG  �  s�  �  s�����  rG����      D   ,  t�����  t�  �  v  �  v����  t�����      D   ,  v�����  v�  �  xK  �  xK����  v�����      D   ,  y;����  y;  �  z�  �  z�����  y;����      D   ,  {����  {  �  |�  �  |�����  {����      D   ,  q  �  q  
�  r�  
�  r�  �  q  �      D   ,  si  �  si  
�  t�  
�  t�  �  si  �      D   ,  u�  �  u�  
�  w=  
�  w=  �  u�  �      D   ,  x  �  x  
�  y�  
�  y�  �  x  �      D   ,  zS  �  zS  
�  {�  
�  {�  �  zS  �      D   ,  k�  �  k�  �  l�  �  l�  �  k�  �      D   ,  m�  �  m�  �  n�  �  n�  �  m�  �      D   ,  pD  �  pD  �  q*  �  q*  �  pD  �      D   ,  r�  �  r�  �  sx  �  sx  �  r�  �      D   ,  ]�  �  ]�  >  ^�  >  ^�  �  ]�  �      D   ,  `"  �  `"  >  a  >  a  �  `"  �      D   ,  bp  �  bp  >  cV  >  cV  �  bp  �      D   ,  d�  �  d�  >  e�  >  e�  �  d�  �      D   ,  g  �  g  >  g�  >  g�  �  g  �      D   ,  iZ  �  iZ  >  j@  >  j@  �  iZ  �      D   ,  ]����2  ]�����  ^�����  ^����2  ]����2      D   ,  `"���2  `"����  a����  a���2  `"���2      D   ,  bp���2  bp����  cV����  cV���2  bp���2      D   ,  d����2  d�����  e�����  e����2  d����2      D   ,  g���2  g����  g�����  g����2  g���2      D   ,  iZ���2  iZ����  j@����  j@���2  iZ���2      D   ,  k����2  k�����  l�����  l����2  k����2      D   ,  m����2  m�����  n�����  n����2  m����2      D   ,  pD���2  pD����  q*����  q*���2  pD���2      D   ,  r����2  r�����  sx����  sx���2  r����2      D   ,  t����2  t�����  u�����  u����2  t����2      D   ,  w.���2  w.����  x����  x���2  w.���2      D   ,  y|���2  y|����  zb����  zb���2  y|���2      D   ,  {����2  {�����  |�����  |����2  {����2      D   ,  k�  �  k�  >  l�  >  l�  �  k�  �      D   ,  m�  �  m�  >  n�  >  n�  �  m�  �      D   ,  pD  �  pD  >  q*  >  q*  �  pD  �      D   ,  r�  �  r�  >  sx  >  sx  �  r�  �      D   ,  t�  �  t�  >  u�  >  u�  �  t�  �      D   ,  w.  �  w.  >  x  >  x  �  w.  �      D   ,  y|  �  y|  >  zb  >  zb  �  y|  �      D   ,  {�  �  {�  >  |�  >  |�  �  {�  �      D   ,  t�  �  t�  �  u�  �  u�  �  t�  �      D   ,  w.  �  w.  �  x  �  x  �  w.  �      D   ,  y|  �  y|  �  zb  �  zb  �  y|  �      D   ,  {�  �  {�  �  |�  �  |�  �  {�  �      D   ,  v�  �  v�  �  xK  �  xK  �  v�  �      D   ,  y;  �  y;  �  z�  �  z�  �  y;  �      D   ,  {  �  {  �  |�  �  |�  �  {  �      D   ,  i  �  i  �  jw  �  jw  �  i  �      D   ,  kg  �  kg  �  l�  �  l�  �  kg  �      D   ,  m�  �  m�  �  o  �  o  �  m�  �      D   ,  p  �  p  �  qk  �  qk  �  p  �      D   ,  rG  �  rG  �  s�  �  s�  �  rG  �      D   ,  ]�  �  ]�  �  ^�  �  ^�  �  ]�  �      D   ,  `"  �  `"  �  a  �  a  �  `"  �      D   ,  bp  �  bp  �  cV  �  cV  �  bp  �      D   ,  d�  �  d�  �  e�  �  e�  �  d�  �      D   ,  g  �  g  �  g�  �  g�  �  g  �      D   ,  iZ  �  iZ  �  j@  �  j@  �  iZ  �      D   ,  k�  �  k�  �  l�  �  l�  �  k�  �      D   ,  m�  �  m�  �  n�  �  n�  �  m�  �      D   ,  pD  �  pD  �  q*  �  q*  �  pD  �      D   ,  r�  �  r�  �  sx  �  sx  �  r�  �      D   ,  t�  �  t�  �  u�  �  u�  �  t�  �      D   ,  w.  �  w.  �  x  �  x  �  w.  �      D   ,  y|  �  y|  �  zb  �  zb  �  y|  �      D   ,  {�  �  {�  �  |�  �  |�  �  {�  �      D   ,  t�  �  t�  �  v  �  v  �  t�  �      D   ,  ]�  �  ]�  �  ^�  �  ^�  �  ]�  �      D   ,  `"  �  `"  �  a  �  a  �  `"  �      D   ,  bp  �  bp  �  cV  �  cV  �  bp  �      D   ,  d�  �  d�  �  e�  �  e�  �  d�  �      D   ,  g  �  g  �  g�  �  g�  �  g  �      D   ,  iZ  �  iZ  �  j@  �  j@  �  iZ  �      D   ,  ^�  �  ^�  
�  `1  
�  `1  �  ^�  �      D   ,  `�  �  `�  
�  b  
�  b  �  `�  �      D   ,  ]�  �  ]�  �  ^�  �  ^�  �  ]�  �      D   ,  _�  �  _�  �  a?  �  a?  �  _�  �      D   ,  b/  �  b/  �  c�  �  c�  �  b/  �      D   ,  ds  �  ds  �  e�  �  e�  �  ds  �      D   ,  f�  �  f�  �  h3  �  h3  �  f�  �      D   ,  �'  �  �'  
�  ��  
�  ��  �  �'  �      D   ,  �u  �  �u  
�  ��  
�  ��  �  �u  �      D   ,  ��  �  ��  
�  �I  
�  �I  �  ��  �      D   ,  �  �  �  
�  ��  
�  ��  �  �  �      D   ,  �_  �  �_  
�  ��  
�  ��  �  �_  �      D   ,  ��  �  ��  
�  �3  
�  �3  �  ��  �      D   ,  ��  �  ��  
�  ��  
�  ��  �  ��  �      D   ,  �I  �  �I  
�  ��  
�  ��  �  �I  �      D   ,  ��  �  ��  
�  �  
�  �  �  ��  �      D   ,  ��  �  ��  
�  �k  
�  �k  �  ��  �      D   ,  �3  �  �3  
�  ��  
�  ��  �  �3  �      D   ,  ��  �  ��  
�  �  
�  �  �  ��  �      D   ,  ��  �  ��  
�  �U  
�  �U  �  ��  �      D   ,  �  �  �  
�  ��  
�  ��  �  �  �      D   ,  �k  �  �k  
�  ��  
�  ��  �  �k  �      D   ,  ��  �  ��  
�  �?  
�  �?  �  ��  �      D   ,  �  �  �  
�  ��  
�  ��  �  �  �      D   ,  ~�  �  ~�  
�  �u  
�  �u  �  ~�  �      D   ,  �=  �  �=  
�  ��  
�  ��  �  �=  �      D   ,  ��  �  ��  
�  �  
�  �  �  ��  �      D   ,  ��  �  ��  
�  �_  
�  �_  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �F  �  �F  �  �,  �  �,  �  �F  �      D   ,  ��  �  ��  �  �z  �  �z  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �0  �  �0  �  �  �  �  �  �0  �      D   ,  �~  �  �~  �  �d  �  �d  �  �~  �      D   ,  �'  �  �'  �  ��  �  ��  �  �'  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  ��  �  ��  �  �+  �  �+  �  ��  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  �_  �  �_  �  ��  �  ��  �  �_  �      D   ,  ��  �  ��  �  �  �  �  �  ��  �      D   ,  ��  �  ��  �  �c  �  �c  �  ��  �      D   ,  �S  �  �S  �  ��  �  ��  �  �S  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  ��  �  ��  �  �W  �  �W  �  ��  �      D   ,  �r  �  �r  >  �X  >  �X  �  �r  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  �  �  �  >  ��  >  ��  �  �  �      D   ,  �\  �  �\  >  �B  >  �B  �  �\  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  �F  �  �F  >  �,  >  �,  �  �F  �      D   ,  ��  �  ��  >  �z  >  �z  �  ��  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  �0  �  �0  >  �  >  �  �  �0  �      D   ,  �~  �  �~  >  �d  >  �d  �  �~  �      D   ,  �3  �  �3  �  ��  �  ��  �  �3  �      D   ,  �r  �  �r  �  �X  �  �X  �  �r  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  �\  �  �\  �  �B  �  �B  �  �\  �      D   ,  ��  �  ��  >  �n  >  �n  �  ��  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  �$  �  �$  >  �
  >  �
  �  �$  �      D   ,  ��  �  ��  �  �n  �  �n  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  ��  �  ��  �  �W  �  �W  �  ��  �      D   ,  �G  �  �G  �  ��  �  ��  �  �G  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  ��  �  ��  �  �K  �  �K  �  ��  �      D   ,  �$  �  �$  �  �
  �  �
  �  �$  �      D   ,  �:  �  �:  �  �   �  �   �  �:  �      D   ,  ~  �  ~  >  ~�  >  ~�  �  ~  �      D   ,  �f  �  �f  >  �L  >  �L  �  �f  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  �  �  �  >  ��  >  ��  �  �  �      D   ,  }�  �  }�  �  ?  �  ?  �  }�  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  �s  �  �s  �  ��  �  ��  �  �s  �      D   ,  ��  �  ��  �  �  �  �  �  ��  �      D   ,  �  �  �  �  �w  �  �w  �  �  �      D   ,  �S  �  �S  �  ��  �  ��  �  �S  �      D   ,  ��  �  ��  �  �  �  �  �  ��  �      D   ,  ~  �  ~  �  ~�  �  ~�  �  ~  �      D   ,  �f  �  �f  �  �L  �  �L  �  �f  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  �P  �  �P  �  �6  �  �6  �  �P  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �P  �  �P  >  �6  >  �6  �  �P  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  ��  �  ��  >  ��  >  ��  �  ��  �      D   ,  �:  �  �:  >  �   >  �   �  �:  �      D   ,  ������  ��  �  ��  �  ������  ������      D   ,  ������  ��  �  �K  �  �K����  ������      D   ,  }�����  }�  �  ?  �  ?����  }�����      D   ,  �����  �  �  ��  �  ������  �����      D   ,  �s����  �s  �  ��  �  ������  �s����      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  �P  �  �P  �  �6  �  �6  �  �P  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �:  �  �:  �  �   �  �   �  �:  �      D   ,  ��  �  ��  �  �n  �  �n  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �$  �  �$  �  �
  �  �
  �  �$  �      D   ,  ~  �  ~  �  ~�  �  ~�  �  ~  �      D   ,  ������  ��  �  �  �  �����  ������      D   ,  �����  �  �  �w  �  �w����  �����      D   ,  �S����  �S  �  ��  �  ������  �S����      D   ,  ������  ��  �  �  �  �����  ������      D   ,  ~���2  ~����  ~�����  ~����2  ~���2      D   ,  �f���2  �f����  �L����  �L���2  �f���2      D   ,  �����2  ������  ������  �����2  �����2      D   ,  ����2  �����  ������  �����2  ����2      D   ,  �P���2  �P����  �6����  �6���2  �P���2      D   ,  �����2  ������  ������  �����2  �����2      D   ,  �f  �  �f  �  �L  �  �L  �  �f  �      D   ,  �����2  ������  ������  �����2  �����2      D   ,  �:���2  �:����  � ����  � ���2  �:���2      D   ,  �����2  ������  �n����  �n���2  �����2      D   ,  �����2  ������  ������  �����2  �����2      D   ,  �$���2  �$����  �
����  �
���2  �$���2      D   ,  ������  ��  �  �W  �  �W����  ������      D   ,  �G����  �G  �  ��  �  ������  �G����      D   ,  �����2  ������  ������  �����2  �����2      D   ,  �����2  ������  ������  �����2  �����2      D   ,  �F���2  �F����  �,����  �,���2  �F���2      D   ,  �r  �  �r  �  �X  �  �X  �  �r  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �  �  �  �  ��  �  ��  �  �  �      D   ,  �\  �  �\  �  �B  �  �B  �  �\  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �F  �  �F  �  �,  �  �,  �  �F  �      D   ,  ��  �  ��  �  �z  �  �z  �  ��  �      D   ,  ��  �  ��  �  ��  �  ��  �  ��  �      D   ,  �0  �  �0  �  �  �  �  �  �0  �      D   ,  �~  �  �~  �  �d  �  �d  �  �~  �      D   ,  �����2  ������  �z����  �z���2  �����2      D   ,  �����2  ������  ������  �����2  �����2      D   ,  �0���2  �0����  �����  ����2  �0���2      D   ,  �~���2  �~����  �d����  �d���2  �~���2      D   ,  �S����  �S  �  ��  �  ������  �S����      D   ,  ������  ��  �  ��  �  ������  ������      D   ,  ������  ��  �  �W  �  �W����  ������      D   ,  �3����  �3  �  ��  �  ������  �3����      D   ,  �'����  �'  �  ��  �  ������  �'����      D   ,  �����  �  �  ��  �  ������  �����      D   ,  ������  ��  �  �+  �  �+����  ������      D   ,  �����  �  �  ��  �  ������  �����      D   ,  �_����  �_  �  ��  �  ������  �_����      D   ,  ������  ��  �  �  �  �����  ������      D   ,  ������  ��  �  �c  �  �c����  ������      D   ,  �r���2  �r����  �X����  �X���2  �r���2      D   ,  �����2  ������  ������  �����2  �����2      D   ,  ����2  �����  ������  �����2  ����2      D   ,  �\���2  �\����  �B����  �B���2  �\���2      D   ,  |���߭  |����  ~'���  ~'��߭  |���߭      D   ,  ]���ӌ  ]����|  ^����|  ^���ӌ  ]���ӌ      D   ,  _���ӌ  _����|  a?���|  a?��ӌ  _���ӌ      D   ,  b/��ӌ  b/���|  c����|  c���ӌ  b/��ӌ      D   ,  ds��ӌ  ds���|  e����|  e���ӌ  ds��ӌ      D   ,  f���ӌ  f����|  h3���|  h3��ӌ  f���ӌ      D   ,  i��ӌ  i���|  jw���|  jw��ӌ  i��ӌ      D   ,  kg��ӌ  kg���|  l����|  l���ӌ  kg��ӌ      D   ,  m���ӌ  m����|  o���|  o��ӌ  m���ӌ      D   ,  p��ӌ  p���|  qk���|  qk��ӌ  p��ӌ      D   ,  rG��ӌ  rG���|  s����|  s���ӌ  rG��ӌ      D   ,  t���ӌ  t����|  v���|  v��ӌ  t���ӌ      D   ,  v���ӌ  v����|  xK���|  xK��ӌ  v���ӌ      D   ,  y;��ӌ  y;���|  z����|  z���ӌ  y;��ӌ      D   ,  {��ӌ  {���|  |����|  |���ӌ  {��ӌ      D   ,  }���ӌ  }����|  ?���|  ?��ӌ  }���ӌ      D   ,  ���ӌ  ����|  �����|  ����ӌ  ���ӌ      D   ,  �s��ӌ  �s���|  �����|  ����ӌ  �s��ӌ      D   ,  ����ӌ  �����|  ����|  ���ӌ  ����ӌ      D   ,  ���ӌ  ����|  �w���|  �w��ӌ  ���ӌ      D   ,  �S��ӌ  �S���|  �����|  ����ӌ  �S��ӌ      D   ,  ����ӌ  �����|  ����|  ���ӌ  ����ӌ      D   ,  ����ӌ  �����|  �W���|  �W��ӌ  ����ӌ      D   ,  �G��ӌ  �G���|  �����|  ����ӌ  �G��ӌ      D   ,  ����ӌ  �����|  �����|  ����ӌ  ����ӌ      D   ,  ����ӌ  �����|  �K���|  �K��ӌ  ����ӌ      D   ,  �'��ӌ  �'���|  �����|  ����ӌ  �'��ӌ      D   ,  ���ӌ  ����|  �����|  ����ӌ  ���ӌ      D   ,  ����ӌ  �����|  �+���|  �+��ӌ  ����ӌ      D   ,  ���ӌ  ����|  �����|  ����ӌ  ���ӌ      D   ,  �_��ӌ  �_���|  �����|  ����ӌ  �_��ӌ      D   ,  ����ӌ  �����|  ����|  ���ӌ  ����ӌ      D   ,  ����ӌ  �����|  �c���|  �c��ӌ  ����ӌ      D   ,  �S��ӌ  �S���|  �����|  ����ӌ  �S��ӌ      D   ,  ����ӌ  �����|  �����|  ����ӌ  ����ӌ      D   ,  ����ӌ  �����|  �W���|  �W��ӌ  ����ӌ      D   ,  �3��ӌ  �3���|  �����|  ����ӌ  �3��ӌ      D   ,  �����  �����  �w����  �w����  �����      D   ,  ����߭  �����  �����  ����߭  ����߭      D   ,  �S����  �S����  ������  ������  �S����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �W����  �W����  ������      D   ,  �G����  �G����  ������  ������  �G����      D   ,  ������  ������  ������  ������  ������      D   ,  ������  ������  �K����  �K����  ������      D   ,  �'����  �'����  ������  ������  �'����      D   ,  �����  �����  ������  ������  �����      D   ,  ������  ������  �+����  �+����  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �_����  �_����  ������  ������  �_����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �c����  �c����  ������      D   ,  �S����  �S����  ������  ������  �S����      D   ,  ������  ������  ������  ������  ������      D   ,  ������  ������  �W����  �W����  ������      D   ,  �3����  �3����  ������  ������  �3����      D   ,  }�����  }�����  ?����  ?����  }�����      D   ,  �����  �����  ������  ������  �����      D   ,  �s����  �s����  ������  ������  �s����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  �����4  �����4  ������  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �F����  �F���4  �,���4  �,����  �F����      D   ,  ������  ������  �\����  �\����  ������      D   ,  ������  �����4  �����4  ������  ������      D   ,  �N����  �N����  ������  ������  �N����      D   ,  �~����  �~���4  �d���4  �d����  �~����      D   ,  �r����  �r���4  �X���4  �X����  �r����      D   ,  ������  ������  ������  ������  ������      D   ,  �����  ����4  �����4  ������  �����      D   ,  �z����  �z����  �$����  �$����  �z����      D   ,  �n����  �n����  �����  �����  �n����      D   ,  ������  �����4  �����4  ������  ������      D   ,  �
����  �
����  ������  ������  �
����      D   ,  �:����  �:���4  � ���4  � ����  �:����      D   ,  ������  ������  �P����  �P����  ������      D   ,  ������  �����4  �����4  ������  ������      D   ,  �B����  �B����  ������  ������  �B����      D   ,  ~6����  ~6����  ~�����  ~�����  ~6����      D   ,  �f����  �f���4  �L���4  �L����  �f����      D   ,  ������  ������  �|����  �|����  ������      D   ,  �����  ����4  �����4  ������  �����      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �:���|  �:����  � ����  � ���|  �:���|      D   ,  �����|  ������  �n����  �n���|  �����|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �$���|  �$����  �
����  �
���|  �$���|      D   ,  �:���|  �:����  � ����  � ���|  �:���|      D   ,  �����|  ������  �n����  �n���|  �����|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �$���|  �$����  �
����  �
���|  �$���|      D   ,  �=��߭  �=���  �����  ����߭  �=��߭      D   ,  ����߭  �����  ����  ���߭  ����߭      D   ,  ����߭  �����  �_���  �_��߭  ����߭      D   ,  �'��߭  �'���  �����  ����߭  �'��߭      D   ,  �u��߭  �u���  �����  ����߭  �u��߭      D   ,  ����߭  �����  �I���  �I��߭  ����߭      D   ,  ���߭  ����  �����  ����߭  ���߭      D   ,  �_��߭  �_���  �����  ����߭  �_��߭      D   ,  ����߭  �����  �3���  �3��߭  ����߭      D   ,  ~���߭  ~����  �u���  �u��߭  ~���߭      D   ,  ~���|  ~����  ~�����  ~����|  ~���|      D   ,  �f���|  �f����  �L����  �L���|  �f���|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  ����|  �����  ������  �����|  ����|      D   ,  �P���|  �P����  �6����  �6���|  �P���|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  ~���|  ~����  ~�����  ~����|  ~���|      D   ,  �f���|  �f����  �L����  �L���|  �f���|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  ����|  �����  ������  �����|  ����|      D   ,  �P���|  �P����  �6����  �6���|  �P���|      D   ,  ����|  �����  ������  �����|  ����|      D   ,  �\���|  �\����  �B����  �B���|  �\���|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �F���|  �F����  �,����  �,���|  �F���|      D   ,  �����|  ������  �z����  �z���|  �����|      D   ,  �~���|  �~����  �d����  �d���|  �~���|      D   ,  �I��߭  �I���  �����  ����߭  �I��߭      D   ,  ����߭  �����  ����  ���߭  ����߭      D   ,  ����߭  �����  �k���  �k��߭  ����߭      D   ,  �3��߭  �3���  �����  ����߭  �3��߭      D   ,  ����߭  �����  ����  ���߭  ����߭      D   ,  ����߭  �����  �U���  �U��߭  ����߭      D   ,  ���߭  ����  �����  ����߭  ���߭      D   ,  �k��߭  �k���  �����  ����߭  �k��߭      D   ,  �r���|  �r����  �X����  �X���|  �r���|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  ����|  �����  ������  �����|  ����|      D   ,  �\���|  �\����  �B����  �B���|  �\���|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �F���|  �F����  �,����  �,���|  �F���|      D   ,  �����|  ������  �z����  �z���|  �����|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �0���|  �0����  �����  ����|  �0���|      D   ,  �~���|  �~����  �d����  �d���|  �~���|      D   ,  ����߭  �����  �?���  �?��߭  ����߭      D   ,  ���߭  ����  �����  ����߭  ���߭      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �0���|  �0����  �����  ����|  �0���|      D   ,  �r���|  �r����  �X����  �X���|  �r���|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  q��߭  q���  r����  r���߭  q��߭      D   ,  si��߭  si���  t����  t���߭  si��߭      D   ,  u���߭  u����  w=���  w=��߭  u���߭      D   ,  x��߭  x���  y����  y���߭  x��߭      D   ,  zS��߭  zS���  {����  {���߭  zS��߭      D   ,  pD���|  pD����  q*����  q*���|  pD���|      D   ,  r����|  r�����  sx����  sx���|  r����|      D   ,  t����|  t�����  u�����  u����|  t����|      D   ,  w.���|  w.����  x����  x���|  w.���|      D   ,  y|���|  y|����  zb����  zb���|  y|���|      D   ,  {����|  {�����  |�����  |����|  {����|      D   ,  ]����|  ]�����  ^�����  ^����|  ]����|      D   ,  `"���|  `"����  a����  a���|  `"���|      D   ,  bp���|  bp����  cV����  cV���|  bp���|      D   ,  d����|  d�����  e�����  e����|  d����|      D   ,  g���|  g����  g�����  g����|  g���|      D   ,  `"����  `"���4  a���4  a����  `"����      D   ,  bp����  bp���4  cV���4  cV����  bp����      D   ,  d�����  d����4  e����4  e�����  d�����      D   ,  g*����  g*����  g�����  g�����  g*����      D   ,  iZ����  iZ���4  j@���4  j@����  iZ����      D   ,  k�����  k�����  lp����  lp����  k�����      D   ,  m�����  m����4  n����4  n�����  m�����      D   ,  pb����  pb����  q����  q����  pb����      D   ,  r�����  r����4  sx���4  sx����  r�����      D   ,  t�����  t�����  u�����  u�����  t�����      D   ,  w.����  w.���4  x���4  x����  w.����      D   ,  y�����  y�����  zD����  zD����  y�����      D   ,  {�����  {����4  |����4  |�����  {�����      D   ,  iZ���|  iZ����  j@����  j@���|  iZ���|      D   ,  k����|  k�����  l�����  l����|  k����|      D   ,  m����|  m�����  n�����  n����|  m����|      D   ,  ^���߭  ^����  `1���  `1��߭  ^���߭      D   ,  `���߭  `����  b���  b��߭  `���߭      D   ,  cG��߭  cG���  d����  d���߭  cG��߭      D   ,  e���߭  e����  g���  g��߭  e���߭      D   ,  g���߭  g����  ii���  ii��߭  g���߭      D   ,  j1��߭  j1���  k����  k���߭  j1��߭      D   ,  l��߭  l���  n���  n��߭  l��߭      D   ,  n���߭  n����  pS���  pS��߭  n���߭      D   ,  ]�����  ]����4  ^����4  ^�����  ]�����      D   ,  ]����|  ]�����  ^�����  ^����|  ]����|      D   ,  `"���|  `"����  a����  a���|  `"���|      D   ,  bp���|  bp����  cV����  cV���|  bp���|      D   ,  d����|  d�����  e�����  e����|  d����|      D   ,  g���|  g����  g�����  g����|  g���|      D   ,  iZ���|  iZ����  j@����  j@���|  iZ���|      D   ,  k����|  k�����  l�����  l����|  k����|      D   ,  m����|  m�����  n�����  n����|  m����|      D   ,  pD���|  pD����  q*����  q*���|  pD���|      D   ,  r����|  r�����  sx����  sx���|  r����|      D   ,  ]�����  ]�����  ^�����  ^�����  ]�����      D   ,  _�����  _�����  a?����  a?����  _�����      D   ,  b/����  b/����  c�����  c�����  b/����      D   ,  ds����  ds����  e�����  e�����  ds����      D   ,  f�����  f�����  h3����  h3����  f�����      D   ,  i����  i����  jw����  jw����  i����      D   ,  kg����  kg����  l�����  l�����  kg����      D   ,  m�����  m�����  o����  o����  m�����      D   ,  p����  p����  qk����  qk����  p����      D   ,  rG����  rG����  s�����  s�����  rG����      D   ,  t�����  t�����  v����  v����  t�����      D   ,  v�����  v�����  xK����  xK����  v�����      D   ,  y;����  y;����  z�����  z�����  y;����      D   ,  {����  {����  |�����  |�����  {����      D   ,  t����|  t�����  u�����  u����|  t����|      D   ,  w.���|  w.����  x����  x���|  w.���|      D   ,  y|���|  y|����  zb����  zb���|  y|���|      D   ,  {����|  {�����  |�����  |����|  {����|      D   ,  t�����  t����*  u����*  u�����  t�����      D   ,  w.����  w.���*  x���*  x����  w.����      D   ,  y|����  y|���*  zb���*  zb����  y|����      D   ,  {�����  {����*  |����*  |�����  {�����      D   ,  `"���(  `"��ӌ  a��ӌ  a���(  `"���(      D   ,  bp���(  bp��ӌ  cV��ӌ  cV���(  bp���(      D   ,  d����(  d���ӌ  e���ӌ  e����(  d����(      D   ,  g���(  g��ӌ  g���ӌ  g����(  g���(      D   ,  iZ���(  iZ��ӌ  j@��ӌ  j@���(  iZ���(      D   ,  k����(  k���ӌ  l���ӌ  l����(  k����(      D   ,  m����(  m���ӌ  n���ӌ  n����(  m����(      D   ,  pD���(  pD��ӌ  q*��ӌ  q*���(  pD���(      D   ,  r����(  r���ӌ  sx��ӌ  sx���(  r����(      D   ,  t����(  t���ӌ  u���ӌ  u����(  t����(      D   ,  w.���(  w.��ӌ  x��ӌ  x���(  w.���(      D   ,  y|���(  y|��ӌ  zb��ӌ  zb���(  y|���(      D   ,  {����(  {���ӌ  |���ӌ  |����(  {����(      D   ,  ]����(  ]���ӌ  ^���ӌ  ^����(  ]����(      D   ,  ]�����  ]����*  ^����*  ^�����  ]�����      D   ,  `"����  `"���*  a���*  a����  `"����      D   ,  bp����  bp���*  cV���*  cV����  bp����      D   ,  d�����  d����*  e����*  e�����  d�����      D   ,  g����  g���*  g����*  g�����  g����      D   ,  iZ����  iZ���*  j@���*  j@����  iZ����      D   ,  k�����  k����*  l����*  l�����  k�����      D   ,  m�����  m����*  n����*  n�����  m�����      D   ,  pD����  pD���*  q*���*  q*����  pD����      D   ,  r�����  r����*  sx���*  sx����  r�����      D   ,  �f���(  �f��ӌ  �L��ӌ  �L���(  �f���(      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  ����(  ���ӌ  ����ӌ  �����(  ����(      D   ,  �P���(  �P��ӌ  �6��ӌ  �6���(  �P���(      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  �:���(  �:��ӌ  � ��ӌ  � ���(  �:���(      D   ,  �����(  ����ӌ  �n��ӌ  �n���(  �����(      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  �$���(  �$��ӌ  �
��ӌ  �
���(  �$���(      D   ,  �r���(  �r��ӌ  �X��ӌ  �X���(  �r���(      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  ����(  ���ӌ  ����ӌ  �����(  ����(      D   ,  �\���(  �\��ӌ  �B��ӌ  �B���(  �\���(      D   ,  ~����  ~���*  ~����*  ~�����  ~����      D   ,  �f����  �f���*  �L���*  �L����  �f����      D   ,  ������  �����*  �����*  ������  ������      D   ,  �����  ����*  �����*  ������  �����      D   ,  �P����  �P���*  �6���*  �6����  �P����      D   ,  ������  �����*  �����*  ������  ������      D   ,  ������  �����*  �����*  ������  ������      D   ,  �:����  �:���*  � ���*  � ����  �:����      D   ,  ������  �����*  �n���*  �n����  ������      D   ,  ������  �����*  �����*  ������  ������      D   ,  �$����  �$���*  �
���*  �
����  �$����      D   ,  �r����  �r���*  �X���*  �X����  �r����      D   ,  ������  �����*  �����*  ������  ������      D   ,  �����  ����*  �����*  ������  �����      D   ,  �\����  �\���*  �B���*  �B����  �\����      D   ,  ������  �����*  �����*  ������  ������      D   ,  ������  �����*  �����*  ������  ������      D   ,  �F����  �F���*  �,���*  �,����  �F����      D   ,  ������  �����*  �z���*  �z����  ������      D   ,  ������  �����*  �����*  ������  ������      D   ,  �0����  �0���*  ����*  �����  �0����      D   ,  �~����  �~���*  �d���*  �d����  �~����      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  �F���(  �F��ӌ  �,��ӌ  �,���(  �F���(      D   ,  �����(  ����ӌ  �z��ӌ  �z���(  �����(      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  �0���(  �0��ӌ  ���ӌ  ����(  �0���(      D   ,  �~���(  �~��ӌ  �d��ӌ  �d���(  �~���(      D   ,  ~���(  ~��ӌ  ~���ӌ  ~����(  ~���(      D   ,  ����ӌ  �����|  �����|  ����ӌ  ����ӌ      D   ,  ����ӌ  �����|  �7���|  �7��ӌ  ����ӌ      D   ,  �'��ӌ  �'���|  �����|  ����ӌ  �'��ӌ      D   ,  �k��ӌ  �k���|  �����|  ����ӌ  �k��ӌ      D   ,  ����ӌ  �����|  �+���|  �+��ӌ  ����ӌ      D   ,  ���ӌ  ����|  �o���|  �o��ӌ  ���ӌ      D   ,  �_��ӌ  �_���|  �����|  ����ӌ  �_��ӌ      D   ,  ����ӌ  �����|  ����|  ���ӌ  ����ӌ      D   ,  ����ӌ  �����|  �c���|  �c��ӌ  ����ӌ      D   ,  �?��ӌ  �?���|  Ƨ���|  Ƨ��ӌ  �?��ӌ      D   ,  Ǘ��ӌ  Ǘ���|  �����|  ����ӌ  Ǘ��ӌ      D   ,  ����ӌ  �����|  �C���|  �C��ӌ  ����ӌ      D   ,  �3��ӌ  �3���|  ͛���|  ͛��ӌ  �3��ӌ      D   ,  �w��ӌ  �w���|  �����|  ����ӌ  �w��ӌ      D   ,  ����ӌ  �����|  �7���|  �7��ӌ  ����ӌ      D   ,  ����߭  �����  �a���  �a��߭  ����߭      D   ,  �)��߭  �)���  �����  ����߭  �)��߭      D   ,  �w��߭  �w���  �����  ����߭  �w��߭      D   ,  ����߭  �����  �K���  �K��߭  ����߭      D   ,  ���߭  ����  ř���  ř��߭  ���߭      D   ,  �a��߭  �a���  �����  ����߭  �a��߭      D   ,  ȯ��߭  ȯ���  �5���  �5��߭  ȯ��߭      D   ,  ����߭  �����  ̃���  ̃��߭  ����߭      D   ,  �K��߭  �K���  �����  ����߭  �K��߭      D   ,  ϙ��߭  ϙ���  ����  ���߭  ϙ��߭      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �<���|  �<����  �"����  �"���|  �<���|      D   ,  Ŋ���|  Ŋ����  �p����  �p���|  Ŋ���|      D   ,  �����|  ������  Ⱦ����  Ⱦ���|  �����|      D   ,  �&���|  �&����  �����  ����|  �&���|      D   ,  �t���|  �t����  �Z����  �Z���|  �t���|      D   ,  �����|  ������  Ϩ����  Ϩ���|  �����|      D   ,  ����|  �����  ������  �����|  ����|      D   ,  ̒����  ̒����  �<����  �<����  ̒����      D   ,  ������  �����4  Ϩ���4  Ϩ����  ������      D   ,  �.����  �.����  ������  ������  �.����      D   ,  ������  ������  ������  ������  ������      D   ,  �����|  ������  Ϩ����  Ϩ���|  �����|      D   ,  ����|  �����  ������  �����|  ����|      D   ,  Ŋ����  Ŋ���4  �p���4  �p����  Ŋ����      D   ,  ������  ������  Ƞ����  Ƞ����  ������      D   ,  �&����  �&���4  ����4  �����  �&����      D   ,  �����|  ������  ������  �����|  �����|      D   ,  ����|  �����  � ����  � ���|  ����|      D   ,  �h���|  �h����  �N����  �N���|  �h���|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  ����|  �����  ������  �����|  ����|      D   ,  �R���|  �R����  �8����  �8���|  �R���|      D   ,  ����߭  �����  �)���  �)��߭  ����߭      D   ,  ����߭  �����  �w���  �w��߭  ����߭      D   ,  �?��߭  �?���  �����  ����߭  �?��߭      D   ,  ����߭  �����  ����  ���߭  ����߭      D   ,  �����  ����4  � ���4  � ����  �����      D   ,  ������  ������  �0����  �0����  ������      D   ,  ������  �����4  �����4  ������  ������      D   ,  �"����  �"����  ������  ������  �"����      D   ,  �R����  �R���4  �8���4  �8����  �R����      D   ,  ������  ������  ������  ������  ������      D   ,  ������  ������  �7����  �7����  ������      D   ,  �'����  �'����  ������  ������  �'����      D   ,  �k����  �k����  ������  ������  �k����      D   ,  ������  ������  �+����  �+����  ������      D   ,  �����  �����  �o����  �o����  �����      D   ,  �_����  �_����  ������  ������  �_����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �c����  �c����  ������      D   ,  �?����  �?����  Ƨ����  Ƨ����  �?����      D   ,  Ǘ����  Ǘ����  ������  ������  Ǘ����      D   ,  ������  ������  �C����  �C����  ������      D   ,  �3����  �3����  ͛����  ͛����  �3����      D   ,  �w����  �w����  ������  ������  �w����      D   ,  ������  ������  �7����  �7����  ������      D   ,  ������  ������  �h����  �h����  ������      D   ,  ������  �����4  �����4  ������  ������      D   ,  �Z����  �Z����  �����  �����  �Z����      D   ,  �����|  ������  ������  �����|  �����|      D   ,  ����|  �����  � ����  � ���|  ����|      D   ,  �h���|  �h����  �N����  �N���|  �h���|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  ����|  �����  ������  �����|  ����|      D   ,  �R���|  �R����  �8����  �8���|  �R���|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �����|  ������  ������  �����|  �����|      D   ,  �<���|  �<����  �"����  �"���|  �<���|      D   ,  Ŋ���|  Ŋ����  �p����  �p���|  Ŋ���|      D   ,  �����|  ������  Ⱦ����  Ⱦ���|  �����|      D   ,  �&���|  �&����  �����  ����|  �&���|      D   ,  �t���|  �t����  �Z����  �Z���|  �t���|      D   ,  ������  �����*  �����*  ������  ������      D   ,  �<����  �<���*  �"���*  �"����  �<����      D   ,  Ŋ����  Ŋ���*  �p���*  �p����  Ŋ����      D   ,  ������  �����*  Ⱦ���*  Ⱦ����  ������      D   ,  �&����  �&���*  ����*  �����  �&����      D   ,  �t����  �t���*  �Z���*  �Z����  �t����      D   ,  ������  �����*  Ϩ���*  Ϩ����  ������      D   ,  �����  ����*  �����*  ������  �����      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  �<���(  �<��ӌ  �"��ӌ  �"���(  �<���(      D   ,  Ŋ���(  Ŋ��ӌ  �p��ӌ  �p���(  Ŋ���(      D   ,  �����(  ����ӌ  Ⱦ��ӌ  Ⱦ���(  �����(      D   ,  �&���(  �&��ӌ  ���ӌ  ����(  �&���(      D   ,  �t���(  �t��ӌ  �Z��ӌ  �Z���(  �t���(      D   ,  �����(  ����ӌ  Ϩ��ӌ  Ϩ���(  �����(      D   ,  ����(  ���ӌ  ����ӌ  �����(  ����(      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  ����(  ���ӌ  � ��ӌ  � ���(  ����(      D   ,  �h���(  �h��ӌ  �N��ӌ  �N���(  �h���(      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  ����(  ���ӌ  ����ӌ  �����(  ����(      D   ,  �R���(  �R��ӌ  �8��ӌ  �8���(  �R���(      D   ,  �����(  ����ӌ  ����ӌ  �����(  �����(      D   ,  ������  �����*  �����*  ������  ������      D   ,  �����  ����*  � ���*  � ����  �����      D   ,  �h����  �h���*  �N���*  �N����  �h����      D   ,  ������  �����*  �����*  ������  ������      D   ,  �����  ����*  �����*  ������  �����      D   ,  �R����  �R���*  �8���*  �8����  �R����      D   ,  ������  �����*  �����*  ������  ������      D   ,  �U����  �U����  ������  ������  �U����      D   ,  \�����  \�����  �����  �����  \�����      D   ,  �U����  �U����  ������  ������  �U����      D   ,  ]����x  ]����h  ^����h  ^����x  ]����x      D   ,  _����x  _����h  aS���h  aS���x  _����x      D   ,  b/���x  b/���h  c����h  c����x  b/���x      D   ,  d����x  d����h  e����h  e����x  d����x      D   ,  f����x  f����h  h3���h  h3���x  f����x      D   ,  i#���x  i#���h  j����h  j����x  i#���x      D   ,  kg���x  kg���h  l����h  l����x  kg���x      D   ,  m����x  m����h  o'���h  o'���x  m����x      D   ,  p���x  p���h  qk���h  qk���x  p���x      D   ,  r[���x  r[���h  s����h  s����x  r[���x      D   ,  t����x  t����h  v���h  v���x  t����x      D   ,  v����x  v����h  x_���h  x_���x  v����x      D   ,  y;���x  y;���h  z����h  z����x  y;���x      D   ,  {����x  {����h  |����h  |����x  {����x      D   ,  }����x  }����h  ?���h  ?���x  }����x      D   ,  �/���x  �/���h  �����h  �����x  �/���x      D   ,  �s���x  �s���h  �����h  �����x  �s���x      D   ,  �����x  �����h  �3���h  �3���x  �����x      D   ,  ����x  ����h  �w���h  �w���x  ����x      D   ,  �g���x  �g���h  �����h  �����x  �g���x      D   ,  �����x  �����h  ����h  ����x  �����x      D   ,  ����x  ����h  �k���h  �k���x  ����x      D   ,  �G���x  �G���h  �����h  �����x  �G���x      D   ,  �����x  �����h  ����h  ����x  �����x      D   ,  �����x  �����h  �K���h  �K���x  �����x      D   ,  �;���x  �;���h  �����h  �����x  �;���x      D   ,  ����x  ����h  �����h  �����x  ����x      D   ,  �����x  �����h  �?���h  �?���x  �����x      D   ,  ����x  ����h  �����h  �����x  ����x      D   ,  �s���x  �s���h  �����h  �����x  �s���x      D   ,  �����x  �����h  ����h  ����x  �����x      D   ,  ����x  ����h  �w���h  �w���x  ����x      D   ,  �S���x  �S���h  �����h  �����x  �S���x      D   ,  �����x  �����h  ����h  ����x  �����x      D   ,  �����x  �����h  �W���h  �W���x  �����x      D   ,  �G���x  �G���h  �����h  �����x  �G���x      D   ,  �����x  �����h  �����h  �����x  �����x      D   ,  �����x  �����h  �K���h  �K���x  �����x      D   ,  �'���x  �'���h  �����h  �����x  �'���x      D   ,  ����x  ����h  �����h  �����x  ����x      D   ,  �����x  �����h  �+���h  �+���x  �����x      D   ,  ����x  ����h  �����h  �����x  ����x      D   ,  �_���x  �_���h  �����h  �����x  �_���x      D   ,  �����x  �����h  ����h  ����x  �����x      D   ,  �����x  �����h  �c���h  �c���x  �����x      D   ,  �S���x  �S���h  ƻ���h  ƻ���x  �S���x      D   ,  Ǘ���x  Ǘ���h  �����h  �����x  Ǘ���x      D   ,  �����x  �����h  �W���h  �W���x  �����x      D   ,  �3���x  �3���h  ͛���h  ͛���x  �3���x      D   ,  ΋���x  ΋���h  �����h  �����x  ΋���x      D   ,  �����x  �����h  �7���h  �7���x  �����x      D   ,  \���}  \���  ���  ���}  \���}      D   ,  �w��g�  �w��r�  ����r�  ����g�  �w��g�      D   ,  �A��c�  �A��f�  ����f�  ����c�  �A��c�      D   ,  �w��X  �w��b�  ����b�  ����X  �w��X      D   ,  ΋����  ΋���r  �����r  ������  ΋����      D   ,  ������  �����r  �7���r  �7����  ������      D   ,  �����  ������  ������  �����  �����      D   ,  ����  �����  � ����  � ���  ����      D   ,  �h���  �h����  �N����  �N���  �h���      D   ,  �����  ������  ������  �����  �����      D   ,  ����  �����  ������  �����  ����      D   ,  �R���  �R����  �8����  �8���  �R���      D   ,  �����  ������  ������  �����  �����      D   ,  �����  ������  ������  �����  �����      D   ,  �<���  �<����  �"����  �"���  �<���      D   ,  Ŋ���  Ŋ����  �p����  �p���  Ŋ���      D   ,  �����  ������  Ⱦ����  Ⱦ���  �����      D   ,  �&���  �&����  �����  ����  �&���      D   ,  �t���  �t����  �Z����  �Z���  �t���      D   ,  �����  ������  Ϩ����  Ϩ���  �����      D   ,  ����  �����  ������  �����  ����      D   ,  ����r  �����  � ����  � ���r  ����r      D   ,  �h���r  �h����  �N����  �N���r  �h���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  ����r  �����  ������  �����r  ����r      D   ,  �R���r  �R����  �8����  �8���r  �R���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �<���r  �<����  �"����  �"���r  �<���r      D   ,  Ŋ���r  Ŋ����  �p����  �p���r  Ŋ���r      D   ,  �����r  ������  Ⱦ����  Ⱦ���r  �����r      D   ,  �&���r  �&����  �����  ����r  �&���r      D   ,  �t���r  �t����  �Z����  �Z���r  �t���r      D   ,  �����r  ������  Ϩ����  Ϩ���r  �����r      D   ,  ����r  �����  ������  �����r  ����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  ������  ������  �)����  �)����  ������      D   ,  ������  ������  �w����  �w����  ������      D   ,  �?����  �?����  ������  ������  �?����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �a����  �a����  ������      D   ,  �)����  �)����  ������  ������  �)����      D   ,  �w����  �w����  ������  ������  �w����      D   ,  ������  ������  �K����  �K����  ������      D   ,  �����  �����  ř����  ř����  �����      D   ,  �a����  �a����  ������  ������  �a����      D   ,  ȯ����  ȯ����  �5����  �5����  ȯ����      D   ,  ������  ������  ̃����  ̃����  ������      D   ,  �K����  �K����  ������  ������  �K����      D   ,  ϙ����  ϙ����  �����  �����  ϙ����      D   ,  �����r  ������  ������  �����r  �����r      D   ,  ����r  �����  � ����  � ���r  ����r      D   ,  �h���r  �h����  �N����  �N���r  �h���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  ����r  �����  ������  �����r  ����r      D   ,  �R���r  �R����  �8����  �8���r  �R���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �<���r  �<����  �"����  �"���r  �<���r      D   ,  Ŋ���r  Ŋ����  �p����  �p���r  Ŋ���r      D   ,  �����r  ������  Ⱦ����  Ⱦ���r  �����r      D   ,  �&���r  �&����  �����  ����r  �&���r      D   ,  �t���r  �t����  �Z����  �Z���r  �t���r      D   ,  �����r  ������  Ϩ����  Ϩ���r  �����r      D   ,  ����r  �����  ������  �����r  ����r      D   ,  ������  �����r  �����r  ������  ������      D   ,  ������  �����r  �K���r  �K����  ������      D   ,  �'����  �'���r  �����r  ������  �'����      D   ,  �����  ����r  �����r  ������  �����      D   ,  ������  �����r  �+���r  �+����  ������      D   ,  �����  ����r  �����r  ������  �����      D   ,  �_����  �_���r  �����r  ������  �_����      D   ,  ������  �����r  ����r  �����  ������      D   ,  ������  �����r  �c���r  �c����  ������      D   ,  �S����  �S���r  ƻ���r  ƻ����  �S����      D   ,  Ǘ����  Ǘ���r  �����r  ������  Ǘ����      D   ,  ������  �����r  �W���r  �W����  ������      D   ,  �3����  �3���r  ͛���r  ͛����  �3����      D   ,  ȯ����  ȯ����  �5����  �5����  ȯ����      D   ,  ������  ������  ̃����  ̃����  ������      D   ,  �K����  �K����  ������  ������  �K����      D   ,  ϙ����  ϙ����  �����  �����  ϙ����      D   ,  �����h  ������  ������  �����h  �����h      D   ,  ����h  �����  � ����  � ���h  ����h      D   ,  �h���h  �h����  �N����  �N���h  �h���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  ����h  �����  ������  �����h  ����h      D   ,  �R���h  �R����  �8����  �8���h  �R���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �<���h  �<����  �"����  �"���h  �<���h      D   ,  Ŋ���h  Ŋ����  �p����  �p���h  Ŋ���h      D   ,  �����h  ������  Ⱦ����  Ⱦ���h  �����h      D   ,  �&���h  �&����  �����  ����h  �&���h      D   ,  �t���h  �t����  �Z����  �Z���h  �t���h      D   ,  �����h  ������  Ϩ����  Ϩ���h  �����h      D   ,  ����h  �����  ������  �����h  ����h      D   ,  �����  ����   � ���   � ����  �����      D   ,  �h����  �h���   �N���   �N����  �h����      D   ,  ������  �����   �����   ������  ������      D   ,  �����  ����   �����   ������  �����      D   ,  �R����  �R���   �8���   �8����  �R����      D   ,  ������  �����   �����   ������  ������      D   ,  ������  �����   �����   ������  ������      D   ,  �<����  �<���   �"���   �"����  �<����      D   ,  Ŋ����  Ŋ���   �p���   �p����  Ŋ����      D   ,  ������  �����   Ⱦ���   Ⱦ����  ������      D   ,  �&����  �&���   ����   �����  �&����      D   ,  �t����  �t���   �Z���   �Z����  �t����      D   ,  ������  �����   Ϩ���   Ϩ����  ������      D   ,  �����  ����   �����   ������  �����      D   ,  ������  ������  ������  ������  ������      D   ,  ������  ������  �K����  �K����  ������      D   ,  �'����  �'����  ������  ������  �'����      D   ,  �����  �����  ������  ������  �����      D   ,  ������  ������  �+����  �+����  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �_����  �_����  ������  ������  �_����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �c����  �c����  ������      D   ,  �S����  �S����  ƻ����  ƻ����  �S����      D   ,  Ǘ����  Ǘ����  ������  ������  Ǘ����      D   ,  ������  ������  �W����  �W����  ������      D   ,  �3����  �3����  ͛����  ͛����  �3����      D   ,  ΋����  ΋����  ������  ������  ΋����      D   ,  ������  ������  �7����  �7����  ������      D   ,  �����h  ������  ������  �����h  �����h      D   ,  ����h  �����  � ����  � ���h  ����h      D   ,  �h���h  �h����  �N����  �N���h  �h���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  ����h  �����  ������  �����h  ����h      D   ,  �R���h  �R����  �8����  �8���h  �R���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �<���h  �<����  �"����  �"���h  �<���h      D   ,  Ŋ���h  Ŋ����  �p����  �p���h  Ŋ���h      D   ,  �����h  ������  Ⱦ����  Ⱦ���h  �����h      D   ,  �&���h  �&����  �����  ����h  �&���h      D   ,  �t���h  �t����  �Z����  �Z���h  �t���h      D   ,  �����h  ������  Ϩ����  Ϩ���h  �����h      D   ,  ����h  �����  ������  �����h  ����h      D   ,  ������  �����   �����   ������  ������      D   ,  ������  ������  �)����  �)����  ������      D   ,  ������  ������  �w����  �w����  ������      D   ,  �?����  �?����  ������  ������  �?����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �a����  �a����  ������      D   ,  �)����  �)����  ������  ������  �)����      D   ,  �w����  �w����  ������  ������  �w����      D   ,  ������  ������  �K����  �K����  ������      D   ,  �����  �����  ř����  ř����  �����      D   ,  �a����  �a����  ������  ������  �a����      D   ,  |�����  |�����  ~'����  ~'����  |�����      D   ,  |�����  |�����  ~'����  ~'����  |�����      D   ,  ������  ������  ������  ������  ������      D   ,  }�����  }����r  ?���r  ?����  }�����      D   ,  �/����  �/���r  �����r  ������  �/����      D   ,  �s����  �s���r  �����r  ������  �s����      D   ,  ������  �����r  �3���r  �3����  ������      D   ,  �����  ����r  �w���r  �w����  �����      D   ,  �g����  �g���r  �����r  ������  �g����      D   ,  ������  �����r  ����r  �����  ������      D   ,  �����  ����r  �k���r  �k����  �����      D   ,  �G����  �G���r  �����r  ������  �G����      D   ,  ������  �����r  ����r  �����  ������      D   ,  ������  �����r  �K���r  �K����  ������      D   ,  �;����  �;���r  �����r  ������  �;����      D   ,  �����  ����r  �����r  ������  �����      D   ,  ������  �����r  �?���r  �?����  ������      D   ,  �����  ����r  �����r  ������  �����      D   ,  �s����  �s���r  �����r  ������  �s����      D   ,  ������  �����r  ����r  �����  ������      D   ,  �����  ����r  �w���r  �w����  �����      D   ,  �S����  �S���r  �����r  ������  �S����      D   ,  ������  �����r  ����r  �����  ������      D   ,  ������  �����r  �W���r  �W����  ������      D   ,  �G����  �G���r  �����r  ������  �G����      D   ,  �F���r  �F����  �,����  �,���r  �F���r      D   ,  �����r  ������  �z����  �z���r  �����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �0���r  �0����  �����  ����r  �0���r      D   ,  �~���r  �~����  �d����  �d���r  �~���r      D   ,  �F���r  �F����  �,����  �,���r  �F���r      D   ,  �����r  ������  �z����  �z���r  �����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �0���r  �0����  �����  ����r  �0���r      D   ,  �~���r  �~����  �d����  �d���r  �~���r      D   ,  �I����  �I����  ������  ������  �I����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �k����  �k����  ������      D   ,  �3����  �3����  ������  ������  �3����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �U����  �U����  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �k����  �k����  ������  ������  �k����      D   ,  ������  ������  �?����  �?����  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �r���r  �r����  �X����  �X���r  �r���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  ����r  �����  ������  �����r  ����r      D   ,  �\���r  �\����  �B����  �B���r  �\���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �r���r  �r����  �X����  �X���r  �r���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  ����r  �����  ������  �����r  ����r      D   ,  �\���r  �\����  �B����  �B���r  �\���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �:���r  �:����  � ����  � ���r  �:���r      D   ,  �����r  ������  �n����  �n���r  �����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �$���r  �$����  �
����  �
���r  �$���r      D   ,  �=����  �=����  ������  ������  �=����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �_����  �_����  ������      D   ,  �'����  �'����  ������  ������  �'����      D   ,  �u����  �u����  ������  ������  �u����      D   ,  ������  ������  �I����  �I����  ������      D   ,  ~���r  ~����  ~�����  ~����r  ~���r      D   ,  �f���r  �f����  �L����  �L���r  �f���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  ����r  �����  ������  �����r  ����r      D   ,  �P���r  �P����  �6����  �6���r  �P���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �:���r  �:����  � ����  � ���r  �:���r      D   ,  �����r  ������  �n����  �n���r  �����r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  �$���r  �$����  �
����  �
���r  �$���r      D   ,  �����  �����  ������  ������  �����      D   ,  �_����  �_����  ������  ������  �_����      D   ,  ������  ������  �3����  �3����  ������      D   ,  ~�����  ~�����  �u����  �u����  ~�����      D   ,  �����r  ������  ������  �����r  �����r      D   ,  ����r  �����  ������  �����r  ����r      D   ,  �P���r  �P����  �6����  �6���r  �P���r      D   ,  �����r  ������  ������  �����r  �����r      D   ,  ~���r  ~����  ~�����  ~����r  ~���r      D   ,  �f���r  �f����  �L����  �L���r  �f���r      D   ,  �����  ������  ������  �����  �����      D   ,  �����  ������  ������  �����  �����      D   ,  �:���  �:����  � ����  � ���  �:���      D   ,  �����  ������  �n����  �n���  �����      D   ,  �����  ������  ������  �����  �����      D   ,  �$���  �$����  �
����  �
���  �$���      D   ,  ~���  ~����  ~�����  ~����  ~���      D   ,  �����  ������  ������  �����  �����      D   ,  ����  �����  ������  �����  ����      D   ,  �P���  �P����  �6����  �6���  �P���      D   ,  �f���  �f����  �L����  �L���  �f���      D   ,  �����  ������  ������  �����  �����      D   ,  ����  �����  ������  �����  ����      D   ,  �\���  �\����  �B����  �B���  �\���      D   ,  �����  ������  ������  �����  �����      D   ,  �����  ������  ������  �����  �����      D   ,  �F���  �F����  �,����  �,���  �F���      D   ,  �����  ������  �z����  �z���  �����      D   ,  �����  ������  ������  �����  �����      D   ,  �0���  �0����  �����  ����  �0���      D   ,  �~���  �~����  �d����  �d���  �~���      D   ,  �r���  �r����  �X����  �X���  �r���      D   ,  y|���r  y|����  zb����  zb���r  y|���r      D   ,  {����r  {�����  |�����  |����r  {����r      D   ,  x����  x����  y�����  y�����  x����      D   ,  `"���r  `"����  a����  a���r  `"���r      D   ,  bp���r  bp����  cV����  cV���r  bp���r      D   ,  d����r  d�����  e�����  e����r  d����r      D   ,  g���r  g����  g�����  g����r  g���r      D   ,  iZ���r  iZ����  j@����  j@���r  iZ���r      D   ,  k����r  k�����  l�����  l����r  k����r      D   ,  m����r  m�����  n�����  n����r  m����r      D   ,  pD���r  pD����  q*����  q*���r  pD���r      D   ,  r����r  r�����  sx����  sx���r  r����r      D   ,  t����r  t�����  u�����  u����r  t����r      D   ,  ]�����  ]����r  ^����r  ^�����  ]�����      D   ,  _�����  _����r  aS���r  aS����  _�����      D   ,  b/����  b/���r  c����r  c�����  b/����      D   ,  d�����  d����r  e����r  e�����  d�����      D   ,  f�����  f����r  h3���r  h3����  f�����      D   ,  i#����  i#���r  j����r  j�����  i#����      D   ,  kg����  kg���r  l����r  l�����  kg����      D   ,  m�����  m����r  o'���r  o'����  m�����      D   ,  p����  p���r  qk���r  qk����  p����      D   ,  r[����  r[���r  s����r  s�����  r[����      D   ,  t�����  t����r  v���r  v����  t�����      D   ,  v�����  v����r  x_���r  x_����  v�����      D   ,  y;����  y;���r  z����r  z�����  y;����      D   ,  {�����  {����r  |����r  |�����  {�����      D   ,  zS����  zS����  {�����  {�����  zS����      D   ,  k����  k�����  l�����  l����  k����      D   ,  m����  m�����  n�����  n����  m����      D   ,  pD���  pD����  q*����  q*���  pD���      D   ,  r����  r�����  sx����  sx���  r����      D   ,  t����  t�����  u�����  u����  t����      D   ,  w.���  w.����  x����  x���  w.���      D   ,  y|���  y|����  zb����  zb���  y|���      D   ,  {����  {�����  |�����  |����  {����      D   ,  g���  g����  g�����  g����  g���      D   ,  iZ���  iZ����  j@����  j@���  iZ���      D   ,  u�����  u�����  w=����  w=����  u�����      D   ,  ]����r  ]�����  ^�����  ^����r  ]����r      D   ,  `"���r  `"����  a����  a���r  `"���r      D   ,  bp���r  bp����  cV����  cV���r  bp���r      D   ,  d����r  d�����  e�����  e����r  d����r      D   ,  g���r  g����  g�����  g����r  g���r      D   ,  iZ���r  iZ����  j@����  j@���r  iZ���r      D   ,  k����r  k�����  l�����  l����r  k����r      D   ,  m����r  m�����  n�����  n����r  m����r      D   ,  pD���r  pD����  q*����  q*���r  pD���r      D   ,  r����r  r�����  sx����  sx���r  r����r      D   ,  w.���r  w.����  x����  x���r  w.���r      D   ,  y|���r  y|����  zb����  zb���r  y|���r      D   ,  {����r  {�����  |�����  |����r  {����r      D   ,  t����r  t�����  u�����  u����r  t����r      D   ,  w.���r  w.����  x����  x���r  w.���r      D   ,  ^�����  ^�����  `1����  `1����  ^�����      D   ,  `�����  `�����  b����  b����  `�����      D   ,  cG����  cG����  d�����  d�����  cG����      D   ,  e�����  e�����  g����  g����  e�����      D   ,  g�����  g�����  ii����  ii����  g�����      D   ,  j1����  j1����  k�����  k�����  j1����      D   ,  l����  l����  n����  n����  l����      D   ,  n�����  n�����  pS����  pS����  n�����      D   ,  q����  q����  r�����  r�����  q����      D   ,  si����  si����  t�����  t�����  si����      D   ,  ]����  ]�����  ^�����  ^����  ]����      D   ,  `"���  `"����  a����  a���  `"���      D   ,  bp���  bp����  cV����  cV���  bp���      D   ,  d����  d�����  e�����  e����  d����      D   ,  ]����r  ]�����  ^�����  ^����r  ]����r      D   ,  {����h  {�����  |�����  |����h  {����h      D   ,  d�����  d�����  e�����  e�����  d�����      D   ,  f�����  f�����  h3����  h3����  f�����      D   ,  i#����  i#����  j�����  j�����  i#����      D   ,  kg����  kg����  l�����  l�����  kg����      D   ,  m�����  m�����  o'����  o'����  m�����      D   ,  p����  p����  qk����  qk����  p����      D   ,  r[����  r[����  s�����  s�����  r[����      D   ,  t�����  t�����  v����  v����  t�����      D   ,  v�����  v�����  x_����  x_����  v�����      D   ,  y;����  y;����  z�����  z�����  y;����      D   ,  {�����  {�����  |�����  |�����  {�����      D   ,  iZ����  iZ���   j@���   j@����  iZ����      D   ,  k�����  k����   l����   l�����  k�����      D   ,  m�����  m����   n����   n�����  m�����      D   ,  pD����  pD���   q*���   q*����  pD����      D   ,  ^�����  ^�����  `1����  `1����  ^�����      D   ,  `�����  `�����  b����  b����  `�����      D   ,  cG����  cG����  d�����  d�����  cG����      D   ,  e�����  e�����  g����  g����  e�����      D   ,  g�����  g�����  ii����  ii����  g�����      D   ,  j1����  j1����  k�����  k�����  j1����      D   ,  l����  l����  n����  n����  l����      D   ,  n�����  n�����  pS����  pS����  n�����      D   ,  q����  q����  r�����  r�����  q����      D   ,  si����  si����  t�����  t�����  si����      D   ,  u�����  u�����  w=����  w=����  u�����      D   ,  x����  x����  y�����  y�����  x����      D   ,  zS����  zS����  {�����  {�����  zS����      D   ,  r�����  r����   sx���   sx����  r�����      D   ,  t�����  t����   u����   u�����  t�����      D   ,  w.����  w.���   x���   x����  w.����      D   ,  y|����  y|���   zb���   zb����  y|����      D   ,  {�����  {����   |����   |�����  {�����      D   ,  bp����  bp���   cV���   cV����  bp����      D   ,  d�����  d����   e����   e�����  d�����      D   ,  g����  g���   g����   g�����  g����      D   ,  ]�����  ]�����  ^�����  ^�����  ]�����      D   ,  _�����  _�����  aS����  aS����  _�����      D   ,  b/����  b/����  c�����  c�����  b/����      D   ,  bp���h  bp����  cV����  cV���h  bp���h      D   ,  d����h  d�����  e�����  e����h  d����h      D   ,  g���h  g����  g�����  g����h  g���h      D   ,  iZ���h  iZ����  j@����  j@���h  iZ���h      D   ,  k����h  k�����  l�����  l����h  k����h      D   ,  ]����h  ]�����  ^�����  ^����h  ]����h      D   ,  `"���h  `"����  a����  a���h  `"���h      D   ,  bp���h  bp����  cV����  cV���h  bp���h      D   ,  d����h  d�����  e�����  e����h  d����h      D   ,  g���h  g����  g�����  g����h  g���h      D   ,  iZ���h  iZ����  j@����  j@���h  iZ���h      D   ,  k����h  k�����  l�����  l����h  k����h      D   ,  m����h  m�����  n�����  n����h  m����h      D   ,  pD���h  pD����  q*����  q*���h  pD���h      D   ,  r����h  r�����  sx����  sx���h  r����h      D   ,  t����h  t�����  u�����  u����h  t����h      D   ,  w.���h  w.����  x����  x���h  w.���h      D   ,  y|���h  y|����  zb����  zb���h  y|���h      D   ,  {����h  {�����  |�����  |����h  {����h      D   ,  m����h  m�����  n�����  n����h  m����h      D   ,  pD���h  pD����  q*����  q*���h  pD���h      D   ,  r����h  r�����  sx����  sx���h  r����h      D   ,  t����h  t�����  u�����  u����h  t����h      D   ,  w.���h  w.����  x����  x���h  w.���h      D   ,  y|���h  y|����  zb����  zb���h  y|���h      D   ,  ������  ������  �3����  �3����  ������      D   ,  �����  �����  �w����  �w����  �����      D   ,  �g����  �g����  ������  ������  �g����      D   ,  ������  ������  �����  �����  ������      D   ,  �����  �����  �k����  �k����  �����      D   ,  �G����  �G����  ������  ������  �G����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �K����  �K����  ������      D   ,  �;����  �;����  ������  ������  �;����      D   ,  �����  �����  ������  ������  �����      D   ,  ������  ������  �?����  �?����  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �s����  �s����  ������  ������  �s����      D   ,  ������  ������  �����  �����  ������      D   ,  �����  �����  �w����  �w����  �����      D   ,  �S����  �S����  ������  ������  �S����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �W����  �W����  ������      D   ,  �G����  �G����  ������  ������  �G����      D   ,  ������  ������  ������  ������  ������      D   ,  }�����  }�����  ?����  ?����  }�����      D   ,  �/����  �/����  ������  ������  �/����      D   ,  �s����  �s����  ������  ������  �s����      D   ,  ������  �����   �����   ������  ������      D   ,  ������  �����   �����   ������  ������      D   ,  �F����  �F���   �,���   �,����  �F����      D   ,  ������  �����   �z���   �z����  ������      D   ,  �r����  �r���   �X���   �X����  �r����      D   ,  ������  �����   �����   ������  ������      D   ,  �0����  �0���   ����   �����  �0����      D   ,  �~����  �~���   �d���   �d����  �~����      D   ,  ������  �����   �����   ������  ������      D   ,  �����  ����   �����   ������  �����      D   ,  �\����  �\���   �B���   �B����  �\����      D   ,  �$����  �$���   �
���   �
����  �$����      D   ,  ~����  ~���   ~����   ~�����  ~����      D   ,  �f����  �f���   �L���   �L����  �f����      D   ,  ������  �����   �����   ������  ������      D   ,  �����  ����   �����   ������  �����      D   ,  �P����  �P���   �6���   �6����  �P����      D   ,  ������  �����   �����   ������  ������      D   ,  ������  �����   �����   ������  ������      D   ,  �:����  �:���   � ���   � ����  �:����      D   ,  ������  �����   �n���   �n����  ������      D   ,  ������  �����   �����   ������  ������      D   ,  �$���h  �$����  �
����  �
���h  �$���h      D   ,  ~���h  ~����  ~�����  ~����h  ~���h      D   ,  �f���h  �f����  �L����  �L���h  �f���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  ����h  �����  ������  �����h  ����h      D   ,  �P���h  �P����  �6����  �6���h  �P���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  ~�����  ~�����  �u����  �u����  ~�����      D   ,  �=����  �=����  ������  ������  �=����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �_����  �_����  ������      D   ,  �'����  �'����  ������  ������  �'����      D   ,  �u����  �u����  ������  ������  �u����      D   ,  ������  ������  �I����  �I����  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �_����  �_����  ������  ������  �_����      D   ,  ������  ������  �3����  �3����  ������      D   ,  �:���h  �:����  � ����  � ���h  �:���h      D   ,  �����h  ������  �n����  �n���h  �����h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �$���h  �$����  �
����  �
���h  �$���h      D   ,  ~���h  ~����  ~�����  ~����h  ~���h      D   ,  �f���h  �f����  �L����  �L���h  �f���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  ����h  �����  ������  �����h  ����h      D   ,  �P���h  �P����  �6����  �6���h  �P���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �:���h  �:����  � ����  � ���h  �:���h      D   ,  �����h  ������  �n����  �n���h  �����h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �F���h  �F����  �,����  �,���h  �F���h      D   ,  �����h  ������  �z����  �z���h  �����h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �0���h  �0����  �����  ����h  �0���h      D   ,  �~���h  �~����  �d����  �d���h  �~���h      D   ,  �\���h  �\����  �B����  �B���h  �\���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �F���h  �F����  �,����  �,���h  �F���h      D   ,  �I����  �I����  ������  ������  �I����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �k����  �k����  ������      D   ,  �3����  �3����  ������  ������  �3����      D   ,  ������  ������  �����  �����  ������      D   ,  ������  ������  �U����  �U����  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �k����  �k����  ������  ������  �k����      D   ,  ������  ������  �?����  �?����  ������      D   ,  �����  �����  ������  ������  �����      D   ,  �����h  ������  �z����  �z���h  �����h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �0���h  �0����  �����  ����h  �0���h      D   ,  �~���h  �~����  �d����  �d���h  �~���h      D   ,  ����h  �����  ������  �����h  ����h      D   ,  �r���h  �r����  �X����  �X���h  �r���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �r���h  �r����  �X����  �X���h  �r���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  ����h  �����  ������  �����h  ����h      D   ,  �\���h  �\����  �B����  �B���h  �\���h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  �����h  ������  ������  �����h  �����h      D   ,  re��g�  re��r�  s���r�  s���g�  re��g�      D   ,  t���g�  t���r�  v��r�  v��g�  t���g�      D   ,  w��g�  w��r�  xi��r�  xi��g�  w��g�      D   ,  yO��g�  yO��r�  z���r�  z���g�  yO��g�      D   ,  {���g�  {���r�  }��r�  }��g�  {���g�      D   ,  }���g�  }���r�  S��r�  S��g�  }���g�      D   ,  �9��g�  �9��r�  ����r�  ����g�  �9��g�      D   ,  ����g�  ����r�  ����r�  ����g�  ����g�      D   ,  ����g�  ����r�  �=��r�  �=��g�  ����g�      D   ,  �#��g�  �#��r�  ����r�  ����g�  �#��g�      D   ,  �q��g�  �q��r�  ����r�  ����g�  �q��g�      D   ,  ����g�  ����r�  �'��r�  �'��g�  ����g�      D   ,  ���g�  ���r�  �u��r�  �u��g�  ���g�      D   ,  �[��g�  �[��r�  ����r�  ����g�  �[��g�      D   ,  ����g�  ����r�  ���r�  ���g�  ����g�      D   ,  ����g�  ����r�  �_��r�  �_��g�  ����g�      D   ,  �k��g�  �k��r�  ����r�  ����g�  �k��g�      D   ,  ����g�  ����r�  �!��r�  �!��g�  ����g�      D   ,  ���g�  ���r�  �o��r�  �o��g�  ���g�      D   ,  �U��g�  �U��r�  ����r�  ����g�  �U��g�      D   ,  ����g�  ����r�  ���r�  ���g�  ����g�      D   ,  ����g�  ����r�  �Y��r�  �Y��g�  ����g�      D   ,  �?��g�  �?��r�  ����r�  ����g�  �?��g�      D   ,  ����g�  ����r�  ����r�  ����g�  ����g�      D   ,  ����g�  ����r�  �C��r�  �C��g�  ����g�      D   ,  �)��g�  �)��r�  ����r�  ����g�  �)��g�      D   ,  |���c�  |���f�  ~;��f�  ~;��c�  |���c�      D   ,  ���  �����  �����  ���  ���      D   ,  ����  ������  ������  ����  ����      D   ,  �M��  �M����  �Q����  �Q��  �M��      D   ,  ����  ������  ������  ����  ����      D   ,  ����  ������  ������  ����  ����      D   ,  �!��  �!����  �%����  �%��  �!��      D   ,  ~	��{�  ~	��}  ��}  ��{�  ~	��{�      D   ,  ����{�  ����}  ����}  ����{�  ����{�      D   ,  �A��{�  �A��}  �E��}  �E��{�  �A��{�      D   ,  ����{�  ����}  ����}  ����{�  ����{�      D   ,  �y��{�  �y��}  �}��}  �}��{�  �y��{�      D   ,  ���{�  ���}  ���}  ���{�  ���{�      D   ,  ����{�  ����}  ����}  ����{�  ����{�      D   ,  �M��{�  �M��}  �Q��}  �Q��{�  �M��{�      D   ,  ����{�  ����}  ����}  ����{�  ����{�      D   ,  ����{�  ����}  ����}  ����{�  ����{�      D   ,  �!��{�  �!��}  �%��}  �%��{�  �!��{�      D   ,  ~,��r�  ~,��sQ  ��sQ  ��r�  ~,��r�      D   ,  �z��r�  �z��sQ  �`��sQ  �`��r�  �z��r�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  ���r�  ���sQ  ����sQ  ����r�  ���r�      D   ,  �d��r�  �d��sQ  �J��sQ  �J��r�  �d��r�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  � ��r�  � ��sQ  ����sQ  ����r�  � ��r�      D   ,  �N��r�  �N��sQ  �4��sQ  �4��r�  �N��r�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  �8��r�  �8��sQ  ���sQ  ���r�  �8��r�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  �H��r�  �H��sQ  �.��sQ  �.��r�  �H��r�      D   ,  ����r�  ����sQ  �|��sQ  �|��r�  ����r�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  �2��r�  �2��sQ  ���sQ  ���r�  �2��r�      D   ,  ����r�  ����sQ  �f��sQ  �f��r�  ����r�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  ���r�  ���sQ  ���sQ  ���r�  ���r�      D   ,  �j��r�  �j��sQ  �P��sQ  �P��r�  �j��r�      D   ,  ~���  ~���x  ~����x  ~����  ~���      D   ,  �f���  �f���x  �L���x  �L���  �f���      D   ,  �����  �����x  �����x  �����  �����      D   ,  ����  ����x  �����x  �����  ����      D   ,  �P���  �P���x  �6���x  �6���  �P���      D   ,  �����  �����x  �����x  �����  �����      D   ,  �����  �����x  �����x  �����  �����      D   ,  �:���  �:���x  � ���x  � ���  �:���      D   ,  �����  �����x  �n���x  �n���  �����      D   ,  �����  �����x  �����x  �����  �����      D   ,  �$���  �$���x  �
���x  �
���  �$���      D   ,  �r���  �r���x  �X���x  �X���  �r���      D   ,  �����  �����x  �����x  �����  �����      D   ,  ����  ����x  �����x  �����  ����      D   ,  �\���  �\���x  �B���x  �B���  �\���      D   ,  �����  �����x  �����x  �����  �����      D   ,  �����  �����x  �����x  �����  �����      D   ,  �F���  �F���x  �,���x  �,���  �F���      D   ,  �����  �����x  �z���x  �z���  �����      D   ,  �����  �����x  �����x  �����  �����      D   ,  �0���  �0���x  ����x  ����  �0���      D   ,  �~���  �~���x  �d���x  �d���  �~���      D   ,  ~	��  ~	����  ����  ��  ~	��      D   ,  ����  ������  ������  ����  ����      D   ,  �A��  �A����  �E����  �E��  �A��      D   ,  ����  ������  ������  ����  ����      D   ,  �y��  �y����  �}����  �}��  �y��      D   ,  t����  t����x  u����x  u����  t����      D   ,  w.���  w.���x  x���x  x���  w.���      D   ,  y|���  y|���x  zb���x  zb���  y|���      D   ,  {����  {����x  |����x  |����  {����      D   ,  iZ���  iZ���x  j@���x  j@���  iZ���      D   ,  J���p1  J���{!  K���{!  K���p1  J���p1      D   ,  N\��p1  N\��{!  O���{!  O���p1  N\��p1      D   ,  wB��r�  wB��sQ  x(��sQ  x(��r�  wB��r�      D   ,  y���r�  y���sQ  zv��sQ  zv��r�  y���r�      D   ,  {���r�  {���sQ  |���sQ  |���r�  {���r�      D   ,  k����  k����x  l����x  l����  k����      D   ,  m����  m����x  n����x  n����  m����      D   ,  pD���  pD���x  q*���x  q*���  pD���      D   ,  ]���  ]�����  ^�����  ^���  ]���      D   ,  ba��  ba����  ce����  ce��  ba��      D   ,  ]����  ]����x  ^����x  ^����  ]����      D   ,  ]���{�  ]���}  ^���}  ^���{�  ]���{�      D   ,  ba��{�  ba��}  ce��}  ce��{�  ba��{�      D   ,  f���{�  f���}  h��}  h��{�  f���{�      D   ,  k���{�  k���}  l���}  l���{�  k���{�      D   ,  p5��{�  p5��}  q9��}  q9��{�  p5��{�      D   ,  t���{�  t���}  u���}  u���{�  t���{�      D   ,  ym��{�  ym��}  zq��}  zq��{�  ym��{�      D   ,  f���  f�����  h����  h��  f���      D   ,  k���  k�����  l�����  l���  k���      D   ,  p5��  p5����  q9����  q9��  p5��      D   ,  t���  t�����  u�����  u���  t���      D   ,  ym��  ym����  zq����  zq��  ym��      D   ,  `"���  `"���x  a���x  a���  `"���      D   ,  r����  r����x  sx���x  sx���  r����      D   ,  bp���  bp���x  cV���x  cV���  bp���      D   ,  d����  d����x  e����x  e����  d����      D   ,  g���  g���x  g����x  g����  g���      D   ,  u���c�  u���f�  wQ��f�  wQ��c�  u���c�      D   ,  x��c�  x��f�  y���f�  y���c�  x��c�      D   ,  zg��c�  zg��f�  {���f�  {���c�  zg��c�      D   ,  wB��g�  wB��g�  x(��g�  x(��g�  wB��g�      D   ,  y���g�  y���g�  zv��g�  zv��g�  y���g�      D   ,  r���b�  r���cW  s���cW  s���b�  r���b�      D   ,  t���b�  t���cW  u���cW  u���b�  t���b�      D   ,  wB��b�  wB��cW  x(��cW  x(��b�  wB��b�      D   ,  y���b�  y���cW  zv��cW  zv��b�  y���b�      D   ,  {���b�  {���cW  |���cW  |���b�  {���b�      D   ,  re��X  re��b�  s���b�  s���X  re��X      D   ,  t���X  t���b�  v��b�  v��X  t���X      D   ,  w��X  w��b�  xi��b�  xi��X  w��X      D   ,  yO��X  yO��b�  z���b�  z���X  yO��X      D   ,  {���X  {���b�  }��b�  }��X  {���X      D   ,  {���g�  {���g�  |���g�  |���g�  {���g�      D   ,  r���W�  r���X  s���X  s���W�  r���W�      D   ,  t���W�  t���X  u���X  u���W�  t���W�      D   ,  wB��W�  wB��X  x(��X  x(��W�  wB��W�      D   ,  y���W�  y���X  zv��X  zv��W�  y���W�      D   ,  {���W�  {���X  |���X  |���W�  {���W�      D   ,  s}��c�  s}��f�  u��f�  u��c�  s}��c�      D   ,  }���X  }���b�  S��b�  S��X  }���X      D   ,  �9��X  �9��b�  ����b�  ����X  �9��X      D   ,  ����X  ����b�  ����b�  ����X  ����X      D   ,  ����X  ����b�  �=��b�  �=��X  ����X      D   ,  �#��X  �#��b�  ����b�  ����X  �#��X      D   ,  �q��X  �q��b�  ����b�  ����X  �q��X      D   ,  ����X  ����b�  �'��b�  �'��X  ����X      D   ,  ���X  ���b�  �u��b�  �u��X  ���X      D   ,  �[��X  �[��b�  ����b�  ����X  �[��X      D   ,  ����X  ����b�  ���b�  ���X  ����X      D   ,  ����X  ����b�  �_��b�  �_��X  ����X      D   ,  �k��X  �k��b�  ����b�  ����X  �k��X      D   ,  ����X  ����b�  �!��b�  �!��X  ����X      D   ,  ���X  ���b�  �o��b�  �o��X  ���X      D   ,  �U��X  �U��b�  ����b�  ����X  �U��X      D   ,  ����X  ����b�  ���b�  ���X  ����X      D   ,  ����X  ����b�  �Y��b�  �Y��X  ����X      D   ,  �?��X  �?��b�  ����b�  ����X  �?��X      D   ,  ����X  ����b�  ����b�  ����X  ����X      D   ,  ����X  ����b�  �C��b�  �C��X  ����X      D   ,  �)��X  �)��b�  ����b�  ����X  �)��X      D   ,  �H��g�  �H��g�  �.��g�  �.��g�  �H��g�      D   ,  ����g�  ����g�  �|��g�  �|��g�  ����g�      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  ����c�  ����f�  �	��f�  �	��c�  ����c�      D   ,  ����c�  ����f�  �W��f�  �W��c�  ����c�      D   ,  ���c�  ���f�  ����f�  ����c�  ���c�      D   ,  �m��c�  �m��f�  ����f�  ����c�  �m��c�      D   ,  ����c�  ����f�  �A��f�  �A��c�  ����c�      D   ,  �	��c�  �	��f�  ����f�  ����c�  �	��c�      D   ,  �W��c�  �W��f�  ����f�  ����c�  �W��c�      D   ,  ����c�  ����f�  �+��f�  �+��c�  ����c�      D   ,  ����c�  ����f�  �y��f�  �y��c�  ����c�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  �H��b�  �H��cW  �.��cW  �.��b�  �H��b�      D   ,  ����b�  ����cW  �|��cW  �|��b�  ����b�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  �2��b�  �2��cW  ���cW  ���b�  �2��b�      D   ,  ����b�  ����cW  �f��cW  �f��b�  ����b�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  ���b�  ���cW  ���cW  ���b�  ���b�      D   ,  �j��b�  �j��cW  �P��cW  �P��b�  �j��b�      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  �2��g�  �2��g�  ���g�  ���g�  �2��g�      D   ,  ����g�  ����g�  �f��g�  �f��g�  ����g�      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  ���g�  ���g�  ���g�  ���g�  ���g�      D   ,  �j��g�  �j��g�  �P��g�  �P��g�  �j��g�      D   ,  �;��c�  �;��f�  ����f�  ����c�  �;��c�      D   ,  ����c�  ����f�  ���f�  ���c�  ����c�      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  � ��g�  � ��g�  ����g�  ����g�  � ��g�      D   ,  �N��g�  �N��g�  �4��g�  �4��g�  �N��g�      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  �8��g�  �8��g�  ���g�  ���g�  �8��g�      D   ,  ~,��b�  ~,��cW  ��cW  ��b�  ~,��b�      D   ,  �z��b�  �z��cW  �`��cW  �`��b�  �z��b�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  ���b�  ���cW  ����cW  ����b�  ���b�      D   ,  �d��b�  �d��cW  �J��cW  �J��b�  �d��b�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  � ��b�  � ��cW  ����cW  ����b�  � ��b�      D   ,  �N��b�  �N��cW  �4��cW  �4��b�  �N��b�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  �8��b�  �8��cW  ���cW  ���b�  �8��b�      D   ,  ����c�  ����f�  �]��f�  �]��c�  ����c�      D   ,  �%��c�  �%��f�  ����f�  ����c�  �%��c�      D   ,  �s��c�  �s��f�  ����f�  ����c�  �s��c�      D   ,  ����c�  ����f�  �G��f�  �G��c�  ����c�      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  ���g�  ���g�  ����g�  ����g�  ���g�      D   ,  �d��g�  �d��g�  �J��g�  �J��g�  �d��g�      D   ,  ��c�  ��f�  ����f�  ����c�  ��c�      D   ,  �Q��c�  �Q��f�  ����f�  ����c�  �Q��c�      D   ,  ����c�  ����f�  �%��f�  �%��c�  ����c�      D   ,  ����c�  ����f�  �s��f�  �s��c�  ����c�      D   ,  ~,��g�  ~,��g�  ��g�  ��g�  ~,��g�      D   ,  �z��g�  �z��g�  �`��g�  �`��g�  �z��g�      D   ,  �z��W�  �z��X  �`��X  �`��W�  �z��W�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  ���W�  ���X  ����X  ����W�  ���W�      D   ,  �d��W�  �d��X  �J��X  �J��W�  �d��W�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  � ��W�  � ��X  ����X  ����W�  � ��W�      D   ,  �N��W�  �N��X  �4��X  �4��W�  �N��W�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  �8��W�  �8��X  ���X  ���W�  �8��W�      D   ,  ~,��W�  ~,��X  ��X  ��W�  ~,��W�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  �H��W�  �H��X  �.��X  �.��W�  �H��W�      D   ,  ����W�  ����X  �|��X  �|��W�  ����W�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  �2��W�  �2��X  ���X  ���W�  �2��W�      D   ,  ����W�  ����X  �f��X  �f��W�  ����W�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  ���W�  ���X  ���X  ���W�  ���W�      D   ,  �j��W�  �j��X  �P��X  �P��W�  �j��W�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  ����g�  ����r�  �-��r�  �-��g�  ����g�      D   ,  ���g�  ���r�  �{��r�  �{��g�  ���g�      D   ,  �a��g�  �a��r�  ����r�  ����g�  �a��g�      D   ,  ����g�  ����r�  ���r�  ���g�  ����g�      D   ,  ����g�  ����r�  �e��r�  �e��g�  ����g�      D   ,  ̜��U�  ̜��r�  ����r�  ����U�  ̜��U�      D   ,  �o��b�  �o��s  ����s  ����b�  �o��b�      D   ,  �S��b�  �S��s  ����s  ����b�  �S��b�      D   ,  �7��b�  �7��s  ����s  ����b�  �7��b�      D   ,  ���b�  ���s  ����s  ����b�  ���b�      D   ,  ����b�  ����s g��s g��b�  ����b�      D   , ���b� ���s K��s K��b� ���b�      D   , ���b� ���s /��s /��b� ���b�      D   , ���b� ���s 
��s 
��b� ���b�      D   , ���b� ���s ���s ���b� ���b�      D   , s��b� s��s ���s ���b� s��b�      D   , W��b� W��s ���s ���b� W��b�      D   , ;��b� ;��s ���s ���b� ;��b�      D   , ��s ��sQ ���sQ ���s ��s      D   , ���s ���sQ 	���sQ 	���s ���s      D   , ���s ���sQ ���sQ ���s ���s      D   , ���s ���sQ ���sQ ���s ���s      D   , ���s ���sQ ~��sQ ~��s ���s      D   , |��s |��sQ b��sQ b��s |��s      D   ,  ����s  ����sQ  ����sQ  ����s  ����s      D   ,  ����s  ����sQ  �z��sQ  �z��s  ����s      D   ,  �x��s  �x��sQ  �^��sQ  �^��s  �x��s      D   ,  �\��s  �\��sQ  �B��sQ  �B��s  �\��s      D   ,  @��s  @��sQ &��sQ &��s  @��s      D   , $��s $��sQ 
��sQ 
��s $��s      D   ,  �t���  �t���x  �Z���x  �Z���  �t���      D   ,  �����  �����x  Ϩ���x  Ϩ���  �����      D   ,  ����  ����x  �����x  �����  ����      D   ,  �����  �����x  �����x  �����  �����      D   ,  ����  ����x  � ���x  � ���  ����      D   ,  �h���  �h���x  �N���x  �N���  �h���      D   ,  ����  ������  ������  ����  ����      D   ,  �Y��  �Y����  �]����  �]��  �Y��      D   ,  ����  ������  ������  ����  ����      D   ,  ����{�  ����}  ����}  ����{�  ����{�      D   ,  �-��{�  �-��}  �1��}  �1��{�  �-��{�      D   ,  ����{�  ����}  ����}  ����{�  ����{�      D   ,  �e��{�  �e��}  �i��}  �i��{�  �e��{�      D   ,  ���{�  ���}  ���}  ���{�  ���{�      D   ,  ����  ������  ������  ����  ����      D   ,  ����{�  ����}  ����}  ����{�  ����{�      D   ,  �Y��{�  �Y��}  �]��}  �]��{�  �Y��{�      D   ,  ����{�  ����}  ����}  ����{�  ����{�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  ���r�  ���sQ  ����sQ  ����r�  ���r�      D   ,  �T��r�  �T��sQ  �:��sQ  �:��r�  �T��r�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  ����r�  ����sQ  ����sQ  ����r�  ����r�      D   ,  �-��  �-����  �1����  �1��  �-��      D   ,  ����  ������  ������  ����  ����      D   ,  �e��  �e����  �i����  �i��  �e��      D   ,  ���  �����  �����  ���  ���      D   ,  �����  �����x  �����x  �����  �����      D   ,  ����  ����x  �����x  �����  ����      D   ,  �R���  �R���x  �8���x  �8���  �R���      D   ,  �����  �����x  �����x  �����  �����      D   ,  �����  �����x  �����x  �����  �����      D   ,  �<���  �<���x  �"���x  �"���  �<���      D   ,  Ŋ���  Ŋ���x  �p���x  �p���  Ŋ���      D   ,  �����  �����x  Ⱦ���x  Ⱦ���  �����      D   ,  �&���  �&���x  ����x  ����  �&���      D   ,  �>��r�  �>��sQ  �$��sQ  �$��r�  �>��r�      D   ,  ���X  ���b�  �{��b�  �{��X  ���X      D   ,  �a��X  �a��b�  ����b�  ����X  �a��X      D   ,  ����X  ����b�  ���b�  ���X  ����X      D   ,  ����X  ����b�  �e��b�  �e��X  ����X      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  ���g�  ���g�  ����g�  ����g�  ���g�      D   ,  �T��g�  �T��g�  �:��g�  �:��g�  �T��g�      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  ���W�  ���X  ����X  ����W�  ���W�      D   ,  �T��W�  �T��X  �:��X  �:��W�  �T��W�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  ����W�  ����X  ����X  ����W�  ����W�      D   ,  �>��W�  �>��X  �$��X  �$��W�  �>��W�      D   ,  ����g�  ����g�  ����g�  ����g�  ����g�      D   ,  �>��g�  �>��g�  �$��g�  �$��g�  �>��g�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  ����c�  ����f�  ���f�  ���c�  ����c�      D   ,  ����c�  ����f�  �c��f�  �c��c�  ����c�      D   ,  �+��c�  �+��f�  ����f�  ����c�  �+��c�      D   ,  �y��c�  �y��f�  ����f�  ����c�  �y��c�      D   ,  ����c�  ����f�  �M��f�  �M��c�  ����c�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  �>��b�  �>��cW  �$��cW  �$��b�  �>��b�      D   ,  ����b�  ����cW  ����cW  ����b�  ����b�      D   ,  ���b�  ���cW  ����cW  ����b�  ���b�      D   ,  �T��b�  �T��cW  �:��cW  �:��b�  �T��b�      D   ,  ����X  ����b�  �-��b�  �-��X  ����X      D   ,  ����a�  ����b�  �z��b�  �z��a�  ����a�      D   ,  �x��a�  �x��b�  �^��b�  �^��a�  �x��a�      D   ,  �\��a�  �\��b�  �B��b�  �B��a�  �\��a�      D   ,  @��a�  @��b� &��b� &��a�  @��a�      D   , $��a� $��b� 
��b� 
��a� $��a�      D   , ��a� ��b� ���b� ���a� ��a�      D   , ���a� ���b� 	���b� 	���a� ���a�      D   , ���a� ���b� ���b� ���a� ���a�      D   , ���a� ���b� ���b� ���a� ���a�      D   , ���a� ���b� ~��b� ~��a� ���a�      D   , |��a� |��b� b��b� b��a� |��a�      D   ,  ����^  ����a  ����a  ����^  ����^      D   ,  �f��^  �f��a  ����a  ����^  �f��^      D   ,  �J��^  �J��a  �p��a  �p��^  �J��^      D   ,  �.��^  �.��a  T��a  T��^  �.��^      D   , ��^ ��a 8��a 8��^ ��^      D   , ���^ ���a ��a ��^ ���^      D   , ���^ ���a 	 ��a 	 ��^ ���^      D   , 	���^ 	���a ���a ���^ 	���^      D   , ���^ ���a ���a ���^ ���^      D   , ���^ ���a ���a ���^ ���^      D   , j��^ j��a ���a ���^ j��^      D   ,  ����a�  ����b�  ����b�  ����a�  ����a�      D   ,  ����\�  ����]{  ����]{  ����\�  ����\�      D   ,  ����\�  ����]{  �z��]{  �z��\�  ����\�      D   ,  �x��\�  �x��]{  �^��]{  �^��\�  �x��\�      D   ,  �\��\�  �\��]{  �B��]{  �B��\�  �\��\�      D   ,  @��\�  @��]{ &��]{ &��\�  @��\�      D   , $��\� $��]{ 
��]{ 
��\� $��\�      D   , ��\� ��]{ ���]{ ���\� ��\�      D   , ���\� ���]{ 	���]{ 	���\� ���\�      D   , ���\� ���]{ ���]{ ���\� ���\�      D   , ���\� ���]{ ���]{ ���\� ���\�      D   , ���\� ���]{ ~��]{ ~��\� ���\�      D   , |��\� |��]{ b��]{ b��\� |��\�      D   ,  �o��L7  �o��\�  ����\�  ����L7  �o��L7      D   ,  �S��L7  �S��\�  ����\�  ����L7  �S��L7      D   ,  �7��L7  �7��\�  ����\�  ����L7  �7��L7      D   ,  ���L7  ���\�  ����\�  ����L7  ���L7      D   ,  ����L7  ����\� g��\� g��L7  ����L7      D   , ���L7 ���\� K��\� K��L7 ���L7      D   , ���L7 ���\� /��\� /��L7 ���L7      D   , ���L7 ���\� 
��\� 
��L7 ���L7      D   , ���L7 ���\� ���\� ���L7 ���L7      D   , s��L7 s��\� ���\� ���L7 s��L7      D   , W��L7 W��\� ���\� ���L7 W��L7      D   , ;��L7 ;��\� ���\� ���L7 ;��L7      D   ,  ����K�  ����L7  ����L7  ����K�  ����K�      D   ,  ����K�  ����L7  �z��L7  �z��K�  ����K�      D   ,  �x��K�  �x��L7  �^��L7  �^��K�  �x��K�      D   ,  �\��K�  �\��L7  �B��L7  �B��K�  �\��K�      D   ,  @��K�  @��L7 &��L7 &��K�  @��K�      D   , $��K� $��L7 
��L7 
��K� $��K�      D   , ��K� ��L7 ���L7 ���K� ��K�      D   , ���K� ���L7 	���L7 	���K� ���K�      D   , ���K� ���L7 ���L7 ���K� ���K�      D   , ���K� ���L7 ���L7 ���K� ���K�      D   , ���K� ���L7 ~��L7 ~��K� ���K�      D   , |��K� |��L7 b��L7 b��K� |��K�      D   , |K��b� |K��s }���s }���b� |K��b�      D   , zz��^ zz��a |���a |���^ zz��^      D   , |K��L7 |K��\� }���\� }���L7 |K��L7      D   , ��b� ��s ���s ���b� ��b�      D   , ��b� ��s k��s k��b� ��b�      D   , ���b� ���s O��s O��b� ���b�      D   , ���b� ���s !3��s !3��b� ���b�      D   , "���b� "���s $��s $��b� "���b�      D   , %���b� %���s &���s &���b� %���b�      D   , (w��b� (w��s )���s )���b� (w��b�      D   , +[��b� +[��s ,���s ,���b� +[��b�      D   , .?��b� .?��s /���s /���b� .?��b�      D   , 1#��b� 1#��s 2���s 2���b� 1#��b�      D   , 4��b� 4��s 5o��s 5o��b� 4��b�      D   , 6���b� 6���s 8S��s 8S��b� 6���b�      D   , 9���b� 9���s ;7��s ;7��b� 9���b�      D   , <���b� <���s >��s >��b� <���b�      D   , ?���b� ?���s @���s @���b� ?���b�      D   , B{��b� B{��s C���s C���b� B{��b�      D   , E_��b� E_��s F���s F���b� E_��b�      D   , HC��b� HC��s I���s I���b� HC��b�      D   , K'��b� K'��s L���s L���b� K'��b�      D   , N��b� N��s Os��s Os��b� N��b�      D   , P���b� P���s RW��s RW��b� P���b�      D   , S���b� S���s U;��s U;��b� S���b�      D   , V���b� V���s X��s X��b� V���b�      D   , Y���b� Y���s [��s [��b� Y���b�      D   , \��b� \��s ]���s ]���b� \��b�      D   , _c��b� _c��s `���s `���b� _c��b�      D   , bG��b� bG��s c���s c���b� bG��b�      D   , e+��b� e+��s f���s f���b� e+��b�      D   , h��b� h��s iw��s iw��b� h��b�      D   , j���b� j���s l[��s l[��b� j���b�      D   , m���b� m���s o?��s o?��b� m���b�      D   , p���b� p���s r#��s r#��b� p���b�      D   , s���b� s���s u��s u��b� s���b�      D   , v���b� v���s w���s w���b� v���b�      D   , yg��b� yg��s z���s z���b� yg��b�      D   , IV��^ IV��a K|��a K|��^ IV��^      D   , HC��L7 HC��\� I���\� I���L7 HC��L7      D   , Q0��s Q0��sQ R��sQ R��s Q0��s      D   , T��s T��sQ T���sQ T���s T��s      D   , V���s V���sQ W���sQ W���s V���s      D   , Y���s Y���sQ Z���sQ Z���s Y���s      D   , \���s \���sQ ]���sQ ]���s \���s      D   , _���s _���sQ `���sQ `���s _���s      D   , b���s b���sQ cn��sQ cn��s b���s      D   , el��s el��sQ fR��sQ fR��s el��s      D   , hP��s hP��sQ i6��sQ i6��s hP��s      D   , k4��s k4��sQ l��sQ l��s k4��s      D   , n��s n��sQ n���sQ n���s n��s      D   , p���s p���sQ q���sQ q���s p���s      D   , s���s s���sQ t���sQ t���s s���s      D   , v���s v���sQ w���sQ w���s v���s      D   , y���s y���sQ z���sQ z���s y���s      D   , Kh��s Kh��sQ LN��sQ LN��s Kh��s      D   , NL��s NL��sQ O2��sQ O2��s NL��s      D   , E���s E���sQ F���sQ F���s E���s      D   , H���s H���sQ Ij��sQ Ij��s H���s      D   , 1d��s 1d��sQ 2J��sQ 2J��s 1d��s      D   , :��s :��sQ :���sQ :���s :��s      D   , <���s <���sQ =���sQ =���s <���s      D   , ?���s ?���sQ @���sQ @���s ?���s      D   , 4H��s 4H��sQ 5.��sQ 5.��s 4H��s      D   , B���s B���sQ C���sQ C���s B���s      D   , 7,��s 7,��sQ 8��sQ 8��s 7,��s      D   , `��s `��sQ F��sQ F��s `��s      D   , D��s D��sQ *��sQ *��s D��s      D   , (��s (��sQ ��sQ ��s (��s      D   ,  ��s  ��sQ  ���sQ  ���s  ��s      D   , "���s "���sQ #���sQ #���s "���s      D   , %���s %���sQ &���sQ &���s %���s      D   , (���s (���sQ )���sQ )���s (���s      D   , +���s +���sQ ,���sQ ,���s +���s      D   , .���s .���sQ /f��sQ /f��s .���s      D   , (���a� (���b� )���b� )���a� (���a�      D   , +���a� +���b� ,���b� ,���a� +���a�      D   , .���a� .���b� /f��b� /f��a� .���a�      D   , 1d��a� 1d��b� 2J��b� 2J��a� 1d��a�      D   , 4H��a� 4H��b� 5.��b� 5.��a� 4H��a�      D   , 2��^ 2��a X��a X��^ 2��^      D   , ��^ ��a <��a <��^ ��^      D   , ���^ ���a   ��a   ��^ ���^      D   ,  ���^  ���a #��a #��^  ���^      D   , #���^ #���a %���a %���^ #���^      D   , &���^ &���a (���a (���^ &���^      D   , )���^ )���a +���a +���^ )���^      D   , ,n��^ ,n��a .���a .���^ ,n��^      D   , /R��^ /R��a 1x��a 1x��^ /R��^      D   , 26��^ 26��a 4\��a 4\��^ 26��^      D   , 5��^ 5��a 7@��a 7@��^ 5��^      D   , 7���^ 7���a :$��a :$��^ 7���^      D   , :���^ :���a =��a =��^ :���^      D   , =���^ =���a ?���a ?���^ =���^      D   , @���^ @���a B���a B���^ @���^      D   , C���^ C���a E���a E���^ C���^      D   , Fr��^ Fr��a H���a H���^ Fr��^      D   , 7,��a� 7,��b� 8��b� 8��a� 7,��a�      D   , :��a� :��b� :���b� :���a� :��a�      D   , `��\� `��]{ F��]{ F��\� `��\�      D   , D��\� D��]{ *��]{ *��\� D��\�      D   , (��\� (��]{ ��]{ ��\� (��\�      D   ,  ��\�  ��]{  ���]{  ���\�  ��\�      D   , "���\� "���]{ #���]{ #���\� "���\�      D   , %���\� %���]{ &���]{ &���\� %���\�      D   , (���\� (���]{ )���]{ )���\� (���\�      D   , +���\� +���]{ ,���]{ ,���\� +���\�      D   , .���\� .���]{ /f��]{ /f��\� .���\�      D   , 1d��\� 1d��]{ 2J��]{ 2J��\� 1d��\�      D   , 4H��\� 4H��]{ 5.��]{ 5.��\� 4H��\�      D   , 7,��\� 7,��]{ 8��]{ 8��\� 7,��\�      D   , :��\� :��]{ :���]{ :���\� :��\�      D   , <���\� <���]{ =���]{ =���\� <���\�      D   , ?���\� ?���]{ @���]{ @���\� ?���\�      D   , B���\� B���]{ C���]{ C���\� B���\�      D   , E���\� E���]{ F���]{ F���\� E���\�      D   , H���\� H���]{ Ij��]{ Ij��\� H���\�      D   , ��L7 ��\� ���\� ���L7 ��L7      D   , ��L7 ��\� k��\� k��L7 ��L7      D   , ���L7 ���\� O��\� O��L7 ���L7      D   , ���L7 ���\� !3��\� !3��L7 ���L7      D   , "���L7 "���\� $��\� $��L7 "���L7      D   , %���L7 %���\� &���\� &���L7 %���L7      D   , (w��L7 (w��\� )���\� )���L7 (w��L7      D   , +[��L7 +[��\� ,���\� ,���L7 +[��L7      D   , .?��L7 .?��\� /���\� /���L7 .?��L7      D   , 1#��L7 1#��\� 2���\� 2���L7 1#��L7      D   , 4��L7 4��\� 5o��\� 5o��L7 4��L7      D   , 6���L7 6���\� 8S��\� 8S��L7 6���L7      D   , 9���L7 9���\� ;7��\� ;7��L7 9���L7      D   , <���L7 <���\� >��\� >��L7 <���L7      D   , ?���L7 ?���\� @���\� @���L7 ?���L7      D   , B{��L7 B{��\� C���\� C���L7 B{��L7      D   , E_��L7 E_��\� F���\� F���L7 E_��L7      D   , <���a� <���b� =���b� =���a� <���a�      D   , ?���a� ?���b� @���b� @���a� ?���a�      D   , B���a� B���b� C���b� C���a� B���a�      D   , E���a� E���b� F���b� F���a� E���a�      D   , H���a� H���b� Ij��b� Ij��a� H���a�      D   , `��a� `��b� F��b� F��a� `��a�      D   , D��a� D��b� *��b� *��a� D��a�      D   , (��a� (��b� ��b� ��a� (��a�      D   ,  ��a�  ��b�  ���b�  ���a�  ��a�      D   , "���a� "���b� #���b� #���a� "���a�      D   , %���a� %���b� &���b� &���a� %���a�      D   , `��K� `��L7 F��L7 F��K� `��K�      D   , D��K� D��L7 *��L7 *��K� D��K�      D   , (��K� (��L7 ��L7 ��K� (��K�      D   ,  ��K�  ��L7  ���L7  ���K�  ��K�      D   , "���K� "���L7 #���L7 #���K� "���K�      D   , %���K� %���L7 &���L7 &���K� %���K�      D   , (���K� (���L7 )���L7 )���K� (���K�      D   , +���K� +���L7 ,���L7 ,���K� +���K�      D   , .���K� .���L7 /f��L7 /f��K� .���K�      D   , 1d��K� 1d��L7 2J��L7 2J��K� 1d��K�      D   , 4H��K� 4H��L7 5.��L7 5.��K� 4H��K�      D   , 7,��K� 7,��L7 8��L7 8��K� 7,��K�      D   , :��K� :��L7 :���L7 :���K� :��K�      D   , <���K� <���L7 =���L7 =���K� <���K�      D   , ?���K� ?���L7 @���L7 @���K� ?���K�      D   , B���K� B���L7 C���L7 C���K� B���K�      D   , E���K� E���L7 F���L7 F���K� E���K�      D   , H���K� H���L7 Ij��L7 Ij��K� H���K�      D   , p���\� p���]{ q���]{ q���\� p���\�      D   , s���\� s���]{ t���]{ t���\� s���\�      D   , v���\� v���]{ w���]{ w���\� v���\�      D   , y���\� y���]{ z���]{ z���\� y���\�      D   , R��^ R��a T(��a T(��^ R��^      D   , T���^ T���a W��a W��^ T���^      D   , W���^ W���a Y���a Y���^ W���^      D   , Z���^ Z���a \���a \���^ Z���^      D   , ]���^ ]���a _���a _���^ ]���^      D   , `v��^ `v��a b���a b���^ `v��^      D   , cZ��^ cZ��a e���a e���^ cZ��^      D   , f>��^ f>��a hd��a hd��^ f>��^      D   , i"��^ i"��a kH��a kH��^ i"��^      D   , l��^ l��a n,��a n,��^ l��^      D   , n���^ n���a q��a q��^ n���^      D   , q���^ q���a s���a s���^ q���^      D   , t���^ t���a v���a v���^ t���^      D   , w���^ w���a y���a y���^ w���^      D   , n��a� n��b� n���b� n���a� n��a�      D   , p���a� p���b� q���b� q���a� p���a�      D   , s���a� s���b� t���b� t���a� s���a�      D   , v���a� v���b� w���b� w���a� v���a�      D   , K'��L7 K'��\� L���\� L���L7 K'��L7      D   , N��L7 N��\� Os��\� Os��L7 N��L7      D   , P���L7 P���\� RW��\� RW��L7 P���L7      D   , S���L7 S���\� U;��\� U;��L7 S���L7      D   , V���L7 V���\� X��\� X��L7 V���L7      D   , Y���L7 Y���\� [��\� [��L7 Y���L7      D   , \��L7 \��\� ]���\� ]���L7 \��L7      D   , _c��L7 _c��\� `���\� `���L7 _c��L7      D   , bG��L7 bG��\� c���\� c���L7 bG��L7      D   , e+��L7 e+��\� f���\� f���L7 e+��L7      D   , h��L7 h��\� iw��\� iw��L7 h��L7      D   , j���L7 j���\� l[��\� l[��L7 j���L7      D   , m���L7 m���\� o?��\� o?��L7 m���L7      D   , p���L7 p���\� r#��\� r#��L7 p���L7      D   , s���L7 s���\� u��\� u��L7 s���L7      D   , v���L7 v���\� w���\� w���L7 v���L7      D   , yg��L7 yg��\� z���\� z���L7 yg��L7      D   , y���a� y���b� z���b� z���a� y���a�      D   , Kh��a� Kh��b� LN��b� LN��a� Kh��a�      D   , NL��a� NL��b� O2��b� O2��a� NL��a�      D   , Q0��a� Q0��b� R��b� R��a� Q0��a�      D   , T��a� T��b� T���b� T���a� T��a�      D   , V���a� V���b� W���b� W���a� V���a�      D   , Y���a� Y���b� Z���b� Z���a� Y���a�      D   , \���a� \���b� ]���b� ]���a� \���a�      D   , _���a� _���b� `���b� `���a� _���a�      D   , b���a� b���b� cn��b� cn��a� b���a�      D   , el��a� el��b� fR��b� fR��a� el��a�      D   , hP��a� hP��b� i6��b� i6��a� hP��a�      D   , k4��a� k4��b� l��b� l��a� k4��a�      D   , L:��^ L:��a N`��a N`��^ L:��^      D   , O��^ O��a QD��a QD��^ O��^      D   , Kh��\� Kh��]{ LN��]{ LN��\� Kh��\�      D   , NL��\� NL��]{ O2��]{ O2��\� NL��\�      D   , Q0��\� Q0��]{ R��]{ R��\� Q0��\�      D   , T��\� T��]{ T���]{ T���\� T��\�      D   , V���\� V���]{ W���]{ W���\� V���\�      D   , Y���\� Y���]{ Z���]{ Z���\� Y���\�      D   , \���\� \���]{ ]���]{ ]���\� \���\�      D   , _���\� _���]{ `���]{ `���\� _���\�      D   , b���\� b���]{ cn��]{ cn��\� b���\�      D   , el��\� el��]{ fR��]{ fR��\� el��\�      D   , hP��\� hP��]{ i6��]{ i6��\� hP��\�      D   , k4��\� k4��]{ l��]{ l��\� k4��\�      D   , n��\� n��]{ n���]{ n���\� n��\�      D   , Kh��K� Kh��L7 LN��L7 LN��K� Kh��K�      D   , NL��K� NL��L7 O2��L7 O2��K� NL��K�      D   , Q0��K� Q0��L7 R��L7 R��K� Q0��K�      D   , T��K� T��L7 T���L7 T���K� T��K�      D   , V���K� V���L7 W���L7 W���K� V���K�      D   , Y���K� Y���L7 Z���L7 Z���K� Y���K�      D   , \���K� \���L7 ]���L7 ]���K� \���K�      D   , _���K� _���L7 `���L7 `���K� _���K�      D   , b���K� b���L7 cn��L7 cn��K� b���K�      D   , el��K� el��L7 fR��L7 fR��K� el��K�      D   , hP��K� hP��L7 i6��L7 i6��K� hP��K�      D   , k4��K� k4��L7 l��L7 l��K� k4��K�      D   , n��K� n��L7 n���L7 n���K� n��K�      D   , p���K� p���L7 q���L7 q���K� p���K�      D   , s���K� s���L7 t���L7 t���K� s���K�      D   , v���K� v���L7 w���L7 w���K� v���K�      D   , y���K� y���L7 z���L7 z���K� y���K�      D   , �;��b� �;��s Σ��s Σ��b� �;��b�      D   , /��b� /��s ����s ����b� /��b�      D   , ���b� ���s �{��s �{��b� ���b�      D   , ����b� ����s �_��s �_��b� ����b�      D   , ����b� ����s �C��s �C��b� ����b�      D   , ����b� ����s �'��s �'��b� ����b�      D   , ����b� ����s ���s ���b� ����b�      D   , ����b� ����s ����s ����b� ����b�      D   , �k��b� �k��s ����s ����b� �k��b�      D   , �O��b� �O��s ����s ����b� �O��b�      D   , �3��b� �3��s ����s ����b� �3��b�      D   , ���b� ���s ���s ���b� ���b�      D   , ����b� ����s �c��s �c��b� ����b�      D   , ����b� ����s �G��s �G��b� ����b�      D   , ����b� ����s �+��s �+��b� ����b�      D   , ����b� ����s ���s ���b� ����b�      D   , ����b� ����s ����s ����b� ����b�      D   , �o��b� �o��s ����s ����b� �o��b�      D   , �S��b� �S��s ����s ����b� �S��b�      D   , �7��b� �7��s ����s ����b� �7��b�      D   , ҟ��Z ҟ��ji ���ji ���Z ҟ��Z      D   , ���Z ���ji �l��ji �l��Z ���Z      D   , �~��Y� �~��j( ����j( ����Y� �~��Y�      D   , ����^ ����a ����a ����^ ����^      D   , ���b� ���s ����s ����b� ���b�      D   , ����b� ����s �g��s �g��b� ����b�      D   , ����b� ����s �K��s �K��b� ����b�      D   , ����b� ����s �/��s �/��b� ����b�      D   , ����b� ����s ���s ���b� ����b�      D   , ď��b� ď��s ����s ����b� ď��b�      D   , �s��b� �s��s ����s ����b� �s��b�      D   , �W��b� �W��s ˿��s ˿��b� �W��b�      D   , �|��s �|��sQ �b��sQ �b��s �|��s      D   , ����s ����sQ �z��sQ �z��s ����s      D   , �x��s �x��sQ �^��sQ �^��s �x��s      D   , �\��s �\��sQ �B��sQ �B��s �\��s      D   , �@��s �@��sQ �&��sQ �&��s �@��s      D   , �$��s �$��sQ �
��sQ �
��s �$��s      D   , ���s ���sQ ����sQ ����s ���s      D   , ����s ����sQ ����sQ ����s ����s      D   , ����s ����sQ Ŷ��sQ Ŷ��s ����s      D   , Ǵ��s Ǵ��sQ Ț��sQ Ț��s Ǵ��s      D   , �8��s �8��sQ ���sQ ���s �8��s      D   , ���s ���sQ ���sQ ���s ���s      D   , � ��s � ��sQ ����sQ ����s � ��s      D   , ����s ����sQ ����sQ ����s ����s      D   , ����s ����sQ ����sQ ����s ����s      D   , ����s ����sQ ����sQ ����s ����s      D   , ����s ����sQ �v��sQ �v��s ����s      D   , �t��s �t��sQ �Z��sQ �Z��s �t��s      D   , �X��s �X��sQ �>��sQ �>��s �X��s      D   , �<��s �<��sQ �"��sQ �"��s �<��s      D   , |���s |���sQ }r��sQ }r��s |���s      D   , � ��s � ��sQ ���sQ ���s � ��s      D   , ���s ���sQ ����sQ ����s ���s      D   , ����s ����sQ ����sQ ����s ����s      D   , ����s ����sQ ����sQ ����s ����s      D   , ����s ����sQ ����sQ ����s ����s      D   , p��s p��sQ �V��sQ �V��s p��s      D   , �T��s �T��sQ �:��sQ �:��s �T��s      D   , ����a� ����b� �v��b� �v��a� ����a�      D   , �t��a� �t��b� �Z��b� �Z��a� �t��a�      D   , �X��a� �X��b� �>��b� �>��a� �X��a�      D   , �<��a� �<��b� �"��b� �"��a� �<��a�      D   , � ��a� � ��b� ���b� ���a� � ��a�      D   , ���a� ���b� ����b� ����a� ���a�      D   , ����a� ����b� ����b� ����a� ����a�      D   , ����a� ����b� ����b� ����a� ����a�      D   , ����a� ����b� ����b� ����a� ����a�      D   , }^��^ }^��a ���a ���^ }^��^      D   , �B��^ �B��a �h��a �h��^ �B��^      D   , �&��^ �&��a �L��a �L��^ �&��^      D   , �
��^ �
��a �0��a �0��^ �
��^      D   , ����^ ����a ���a ���^ ����^      D   , ����^ ����a ����a ����^ ����^      D   , ����^ ����a ����a ����^ ����^      D   , ����^ ����a ����a ����^ ����^      D   , �~��^ �~��a ����a ����^ �~��^      D   , �b��^ �b��a ����a ����^ �b��^      D   , �F��^ �F��a �l��a �l��^ �F��^      D   , �*��^ �*��a �P��a �P��^ �*��^      D   , ���^ ���a �4��a �4��^ ���^      D   , ����^ ����a ���a ���^ ����^      D   , /��L7 /��\� ����\� ����L7 /��L7      D   , ���L7 ���\� �{��\� �{��L7 ���L7      D   , ����L7 ����\� �_��\� �_��L7 ����L7      D   , ����L7 ����\� �C��\� �C��L7 ����L7      D   , ����L7 ����\� �'��\� �'��L7 ����L7      D   , ����L7 ����\� ���\� ���L7 ����L7      D   , ����L7 ����\� ����\� ����L7 ����L7      D   , �k��L7 �k��\� ����\� ����L7 �k��L7      D   , �O��L7 �O��\� ����\� ����L7 �O��L7      D   , �3��L7 �3��\� ����\� ����L7 �3��L7      D   , ���L7 ���\� ���\� ���L7 ���L7      D   , ����L7 ����\� �c��\� �c��L7 ����L7      D   , ����L7 ����\� �G��\� �G��L7 ����L7      D   , ����L7 ����\� �+��\� �+��L7 ����L7      D   , ����L7 ����\� ���\� ���L7 ����L7      D   , ����L7 ����\� ����\� ����L7 ����L7      D   , �o��L7 �o��\� ����\� ����L7 �o��L7      D   , ����\� ����]{ ����]{ ����\� ����\�      D   , ����\� ����]{ ����]{ ����\� ����\�      D   , |���\� |���]{ }r��]{ }r��\� |���\�      D   , p��\� p��]{ �V��]{ �V��\� p��\�      D   , �T��\� �T��]{ �:��]{ �:��\� �T��\�      D   , �8��\� �8��]{ ���]{ ���\� �8��\�      D   , ����^ ����a ����a ����^ ����^      D   , ����^ ����a ����a ����^ ����^      D   , ����^ ����a ����a ����^ ����^      D   , ���\� ���]{ ���]{ ���\� ���\�      D   , � ��\� � ��]{ ����]{ ����\� � ��\�      D   , ����\� ����]{ ����]{ ����\� ����\�      D   , ����\� ����]{ ����]{ ����\� ����\�      D   , ����\� ����]{ ����]{ ����\� ����\�      D   , ����\� ����]{ �v��]{ �v��\� ����\�      D   , �t��\� �t��]{ �Z��]{ �Z��\� �t��\�      D   , �X��\� �X��]{ �>��]{ �>��\� �X��\�      D   , �<��\� �<��]{ �"��]{ �"��\� �<��\�      D   , � ��\� � ��]{ ���]{ ���\� � ��\�      D   , ���\� ���]{ ����]{ ����\� ���\�      D   , ����\� ����]{ ����]{ ����\� ����\�      D   , |���a� |���b� }r��b� }r��a� |���a�      D   , p��a� p��b� �V��b� �V��a� p��a�      D   , �T��a� �T��b� �:��b� �:��a� �T��a�      D   , �8��a� �8��b� ���b� ���a� �8��a�      D   , ���a� ���b� ���b� ���a� ���a�      D   , � ��a� � ��b� ����b� ����a� � ��a�      D   , ����a� ����b� ����b� ����a� ����a�      D   , ����a� ����b� ����b� ����a� ����a�      D   , ����a� ����b� ����b� ����a� ����a�      D   , |���K� |���L7 }r��L7 }r��K� |���K�      D   , p��K� p��L7 �V��L7 �V��K� p��K�      D   , �T��K� �T��L7 �:��L7 �:��K� �T��K�      D   , �8��K� �8��L7 ���L7 ���K� �8��K�      D   , ���K� ���L7 ���L7 ���K� ���K�      D   , � ��K� � ��L7 ����L7 ����K� � ��K�      D   , ����K� ����L7 ����L7 ����K� ����K�      D   , ����K� ����L7 ����L7 ����K� ����K�      D   , ����K� ����L7 ����L7 ����K� ����K�      D   , ����K� ����L7 �v��L7 �v��K� ����K�      D   , �t��K� �t��L7 �Z��L7 �Z��K� �t��K�      D   , �X��K� �X��L7 �>��L7 �>��K� �X��K�      D   , �<��K� �<��L7 �"��L7 �"��K� �<��K�      D   , � ��K� � ��L7 ���L7 ���K� � ��K�      D   , ���K� ���L7 ����L7 ����K� ���K�      D   , ����K� ����L7 ����L7 ����K� ����K�      D   , ����K� ����L7 ����L7 ����K� ����K�      D   , ����K� ����L7 ����L7 ����K� ����K�      D   , �W��L7 �W��\� ˿��\� ˿��L7 �W��L7      D   , �;��L7 �;��\� Σ��\� Σ��L7 �;��L7      D   , �\��\� �\��]{ �B��]{ �B��\� �\��\�      D   , �@��\� �@��]{ �&��]{ �&��\� �@��\�      D   , ����a� ����b� �z��b� �z��a� ����a�      D   , �x��a� �x��b� �^��b� �^��a� �x��a�      D   , �\��a� �\��b� �B��b� �B��a� �\��a�      D   , �@��a� �@��b� �&��b� �&��a� �@��a�      D   , �$��a� �$��b� �
��b� �
��a� �$��a�      D   , ���a� ���b� ����b� ����a� ���a�      D   , ����a� ����b� ����b� ����a� ����a�      D   , ����a� ����b� Ŷ��b� Ŷ��a� ����a�      D   , Ǵ��a� Ǵ��b� Ț��b� Ț��a� Ǵ��a�      D   , �|��a� �|��b� �b��b� �b��a� �|��a�      D   , �$��\� �$��]{ �
��]{ �
��\� �$��\�      D   , ���\� ���]{ ����]{ ����\� ���\�      D   , ����\� ����]{ ����]{ ����\� ����\�      D   , ����\� ����]{ Ŷ��]{ Ŷ��\� ����\�      D   , Ǵ��\� Ǵ��]{ Ț��]{ Ț��\� Ǵ��\�      D   , ����\� ����]{ �z��]{ �z��\� ����\�      D   , �x��\� �x��]{ �^��]{ �^��\� �x��\�      D   , �S��L7 �S��\� ����\� ����L7 �S��L7      D   , �f��^ �f��a ����a ����^ �f��^      D   , �J��^ �J��a �p��a �p��^ �J��^      D   , �.��^ �.��a �T��a �T��^ �.��^      D   , ���^ ���a �8��a �8��^ ���^      D   , ����^ ����a ���a ���^ ����^      D   , ����^ ����a � ��a � ��^ ����^      D   , ¾��^ ¾��a ����a ����^ ¾��^      D   , Ţ��^ Ţ��a ����a ����^ Ţ��^      D   , Ȇ��^ Ȇ��a ʬ��a ʬ��^ Ȇ��^      D   , �j��^ �j��a ͐��a ͐��^ �j��^      D   , �7��L7 �7��\� ����\� ����L7 �7��L7      D   , ���L7 ���\� ����\� ����L7 ���L7      D   , ����L7 ����\� �g��\� �g��L7 ����L7      D   , ����L7 ����\� �K��\� �K��L7 ����L7      D   , ����L7 ����\� �/��\� �/��L7 ����L7      D   , ����L7 ����\� ���\� ���L7 ����L7      D   , ď��L7 ď��\� ����\� ����L7 ď��L7      D   , �s��L7 �s��\� ����\� ����L7 �s��L7      D   , ����K� ����L7 �z��L7 �z��K� ����K�      D   , �x��K� �x��L7 �^��L7 �^��K� �x��K�      D   , �\��K� �\��L7 �B��L7 �B��K� �\��K�      D   , �@��K� �@��L7 �&��L7 �&��K� �@��K�      D   , �$��K� �$��L7 �
��L7 �
��K� �$��K�      D   , ���K� ���L7 ����L7 ����K� ���K�      D   , ����K� ����L7 ����L7 ����K� ����K�      D   , ����K� ����L7 Ŷ��L7 Ŷ��K� ����K�      D   , Ǵ��K� Ǵ��L7 Ț��L7 Ț��K� Ǵ��K�      @   , 1U  (2 1U  8� A�  8� A�  (2 1U  (2      @   , ��  (2 ��  8� �D  8� �D  (2 ��  (2      @   ,  �  %�  �  (  �  (  �  %�  �  %�      @   ,  ��  %�  ��  (  �!  (  �!  %�  ��  %�      @   ,  �6  $�  �6  (2  ��  (2  ��  $�  �6  $�      @   ,  ��  $�  ��  (2  ��  (2  ��  $�  ��  $�      @   ,  ��  $�  ��  (2 g  (2 g  $�  ��  $�      @   , /  $� /  (2 .:  (2 .:  $� /  $�      @   , 1U  $� 1U  (2 EF  (2 EF  $� 1U  $�      @   , F  $� F  (2 N~  (2 N~  $� F  $�      @   , OF  $� OF  (2 `�  (2 `�  $� OF  $�      @   , a�  $� a�  (2 ~�  (2 ~�  $� a�  $�      @   , ��  $� ��  (2 ��  (2 ��  $� ��  $�      @   , ��  $� ��  (2 �  (2 �  $� ��  $�      @   , ��  $� ��  (2 �u  (2 �u  $� ��  $�      @   , �=  $� �=  (2 �H  (2 �H  $� �=  $�      @   ,  [���g  [  �  ��  �  �����g  [���g      @   , 1U  # 1U  $� A�  $� A�  # 1U  #      @   , ��  # ��  $� �D  $� �D  # ��  #      @   , �c  # �c  8� ��  8� ��  # �c  #      @   ,  \���~�  \�����  bH����  bH��~�  \���~�      @   ,  [��{]  [��~�  ����~�  ����{]  [��{]      F  , , ���q� ���rR S��rR S��q� ���q�      F  , , ���o� ���p� S��p� S��o� ���o�      F  , , ���nj ���o2 S��o2 S��nj ���nj      F  , , ���l� ���m� S��m� S��l� ���l�      F  , , ���kJ ���l S��l S��kJ ���kJ      F  , , ���i� ���j� S��j� S��i� ���i�      F  , , ���h* ���h� S��h� S��h* ���h*      F  , , ���f� ���gb S��gb S��f� ���f�      F  , , ���e
 ���e� S��e� S��e
 ���e
      F  , , ���cz ���dB S��dB S��cz ���cz      F  , , ���Z� ���[� S��[� S��Z� ���Z�      F  , , ���Yf ���Z. S��Z. S��Yf ���Yf      F  , , ���W� ���X� S��X� S��W� ���W�      F  , , ���VF ���W S��W S��VF ���VF      F  , , ���T� ���U~ S��U~ S��T� ���T�      F  , , ���S& ���S� S��S� S��S& ���S&      F  , , ���Q� ���R^ S��R^ S��Q� ���Q�      F  , , ���P ���P� S��P� S��P ���P      F  , , ���Nv ���O> S��O> S��Nv ���Nv      F  , , ���L� ���M� S��M� S��L� ���L�      F  , , ��  2� ��  3� ��  3� ��  2� ��  2�      F  , , ��  1V ��  2 ��  2 ��  1V ��  1V      F  , , ��  /� ��  0� ��  0� ��  /� ��  /�      F  , , ��  .6 ��  .� ��  .� ��  .6 ��  .6      F  , , ��  ,� ��  -n ��  -n ��  ,� ��  ,�      F  , , ��  + ��  +� ��  +� ��  + ��  +      F  , , ��  )� ��  *N ��  *N ��  )� ��  )�      F  , , ��  "� ��  #Z ��  #Z ��  "� ��  "�      F  , , ��  ! ��  !� ��  !� ��  ! ��  !      F  , , ��  r ��   : ��   : ��  r ��  r      F  , , ��  � ��  � ��  � ��  � ��  �      F  , , ��  R ��   ��   ��  R ��  R      F  , , ��  � ��  � ��  � ��  � ��  �      F  , , ��  2 ��  � ��  � ��  2 ��  2      F  , , ŉ  1V ŉ  2 �Q  2 �Q  1V ŉ  1V      F  , , �%  1V �%  2 ��  2 ��  1V �%  1V      F  , , ��  1V ��  2 ω  2 ω  1V ��  1V      F  , , ŉ  /� ŉ  0� �Q  0� �Q  /� ŉ  /�      F  , , �%  /� �%  0� ��  0� ��  /� �%  /�      F  , , ��  /� ��  0� ω  0� ω  /� ��  /�      F  , , ŉ  .6 ŉ  .� �Q  .� �Q  .6 ŉ  .6      F  , , �%  .6 �%  .� ��  .� ��  .6 �%  .6      F  , , ��  .6 ��  .� ω  .� ω  .6 ��  .6      F  , , ŉ  ,� ŉ  -n �Q  -n �Q  ,� ŉ  ,�      F  , , �%  ,� �%  -n ��  -n ��  ,� �%  ,�      F  , , ��  ,� ��  -n ω  -n ω  ,� ��  ,�      F  , , ŉ  + ŉ  +� �Q  +� �Q  + ŉ  +      F  , , �%  + �%  +� ��  +� ��  + �%  +      F  , , ��  + ��  +� ω  +� ω  + ��  +      F  , , ŉ  2� ŉ  3� �Q  3� �Q  2� ŉ  2�      F  , , ŉ  )� ŉ  *N �Q  *N �Q  )� ŉ  )�      F  , , �%  )� �%  *N ��  *N ��  )� �%  )�      F  , , ��  )� ��  *N ω  *N ω  )� ��  )�      F  , , �%  2� �%  3� ��  3� ��  2� �%  2�      F  , , ��  2� ��  3� ω  3� ω  2� ��  2�      F  , , �Q  /� �Q  0� �  0� �  /� �Q  /�      F  , , �Q  2� �Q  3� �  3� �  2� �Q  2�      F  , , �}  ,� �}  -n �E  -n �E  ,� �}  ,�      F  , , �  ,� �  -n ��  -n ��  ,� �  ,�      F  , , ��  ,� ��  -n �}  -n �}  ,� ��  ,�      F  , , �Q  ,� �Q  -n �  -n �  ,� �Q  ,�      F  , , ��  ,� ��  -n ��  -n ��  ,� ��  ,�      F  , , ��  /� ��  0� ��  0� ��  /� ��  /�      F  , , ��  1V ��  2 ��  2 ��  1V ��  1V      F  , , �  2� �  3� ��  3� ��  2� �  2�      F  , , ��  2� ��  3� ��  3� ��  2� ��  2�      F  , , �}  + �}  +� �E  +� �E  + �}  +      F  , , �  + �  +� ��  +� ��  + �  +      F  , , ��  + ��  +� �}  +� �}  + ��  +      F  , , �Q  + �Q  +� �  +� �  + �Q  +      F  , , ��  + ��  +� ��  +� ��  + ��  +      F  , , �}  /� �}  0� �E  0� �E  /� �}  /�      F  , , ��  2� ��  3� �}  3� �}  2� ��  2�      F  , , �}  .6 �}  .� �E  .� �E  .6 �}  .6      F  , , �  .6 �  .� ��  .� ��  .6 �  .6      F  , , �}  )� �}  *N �E  *N �E  )� �}  )�      F  , , �  )� �  *N ��  *N ��  )� �  )�      F  , , ��  )� ��  *N �}  *N �}  )� ��  )�      F  , , �Q  )� �Q  *N �  *N �  )� �Q  )�      F  , , ��  )� ��  *N ��  *N ��  )� ��  )�      F  , , ��  .6 ��  .� �}  .� �}  .6 ��  .6      F  , , �Q  .6 �Q  .� �  .� �  .6 �Q  .6      F  , , ��  .6 ��  .� ��  .� ��  .6 ��  .6      F  , , �  /� �  0� ��  0� ��  /� �  /�      F  , , ��  /� ��  0� �}  0� �}  /� ��  /�      F  , , �}  2� �}  3� �E  3� �E  2� �}  2�      F  , , �}  1V �}  2 �E  2 �E  1V �}  1V      F  , , �  1V �  2 ��  2 ��  1V �  1V      F  , , ��  1V ��  2 �}  2 �}  1V ��  1V      F  , , �Q  1V �Q  2 �  2 �  1V �Q  1V      F  , , �}  ! �}  !� �E  !� �E  ! �}  !      F  , , �  ! �  !� ��  !� ��  ! �  !      F  , , ��  ! ��  !� �}  !� �}  ! ��  !      F  , , �Q  ! �Q  !� �  !� �  ! �Q  !      F  , , ��  ! ��  !� ��  !� ��  ! ��  !      F  , , �  "� �  #Z ��  #Z ��  "� �  "�      F  , , �}  r �}   : �E   : �E  r �}  r      F  , , �  r �   : ��   : ��  r �  r      F  , , ��  r ��   : �}   : �}  r ��  r      F  , , �Q  r �Q   : �   : �  r �Q  r      F  , , ��  r ��   : ��   : ��  r ��  r      F  , , ��  "� ��  #Z �}  #Z �}  "� ��  "�      F  , , �}  � �}  � �E  � �E  � �}  �      F  , , �  � �  � ��  � ��  � �  �      F  , , ��  � ��  � �}  � �}  � ��  �      F  , , �Q  � �Q  � �  � �  � �Q  �      F  , , ��  � ��  � ��  � ��  � ��  �      F  , , �Q  "� �Q  #Z �  #Z �  "� �Q  "�      F  , , �}  R �}   �E   �E  R �}  R      F  , , �  R �   ��   ��  R �  R      F  , , ��  R ��   �}   �}  R ��  R      F  , , �Q  R �Q   �   �  R �Q  R      F  , , ��  R ��   ��   ��  R ��  R      F  , , ��  "� ��  #Z ��  #Z ��  "� ��  "�      F  , , �}  � �}  � �E  � �E  � �}  �      F  , , �  � �  � ��  � ��  � �  �      F  , , ��  � ��  � �}  � �}  � ��  �      F  , , �Q  � �Q  � �  � �  � �Q  �      F  , , ��  � ��  � ��  � ��  � ��  �      F  , , �}  "� �}  #Z �E  #Z �E  "� �}  "�      F  , , �}  2 �}  � �E  � �E  2 �}  2      F  , , �  2 �  � ��  � ��  2 �  2      F  , , ��  2 ��  � �}  � �}  2 ��  2      F  , , �Q  2 �Q  � �  � �  2 �Q  2      F  , , ��  2 ��  � ��  � ��  2 ��  2      F  , , ŉ  R ŉ   �Q   �Q  R ŉ  R      F  , , �%  R �%   ��   ��  R �%  R      F  , , ��  R ��   ω   ω  R ��  R      F  , , ŉ  ! ŉ  !� �Q  !� �Q  ! ŉ  !      F  , , �%  ! �%  !� ��  !� ��  ! �%  !      F  , , ��  ! ��  !� ω  !� ω  ! ��  !      F  , , ŉ  � ŉ  � �Q  � �Q  � ŉ  �      F  , , �%  � �%  � ��  � ��  � �%  �      F  , , ��  � ��  � ω  � ω  � ��  �      F  , , ŉ  � ŉ  � �Q  � �Q  � ŉ  �      F  , , �%  � �%  � ��  � ��  � �%  �      F  , , ��  � ��  � ω  � ω  � ��  �      F  , , ŉ  r ŉ   : �Q   : �Q  r ŉ  r      F  , , �%  r �%   : ��   : ��  r �%  r      F  , , ��  r ��   : ω   : ω  r ��  r      F  , , ŉ  "� ŉ  #Z �Q  #Z �Q  "� ŉ  "�      F  , , �%  "� �%  #Z ��  #Z ��  "� �%  "�      F  , , ��  "� ��  #Z ω  #Z ω  "� ��  "�      F  , , ŉ  2 ŉ  � �Q  � �Q  2 ŉ  2      F  , , �%  2 �%  � ��  � ��  2 �%  2      F  , , ��  2 ��  � ω  � ω  2 ��  2      F  , , �  + �  +� ��  +� ��  + �  +      F  , , ��  + ��  +� �q  +� �q  + ��  +      F  , , �E  + �E  +� �  +� �  + �E  +      F  , , �  .6 �  .� ��  .� ��  .6 �  .6      F  , , ��  .6 ��  .� �q  .� �q  .6 ��  .6      F  , , �E  .6 �E  .� �  .� �  .6 �E  .6      F  , , y�  r y�   : zf   : zf  r y�  r      F  , , ~:  r ~:   :    :   r ~:  r      F  , , �q  r �q   : �9   : �9  r �q  r      F  , , �  r �   : ��   : ��  r �  r      F  , , ��  r ��   : �q   : �q  r ��  r      F  , , �E  r �E   : �   : �  r �E  r      F  , , y�  /� y�  0� zf  0� zf  /� y�  /�      F  , , ~:  /� ~:  0�   0�   /� ~:  /�      F  , , �q  /� �q  0� �9  0� �9  /� �q  /�      F  , , �  /� �  0� ��  0� ��  /� �  /�      F  , , ��  /� ��  0� �q  0� �q  /� ��  /�      F  , , �E  /� �E  0� �  0� �  /� �E  /�      F  , , y�  )� y�  *N zf  *N zf  )� y�  )�      F  , , ~:  )� ~:  *N   *N   )� ~:  )�      F  , , �q  )� �q  *N �9  *N �9  )� �q  )�      F  , , y�  � y�  � zf  � zf  � y�  �      F  , , ~:  � ~:  �   �   � ~:  �      F  , , �q  � �q  � �9  � �9  � �q  �      F  , , �  � �  � ��  � ��  � �  �      F  , , ��  � ��  � �q  � �q  � ��  �      F  , , �E  � �E  � �  � �  � �E  �      F  , , �  )� �  *N ��  *N ��  )� �  )�      F  , , ��  )� ��  *N �q  *N �q  )� ��  )�      F  , , �E  )� �E  *N �  *N �  )� �E  )�      F  , , �  2� �  3� ��  3� ��  2� �  2�      F  , , ��  2� ��  3� �q  3� �q  2� ��  2�      F  , , �E  2� �E  3� �  3� �  2� �E  2�      F  , , y�  ,� y�  -n zf  -n zf  ,� y�  ,�      F  , , ~:  ,� ~:  -n   -n   ,� ~:  ,�      F  , , �q  ,� �q  -n �9  -n �9  ,� �q  ,�      F  , , y�  R y�   zf   zf  R y�  R      F  , , ~:  R ~:        R ~:  R      F  , , �q  R �q   �9   �9  R �q  R      F  , , �  R �   ��   ��  R �  R      F  , , ��  R ��   �q   �q  R ��  R      F  , , �E  R �E   �   �  R �E  R      F  , , �  ,� �  -n ��  -n ��  ,� �  ,�      F  , , ��  ,� ��  -n �q  -n �q  ,� ��  ,�      F  , , �E  ,� �E  -n �  -n �  ,� �E  ,�      F  , , y�  "� y�  #Z zf  #Z zf  "� y�  "�      F  , , ~:  "� ~:  #Z   #Z   "� ~:  "�      F  , , �q  "� �q  #Z �9  #Z �9  "� �q  "�      F  , , �  "� �  #Z ��  #Z ��  "� �  "�      F  , , ��  "� ��  #Z �q  #Z �q  "� ��  "�      F  , , �E  "� �E  #Z �  #Z �  "� �E  "�      F  , , y�  � y�  � zf  � zf  � y�  �      F  , , ~:  � ~:  �   �   � ~:  �      F  , , �q  � �q  � �9  � �9  � �q  �      F  , , �  � �  � ��  � ��  � �  �      F  , , ��  � ��  � �q  � �q  � ��  �      F  , , �E  � �E  � �  � �  � �E  �      F  , , y�  1V y�  2 zf  2 zf  1V y�  1V      F  , , ~:  1V ~:  2   2   1V ~:  1V      F  , , �q  1V �q  2 �9  2 �9  1V �q  1V      F  , , �  1V �  2 ��  2 ��  1V �  1V      F  , , ��  1V ��  2 �q  2 �q  1V ��  1V      F  , , �E  1V �E  2 �  2 �  1V �E  1V      F  , , y�  .6 y�  .� zf  .� zf  .6 y�  .6      F  , , ~:  .6 ~:  .�   .�   .6 ~:  .6      F  , , �q  .6 �q  .� �9  .� �9  .6 �q  .6      F  , , y�  2 y�  � zf  � zf  2 y�  2      F  , , ~:  2 ~:  �   �   2 ~:  2      F  , , �q  2 �q  � �9  � �9  2 �q  2      F  , , �  2 �  � ��  � ��  2 �  2      F  , , ��  2 ��  � �q  � �q  2 ��  2      F  , , �E  2 �E  � �  � �  2 �E  2      F  , , y�  ! y�  !� zf  !� zf  ! y�  !      F  , , ~:  ! ~:  !�   !�   ! ~:  !      F  , , �q  ! �q  !� �9  !� �9  ! �q  !      F  , , �  ! �  !� ��  !� ��  ! �  !      F  , , ��  ! ��  !� �q  !� �q  ! ��  !      F  , , �E  ! �E  !� �  !� �  ! �E  !      F  , , y�  + y�  +� zf  +� zf  + y�  +      F  , , ~:  + ~:  +�   +�   + ~:  +      F  , , �q  + �q  +� �9  +� �9  + �q  +      F  , , y�  2� y�  3� zf  3� zf  2� y�  2�      F  , , ~:  2� ~:  3�   3�   2� ~:  2�      F  , , �q  2� �q  3� �9  3� �9  2� �q  2�      F  , , b�  /� b�  0� cZ  0� cZ  /� b�  /�      F  , , b�  ,� b�  -n cZ  -n cZ  ,� b�  ,�      F  , , g.  ,� g.  -n g�  -n g�  ,� g.  ,�      F  , , k�  ,� k�  -n l�  -n l�  ,� k�  ,�      F  , , pf  ,� pf  -n q.  -n q.  ,� pf  ,�      F  , , u  ,� u  -n u�  -n u�  ,� u  ,�      F  , , g.  /� g.  0� g�  0� g�  /� g.  /�      F  , , k�  /� k�  0� l�  0� l�  /� k�  /�      F  , , pf  /� pf  0� q.  0� q.  /� pf  /�      F  , , u  /� u  0� u�  0� u�  /� u  /�      F  , , pf  1V pf  2 q.  2 q.  1V pf  1V      F  , , u  1V u  2 u�  2 u�  1V u  1V      F  , , b�  + b�  +� cZ  +� cZ  + b�  +      F  , , g.  + g.  +� g�  +� g�  + g.  +      F  , , k�  + k�  +� l�  +� l�  + k�  +      F  , , pf  + pf  +� q.  +� q.  + pf  +      F  , , u  + u  +� u�  +� u�  + u  +      F  , , b�  1V b�  2 cZ  2 cZ  1V b�  1V      F  , , b�  )� b�  *N cZ  *N cZ  )� b�  )�      F  , , g.  )� g.  *N g�  *N g�  )� g.  )�      F  , , k�  )� k�  *N l�  *N l�  )� k�  )�      F  , , pf  )� pf  *N q.  *N q.  )� pf  )�      F  , , u  )� u  *N u�  *N u�  )� u  )�      F  , , b�  .6 b�  .� cZ  .� cZ  .6 b�  .6      F  , , g.  .6 g.  .� g�  .� g�  .6 g.  .6      F  , , k�  .6 k�  .� l�  .� l�  .6 k�  .6      F  , , pf  .6 pf  .� q.  .� q.  .6 pf  .6      F  , , u  .6 u  .� u�  .� u�  .6 u  .6      F  , , g.  1V g.  2 g�  2 g�  1V g.  1V      F  , , k�  1V k�  2 l�  2 l�  1V k�  1V      F  , , b�  2� b�  3� cZ  3� cZ  2� b�  2�      F  , , g.  2� g.  3� g�  3� g�  2� g.  2�      F  , , k�  2� k�  3� l�  3� l�  2� k�  2�      F  , , pf  2� pf  3� q.  3� q.  2� pf  2�      F  , , u  2� u  3� u�  3� u�  2� u  2�      F  , , ]�  /� ]�  0� ^�  0� ^�  /� ]�  /�      F  , , K�  /� K�  0� LN  0� LN  /� K�  /�      F  , , T�  1V T�  2 U�  2 U�  1V T�  1V      F  , , YZ  1V YZ  2 Z"  2 Z"  1V YZ  1V      F  , , ]�  1V ]�  2 ^�  2 ^�  1V ]�  1V      F  , , F�  ,� F�  -n G�  -n G�  ,� F�  ,�      F  , , F�  .6 F�  .� G�  .� G�  .6 F�  .6      F  , , K�  .6 K�  .� LN  .� LN  .6 K�  .6      F  , , P"  .6 P"  .� P�  .� P�  .6 P"  .6      F  , , T�  .6 T�  .� U�  .� U�  .6 T�  .6      F  , , YZ  .6 YZ  .� Z"  .� Z"  .6 YZ  .6      F  , , F�  )� F�  *N G�  *N G�  )� F�  )�      F  , , K�  )� K�  *N LN  *N LN  )� K�  )�      F  , , P"  )� P"  *N P�  *N P�  )� P"  )�      F  , , T�  )� T�  *N U�  *N U�  )� T�  )�      F  , , YZ  )� YZ  *N Z"  *N Z"  )� YZ  )�      F  , , ]�  )� ]�  *N ^�  *N ^�  )� ]�  )�      F  , , K�  ,� K�  -n LN  -n LN  ,� K�  ,�      F  , , P"  ,� P"  -n P�  -n P�  ,� P"  ,�      F  , , T�  ,� T�  -n U�  -n U�  ,� T�  ,�      F  , , YZ  ,� YZ  -n Z"  -n Z"  ,� YZ  ,�      F  , , ]�  ,� ]�  -n ^�  -n ^�  ,� ]�  ,�      F  , , ]�  .6 ]�  .� ^�  .� ^�  .6 ]�  .6      F  , , F�  1V F�  2 G�  2 G�  1V F�  1V      F  , , K�  1V K�  2 LN  2 LN  1V K�  1V      F  , , P"  1V P"  2 P�  2 P�  1V P"  1V      F  , , F�  + F�  +� G�  +� G�  + F�  +      F  , , K�  + K�  +� LN  +� LN  + K�  +      F  , , P"  + P"  +� P�  +� P�  + P"  +      F  , , T�  + T�  +� U�  +� U�  + T�  +      F  , , F�  /� F�  0� G�  0� G�  /� F�  /�      F  , , F�  2� F�  3� G�  3� G�  2� F�  2�      F  , , K�  2� K�  3� LN  3� LN  2� K�  2�      F  , , P"  2� P"  3� P�  3� P�  2� P"  2�      F  , , T�  2� T�  3� U�  3� U�  2� T�  2�      F  , , YZ  2� YZ  3� Z"  3� Z"  2� YZ  2�      F  , , ]�  2� ]�  3� ^�  3� ^�  2� ]�  2�      F  , , YZ  + YZ  +� Z"  +� Z"  + YZ  +      F  , , ]�  + ]�  +� ^�  +� ^�  + ]�  +      F  , , P"  /� P"  0� P�  0� P�  /� P"  /�      F  , , T�  /� T�  0� U�  0� U�  /� T�  /�      F  , , YZ  /� YZ  0� Z"  0� Z"  /� YZ  /�      F  , , K�  � K�  � LN  � LN  � K�  �      F  , , P"  � P"  � P�  � P�  � P"  �      F  , , T�  � T�  � U�  � U�  � T�  �      F  , , YZ  � YZ  � Z"  � Z"  � YZ  �      F  , , ]�  � ]�  � ^�  � ^�  � ]�  �      F  , , K�  � K�  � LN  � LN  � K�  �      F  , , P"  � P"  � P�  � P�  � P"  �      F  , , T�  � T�  � U�  � U�  � T�  �      F  , , YZ  � YZ  � Z"  � Z"  � YZ  �      F  , , ]�  � ]�  � ^�  � ^�  � ]�  �      F  , , F�  ! F�  !� G�  !� G�  ! F�  !      F  , , K�  ! K�  !� LN  !� LN  ! K�  !      F  , , P"  ! P"  !� P�  !� P�  ! P"  !      F  , , T�  ! T�  !� U�  !� U�  ! T�  !      F  , , YZ  ! YZ  !� Z"  !� Z"  ! YZ  !      F  , , ]�  ! ]�  !� ^�  !� ^�  ! ]�  !      F  , , T�  "� T�  #Z U�  #Z U�  "� T�  "�      F  , , YZ  "� YZ  #Z Z"  #Z Z"  "� YZ  "�      F  , , F�  r F�   : G�   : G�  r F�  r      F  , , F�  2 F�  � G�  � G�  2 F�  2      F  , , K�  2 K�  � LN  � LN  2 K�  2      F  , , P"  2 P"  � P�  � P�  2 P"  2      F  , , T�  2 T�  � U�  � U�  2 T�  2      F  , , YZ  2 YZ  � Z"  � Z"  2 YZ  2      F  , , ]�  2 ]�  � ^�  � ^�  2 ]�  2      F  , , K�  r K�   : LN   : LN  r K�  r      F  , , P"  r P"   : P�   : P�  r P"  r      F  , , T�  r T�   : U�   : U�  r T�  r      F  , , YZ  r YZ   : Z"   : Z"  r YZ  r      F  , , ]�  r ]�   : ^�   : ^�  r ]�  r      F  , , F�  R F�   G�   G�  R F�  R      F  , , K�  R K�   LN   LN  R K�  R      F  , , P"  R P"   P�   P�  R P"  R      F  , , T�  R T�   U�   U�  R T�  R      F  , , YZ  R YZ   Z"   Z"  R YZ  R      F  , , ]�  R ]�   ^�   ^�  R ]�  R      F  , , ]�  "� ]�  #Z ^�  #Z ^�  "� ]�  "�      F  , , F�  "� F�  #Z G�  #Z G�  "� F�  "�      F  , , K�  "� K�  #Z LN  #Z LN  "� K�  "�      F  , , P"  "� P"  #Z P�  #Z P�  "� P"  "�      F  , , F�  � F�  � G�  � G�  � F�  �      F  , , F�  � F�  � G�  � G�  � F�  �      F  , , pf  � pf  � q.  � q.  � pf  �      F  , , u  � u  � u�  � u�  � u  �      F  , , b�  R b�   cZ   cZ  R b�  R      F  , , g.  R g.   g�   g�  R g.  R      F  , , k�  R k�   l�   l�  R k�  R      F  , , pf  R pf   q.   q.  R pf  R      F  , , u  R u   u�   u�  R u  R      F  , , b�  r b�   : cZ   : cZ  r b�  r      F  , , g.  r g.   : g�   : g�  r g.  r      F  , , k�  r k�   : l�   : l�  r k�  r      F  , , pf  r pf   : q.   : q.  r pf  r      F  , , u  r u   : u�   : u�  r u  r      F  , , b�  "� b�  #Z cZ  #Z cZ  "� b�  "�      F  , , b�  2 b�  � cZ  � cZ  2 b�  2      F  , , g.  2 g.  � g�  � g�  2 g.  2      F  , , k�  2 k�  � l�  � l�  2 k�  2      F  , , pf  2 pf  � q.  � q.  2 pf  2      F  , , u  2 u  � u�  � u�  2 u  2      F  , , g.  "� g.  #Z g�  #Z g�  "� g.  "�      F  , , k�  "� k�  #Z l�  #Z l�  "� k�  "�      F  , , pf  "� pf  #Z q.  #Z q.  "� pf  "�      F  , , u  "� u  #Z u�  #Z u�  "� u  "�      F  , , b�  ! b�  !� cZ  !� cZ  ! b�  !      F  , , b�  � b�  � cZ  � cZ  � b�  �      F  , , g.  � g.  � g�  � g�  � g.  �      F  , , k�  � k�  � l�  � l�  � k�  �      F  , , pf  � pf  � q.  � q.  � pf  �      F  , , u  � u  � u�  � u�  � u  �      F  , , g.  ! g.  !� g�  !� g�  ! g.  !      F  , , k�  ! k�  !� l�  !� l�  ! k�  !      F  , , pf  ! pf  !� q.  !� q.  ! pf  !      F  , , u  ! u  !� u�  !� u�  ! u  !      F  , , b�  � b�  � cZ  � cZ  � b�  �      F  , , g.  � g.  � g�  � g�  � g.  �      F  , , k�  � k�  � l�  � l�  � k�  �      F  , , �  � �  � o  � o  � �  �      F  , , C  � C  �   �   � C  �      F  , , �  � �  �  �  �  �  � �  �      F  , , ${  � ${  � %C  � %C  � ${  �      F  , , )  � )  � )�  � )�  � )  �      F  , , -�  � -�  � .{  � .{  � -�  �      F  , , -�  ,� -�  -n .{  -n .{  ,� -�  ,�      F  , , �  ,� �  -n o  -n o  ,� �  ,�      F  , , C  ,� C  -n   -n   ,� C  ,�      F  , , �  ,� �  -n  �  -n  �  ,� �  ,�      F  , , �  ! �  !� o  !� o  ! �  !      F  , , C  ! C  !�   !�   ! C  !      F  , , �  ! �  !�  �  !�  �  ! �  !      F  , , ${  ! ${  !� %C  !� %C  ! ${  !      F  , , )  ! )  !� )�  !� )�  ! )  !      F  , , -�  ! -�  !� .{  !� .{  ! -�  !      F  , , C  1V C  2   2   1V C  1V      F  , , -�  )� -�  *N .{  *N .{  )� -�  )�      F  , , �  1V �  2  �  2  �  1V �  1V      F  , , ${  1V ${  2 %C  2 %C  1V ${  1V      F  , , )  1V )  2 )�  2 )�  1V )  1V      F  , , -�  1V -�  2 .{  2 .{  1V -�  1V      F  , , ${  ,� ${  -n %C  -n %C  ,� ${  ,�      F  , , �  1V �  2 o  2 o  1V �  1V      F  , , �  r �   : o   : o  r �  r      F  , , �  + �  +� o  +� o  + �  +      F  , , C  + C  +�   +�   + C  +      F  , , �  .6 �  .� o  .� o  .6 �  .6      F  , , �  R �   o   o  R �  R      F  , , C  R C        R C  R      F  , , �  R �    �    �  R �  R      F  , , ${  R ${   %C   %C  R ${  R      F  , , �  2 �  � o  � o  2 �  2      F  , , C  2 C  �   �   2 C  2      F  , , �  2 �  �  �  �  �  2 �  2      F  , , ${  2 ${  � %C  � %C  2 ${  2      F  , , )  2 )  � )�  � )�  2 )  2      F  , , -�  2 -�  � .{  � .{  2 -�  2      F  , , )  R )   )�   )�  R )  R      F  , , -�  R -�   .{   .{  R -�  R      F  , , �  + �  +�  �  +�  �  + �  +      F  , , ${  + ${  +� %C  +� %C  + ${  +      F  , , )  + )  +� )�  +� )�  + )  +      F  , , -�  + -�  +� .{  +� .{  + -�  +      F  , , C  r C   :    :   r C  r      F  , , �  � �  � o  � o  � �  �      F  , , C  � C  �   �   � C  �      F  , , �  � �  �  �  �  �  � �  �      F  , , ${  � ${  � %C  � %C  � ${  �      F  , , )  � )  � )�  � )�  � )  �      F  , , -�  � -�  � .{  � .{  � -�  �      F  , , C  .6 C  .�   .�   .6 C  .6      F  , , �  .6 �  .�  �  .�  �  .6 �  .6      F  , , ${  .6 ${  .� %C  .� %C  .6 ${  .6      F  , , �  /� �  0� o  0� o  /� �  /�      F  , , C  /� C  0�   0�   /� C  /�      F  , , �  /� �  0�  �  0�  �  /� �  /�      F  , , ${  /� ${  0� %C  0� %C  /� ${  /�      F  , , )  /� )  0� )�  0� )�  /� )  /�      F  , , -�  /� -�  0� .{  0� .{  /� -�  /�      F  , , )  .6 )  .� )�  .� )�  .6 )  .6      F  , , �  "� �  #Z o  #Z o  "� �  "�      F  , , C  "� C  #Z   #Z   "� C  "�      F  , , �  "� �  #Z  �  #Z  �  "� �  "�      F  , , �  2� �  3� o  3� o  2� �  2�      F  , , C  2� C  3�   3�   2� C  2�      F  , , �  2� �  3�  �  3�  �  2� �  2�      F  , , ${  2� ${  3� %C  3� %C  2� ${  2�      F  , , )  2� )  3� )�  3� )�  2� )  2�      F  , , -�  2� -�  3� .{  3� .{  2� -�  2�      F  , , -�  .6 -�  .� .{  .� .{  .6 -�  .6      F  , , �  r �   :  �   :  �  r �  r      F  , , ${  r ${   : %C   : %C  r ${  r      F  , , )  r )   : )�   : )�  r )  r      F  , , -�  r -�   : .{   : .{  r -�  r      F  , , )  ,� )  -n )�  -n )�  ,� )  ,�      F  , , �  )� �  *N o  *N o  )� �  )�      F  , , C  )� C  *N   *N   )� C  )�      F  , , �  )� �  *N  �  *N  �  )� �  )�      F  , , ${  )� ${  *N %C  *N %C  )� ${  )�      F  , , )  )� )  *N )�  *N )�  )� )  )�      F  , , ${  "� ${  #Z %C  #Z %C  "� ${  "�      F  , , )  "� )  #Z )�  #Z )�  "� )  "�      F  , , -�  "� -�  #Z .{  #Z .{  "� -�  "�      F  , ,  �c  �  �c  �  �+  �  �+  �  �c  �      F  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      F  , ,  ��  �  ��  �  c  �  c  �  ��  �      F  , , 7  � 7  � �  � �  � 7  �      F  , , �  � �  � 	�  � 	�  � �  �      F  , , o  � o  � 7  � 7  � o  �      F  , ,   �   � �  � �  �   �      F  , ,  ��  !  ��  !�  c  !�  c  !  ��  !      F  , , 7  ! 7  !� �  !� �  ! 7  !      F  , , �  ! �  !� 	�  !� 	�  ! �  !      F  , , o  ! o  !� 7  !� 7  ! o  !      F  , ,   !   !� �  !� �  !   !      F  , , 7  /� 7  0� �  0� �  /� 7  /�      F  , ,  �c  �  �c  �  �+  �  �+  �  �c  �      F  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      F  , ,  ��  �  ��  �  c  �  c  �  ��  �      F  , , 7  � 7  � �  � �  � 7  �      F  , , �  � �  � 	�  � 	�  � �  �      F  , , o  � o  � 7  � 7  � o  �      F  , ,   �   � �  � �  �   �      F  , , �  /� �  0� 	�  0� 	�  /� �  /�      F  , , o  /� o  0� 7  0� 7  /� o  /�      F  , ,   /�   0� �  0� �  /�   /�      F  , ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      F  , ,  ��  2�  ��  3�  c  3�  c  2�  ��  2�      F  , , 7  2� 7  3� �  3� �  2� 7  2�      F  , ,  �c  1V  �c  2  �+  2  �+  1V  �c  1V      F  , ,  ��  1V  ��  2  ��  2  ��  1V  ��  1V      F  , ,  ��  1V  ��  2  c  2  c  1V  ��  1V      F  , , 7  1V 7  2 �  2 �  1V 7  1V      F  , , �  1V �  2 	�  2 	�  1V �  1V      F  , , o  1V o  2 7  2 7  1V o  1V      F  , ,   1V   2 �  2 �  1V   1V      F  , , �  2� �  3� 	�  3� 	�  2� �  2�      F  , ,  �c  .6  �c  .�  �+  .�  �+  .6  �c  .6      F  , ,  ��  .6  ��  .�  ��  .�  ��  .6  ��  .6      F  , ,  �c  "�  �c  #Z  �+  #Z  �+  "�  �c  "�      F  , ,  ��  "�  ��  #Z  ��  #Z  ��  "�  ��  "�      F  , ,  ��  "�  ��  #Z  c  #Z  c  "�  ��  "�      F  , ,  �c  2  �c  �  �+  �  �+  2  �c  2      F  , ,  ��  2  ��  �  ��  �  ��  2  ��  2      F  , ,  ��  2  ��  �  c  �  c  2  ��  2      F  , , 7  2 7  � �  � �  2 7  2      F  , , �  2 �  � 	�  � 	�  2 �  2      F  , , o  2 o  � 7  � 7  2 o  2      F  , ,   2   � �  � �  2   2      F  , , 7  "� 7  #Z �  #Z �  "� 7  "�      F  , , �  "� �  #Z 	�  #Z 	�  "� �  "�      F  , , o  "� o  #Z 7  #Z 7  "� o  "�      F  , ,   "�   #Z �  #Z �  "�   "�      F  , ,  ��  .6  ��  .�  c  .�  c  .6  ��  .6      F  , , 7  .6 7  .� �  .� �  .6 7  .6      F  , , �  .6 �  .� 	�  .� 	�  .6 �  .6      F  , , o  .6 o  .� 7  .� 7  .6 o  .6      F  , ,   .6   .� �  .� �  .6   .6      F  , , o  2� o  3� 7  3� 7  2� o  2�      F  , ,   2�   3� �  3� �  2�   2�      F  , ,  �c  2�  �c  3�  �+  3�  �+  2�  �c  2�      F  , ,  �c  r  �c   :  �+   :  �+  r  �c  r      F  , ,  �c  R  �c    �+    �+  R  �c  R      F  , ,  ��  R  ��    ��    ��  R  ��  R      F  , ,  ��  R  ��    c    c  R  ��  R      F  , , 7  R 7   �   �  R 7  R      F  , , �  R �   	�   	�  R �  R      F  , , o  R o   7   7  R o  R      F  , ,   R    �   �  R   R      F  , ,  ��  r  ��   :  ��   :  ��  r  ��  r      F  , ,  ��  r  ��   :  c   :  c  r  ��  r      F  , , 7  r 7   : �   : �  r 7  r      F  , , �  r �   : 	�   : 	�  r �  r      F  , , o  r o   : 7   : 7  r o  r      F  , ,   r    : �   : �  r   r      F  , ,  �c  /�  �c  0�  �+  0�  �+  /�  �c  /�      F  , ,  �c  ,�  �c  -n  �+  -n  �+  ,�  �c  ,�      F  , ,  �c  )�  �c  *N  �+  *N  �+  )�  �c  )�      F  , ,  ��  )�  ��  *N  ��  *N  ��  )�  ��  )�      F  , ,  ��  )�  ��  *N  c  *N  c  )�  ��  )�      F  , , 7  )� 7  *N �  *N �  )� 7  )�      F  , , �  )� �  *N 	�  *N 	�  )� �  )�      F  , , o  )� o  *N 7  *N 7  )� o  )�      F  , ,   )�   *N �  *N �  )�   )�      F  , ,  ��  ,�  ��  -n  ��  -n  ��  ,�  ��  ,�      F  , ,  ��  ,�  ��  -n  c  -n  c  ,�  ��  ,�      F  , , 7  ,� 7  -n �  -n �  ,� 7  ,�      F  , ,  �c  +  �c  +�  �+  +�  �+  +  �c  +      F  , ,  ��  +  ��  +�  ��  +�  ��  +  ��  +      F  , ,  ��  +  ��  +�  c  +�  c  +  ��  +      F  , , 7  + 7  +� �  +� �  + 7  +      F  , , �  + �  +� 	�  +� 	�  + �  +      F  , , o  + o  +� 7  +� 7  + o  +      F  , ,   +   +� �  +� �  +   +      F  , , �  ,� �  -n 	�  -n 	�  ,� �  ,�      F  , , o  ,� o  -n 7  -n 7  ,� o  ,�      F  , ,   ,�   -n �  -n �  ,�   ,�      F  , ,  ��  /�  ��  0�  ��  0�  ��  /�  ��  /�      F  , ,  ��  /�  ��  0�  c  0�  c  /�  ��  /�      F  , ,  �c  !  �c  !�  �+  !�  �+  !  �c  !      F  , ,  ��  !  ��  !�  ��  !�  ��  !  ��  !      F  , ,  `'  �  `'  V  `�  V  `�  �  `'  �      F  , ,  d�  �  d�  V  e�  V  e�  �  d�  �      F  , ,  i_  �  i_  V  j'  V  j'  �  i_  �      F  , ,  m�  �  m�  V  n�  V  n�  �  m�  �      F  , ,  r�  �  r�  V  s_  V  s_  �  r�  �      F  , ,  w3  �  w3  V  w�  V  w�  �  w3  �      F  , ,  {�  �  {�  V  |�  V  |�  �  {�  �      F  , ,  `'  �  `'  �  `�  �  `�  �  `'  �      F  , ,  d�  �  d�  �  e�  �  e�  �  d�  �      F  , ,  i_  �  i_  �  j'  �  j'  �  i_  �      F  , ,  m�  �  m�  �  n�  �  n�  �  m�  �      F  , ,  r�  �  r�  �  s_  �  s_  �  r�  �      F  , ,  w3  �  w3  �  w�  �  w�  �  w3  �      F  , ,  {�  �  {�  �  |�  �  |�  �  {�  �      F  , ,  `'  n  `'  6  `�  6  `�  n  `'  n      F  , ,  d�  n  d�  6  e�  6  e�  n  d�  n      F  , ,  i_  n  i_  6  j'  6  j'  n  i_  n      F  , ,  m�  n  m�  6  n�  6  n�  n  m�  n      F  , ,  r�  n  r�  6  s_  6  s_  n  r�  n      F  , ,  w3  n  w3  6  w�  6  w�  n  w3  n      F  , ,  {�  n  {�  6  |�  6  |�  n  {�  n      F  , ,  `'  �  `'  �  `�  �  `�  �  `'  �      F  , ,  d�  �  d�  �  e�  �  e�  �  d�  �      F  , ,  i_  �  i_  �  j'  �  j'  �  i_  �      F  , ,  m�  �  m�  �  n�  �  n�  �  m�  �      F  , ,  r�  �  r�  �  s_  �  s_  �  r�  �      F  , ,  w3  �  w3  �  w�  �  w�  �  w3  �      F  , ,  {�  �  {�  �  |�  �  |�  �  {�  �      F  , ,  `'  N  `'    `�    `�  N  `'  N      F  , ,  d�  N  d�    e�    e�  N  d�  N      F  , ,  i_  N  i_    j'    j'  N  i_  N      F  , ,  m�  N  m�    n�    n�  N  m�  N      F  , ,  r�  N  r�    s_    s_  N  r�  N      F  , ,  w3  N  w3    w�    w�  N  w3  N      F  , ,  {�  N  {�    |�    |�  N  {�  N      F  , ,  `'  Z  `'  "  `�  "  `�  Z  `'  Z      F  , ,  d�  Z  d�  "  e�  "  e�  Z  d�  Z      F  , ,  i_  Z  i_  "  j'  "  j'  Z  i_  Z      F  , ,  m�  Z  m�  "  n�  "  n�  Z  m�  Z      F  , ,  r�  Z  r�  "  s_  "  s_  Z  r�  Z      F  , ,  w3  Z  w3  "  w�  "  w�  Z  w3  Z      F  , ,  {�  Z  {�  "  |�  "  |�  Z  {�  Z      F  , ,  `'  �  `'  �  `�  �  `�  �  `'  �      F  , ,  d�  �  d�  �  e�  �  e�  �  d�  �      F  , ,  i_  �  i_  �  j'  �  j'  �  i_  �      F  , ,  m�  �  m�  �  n�  �  n�  �  m�  �      F  , ,  r�  �  r�  �  s_  �  s_  �  r�  �      F  , ,  w3  �  w3  �  w�  �  w�  �  w3  �      F  , ,  {�  �  {�  �  |�  �  |�  �  {�  �      F  , ,  `'  :  `'    `�    `�  :  `'  :      F  , ,  d�  :  d�    e�    e�  :  d�  :      F  , ,  i_  :  i_    j'    j'  :  i_  :      F  , ,  m�  :  m�    n�    n�  :  m�  :      F  , ,  r�  :  r�    s_    s_  :  r�  :      F  , ,  w3  :  w3    w�    w�  :  w3  :      F  , ,  {�  :  {�    |�    |�  :  {�  :      F  , ,  `'   �  `'  r  `�  r  `�   �  `'   �      F  , ,  d�   �  d�  r  e�  r  e�   �  d�   �      F  , ,  i_   �  i_  r  j'  r  j'   �  i_   �      F  , ,  m�   �  m�  r  n�  r  n�   �  m�   �      F  , ,  r�   �  r�  r  s_  r  s_   �  r�   �      F  , ,  w3   �  w3  r  w�  r  w�   �  w3   �      F  , ,  {�   �  {�  r  |�  r  |�   �  {�   �      F  , ,  `'���  `'����  `�����  `����  `'���      F  , ,  d����  d�����  e�����  e����  d����      F  , ,  i_���  i_����  j'����  j'���  i_���      F  , ,  m����  m�����  n�����  n����  m����      F  , ,  r����  r�����  s_����  s_���  r����      F  , ,  w3���  w3����  w�����  w����  w3���      F  , ,  {����  {�����  |�����  |����  {����      F  , ,  `'����  `'���R  `����R  `�����  `'����      F  , ,  d�����  d����R  e����R  e�����  d�����      F  , ,  i_����  i_���R  j'���R  j'����  i_����      F  , ,  m�����  m����R  n����R  n�����  m�����      F  , ,  r�����  r����R  s_���R  s_����  r�����      F  , ,  w3����  w3���R  w����R  w�����  w3����      F  , ,  {�����  {����R  |����R  |�����  {�����      F  , ,  `'����  `'����  `�����  `�����  `'����      F  , ,  d�����  d�����  e�����  e�����  d�����      F  , ,  i_����  i_����  j'����  j'����  i_����      F  , ,  m�����  m�����  n�����  n�����  m�����      F  , ,  r�����  r�����  s_����  s_����  r�����      F  , ,  w3����  w3����  w�����  w�����  w3����      F  , ,  {�����  {�����  |�����  |�����  {�����      F  , ,  `'  �  `'  v  `�  v  `�  �  `'  �      F  , ,  d�  �  d�  v  e�  v  e�  �  d�  �      F  , ,  i_  �  i_  v  j'  v  j'  �  i_  �      F  , ,  m�  �  m�  v  n�  v  n�  �  m�  �      F  , ,  r�  �  r�  v  s_  v  s_  �  r�  �      F  , ,  w3  �  w3  v  w�  v  w�  �  w3  �      F  , ,  {�  �  {�  v  |�  v  |�  �  {�  �      F  , ,  `'    `'  �  `�  �  `�    `'        F  , ,  d�    d�  �  e�  �  e�    d�        F  , ,  i_    i_  �  j'  �  j'    i_        F  , ,  m�    m�  �  n�  �  n�    m�        F  , ,  r�    r�  �  s_  �  s_    r�        F  , ,  w3    w3  �  w�  �  w�    w3        F  , ,  {�    {�  �  |�  �  |�    {�        F  , ,  �?  :  �?    �    �  :  �?  :      F  , ,  ��  :  ��    ��    ��  :  ��  :      F  , ,  ��    ��  �  �k  �  �k    ��        F  , ,  �?    �?  �  �  �  �    �?        F  , ,  �k  �  �k  V  �3  V  �3  �  �k  �      F  , ,  �k  N  �k    �3    �3  N  �k  N      F  , ,  �  N  �    ��    ��  N  �  N      F  , ,  ��  N  ��    �k    �k  N  ��  N      F  , ,  �?  N  �?    �    �  N  �?  N      F  , ,  �k   �  �k  r  �3  r  �3   �  �k   �      F  , ,  �   �  �  r  ��  r  ��   �  �   �      F  , ,  ��   �  ��  r  �k  r  �k   �  ��   �      F  , ,  �?   �  �?  r  �  r  �   �  �?   �      F  , ,  ��   �  ��  r  ��  r  ��   �  ��   �      F  , ,  ��  N  ��    ��    ��  N  ��  N      F  , ,  �k  n  �k  6  �3  6  �3  n  �k  n      F  , ,  �  n  �  6  ��  6  ��  n  �  n      F  , ,  ��  n  ��  6  �k  6  �k  n  ��  n      F  , ,  �?  n  �?  6  �  6  �  n  �?  n      F  , ,  ��  n  ��  6  ��  6  ��  n  ��  n      F  , ,  �  �  �  V  ��  V  ��  �  �  �      F  , ,  �k���  �k����  �3����  �3���  �k���      F  , ,  ����  �����  ������  �����  ����      F  , ,  �����  ������  �k����  �k���  �����      F  , ,  �?���  �?����  �����  ����  �?���      F  , ,  �����  ������  ������  �����  �����      F  , ,  ��  �  ��  V  �k  V  �k  �  ��  �      F  , ,  �k  Z  �k  "  �3  "  �3  Z  �k  Z      F  , ,  �  Z  �  "  ��  "  ��  Z  �  Z      F  , ,  ��  Z  ��  "  �k  "  �k  Z  ��  Z      F  , ,  �?  Z  �?  "  �  "  �  Z  �?  Z      F  , ,  ��  Z  ��  "  ��  "  ��  Z  ��  Z      F  , ,  �k  �  �k  �  �3  �  �3  �  �k  �      F  , ,  �k����  �k���R  �3���R  �3����  �k����      F  , ,  �����  ����R  �����R  ������  �����      F  , ,  ������  �����R  �k���R  �k����  ������      F  , ,  �?����  �?���R  ����R  �����  �?����      F  , ,  ������  �����R  �����R  ������  ������      F  , ,  �  �  �  �  ��  �  ��  �  �  �      F  , ,  ��  �  ��  �  �k  �  �k  �  ��  �      F  , ,  �?  �  �?  �  �  �  �  �  �?  �      F  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      F  , ,  �k  �  �k  �  �3  �  �3  �  �k  �      F  , ,  �  �  �  �  ��  �  ��  �  �  �      F  , ,  �k  �  �k  �  �3  �  �3  �  �k  �      F  , ,  �k����  �k����  �3����  �3����  �k����      F  , ,  �����  �����  ������  ������  �����      F  , ,  ������  ������  �k����  �k����  ������      F  , ,  �?����  �?����  �����  �����  �?����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �  �  �  �  ��  �  ��  �  �  �      F  , ,  ��  �  ��  �  �k  �  �k  �  ��  �      F  , ,  �?  �  �?  �  �  �  �  �  �?  �      F  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      F  , ,  ��  �  ��  �  �k  �  �k  �  ��  �      F  , ,  �?  �  �?  �  �  �  �  �  �?  �      F  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      F  , ,  �k  �  �k  v  �3  v  �3  �  �k  �      F  , ,  �  �  �  v  ��  v  ��  �  �  �      F  , ,  ��  �  ��  v  �k  v  �k  �  ��  �      F  , ,  �?  �  �?  v  �  v  �  �  �?  �      F  , ,  ��  �  ��  v  ��  v  ��  �  ��  �      F  , ,  �?  �  �?  V  �  V  �  �  �?  �      F  , ,  ��  �  ��  V  ��  V  ��  �  ��  �      F  , ,  ��    ��  �  ��  �  ��    ��        F  , ,  �    �  �  ��  �  ��    �        F  , ,  �k  :  �k    �3    �3  :  �k  :      F  , ,  �  :  �    ��    ��  :  �  :      F  , ,  ��  :  ��    �k    �k  :  ��  :      F  , ,  �k    �k  �  �3  �  �3    �k        F  , ,  ����  �����  ������  �����  ����      F  , ,  �����  ������  �k����  �k���  �����      F  , ,  �?���  �?����  �����  ����  �?���      F  , ,  �����  ������  ������  �����  �����      F  , ,  �k���  �k���L  �3���L  �3���  �k���      F  , ,  ����  ����L  �����L  �����  ����      F  , ,  �����  �����L  �k���L  �k���  �����      F  , ,  �?���  �?���L  ����L  ����  �?���      F  , ,  �����  �����L  �����L  �����  �����      F  , ,  �k����  �k���  �3���  �3����  �k����      F  , ,  �����  ����  �����  ������  �����      F  , ,  ������  �����  �k���  �k����  ������      F  , ,  �?����  �?���  ����  �����  �?����      F  , ,  ������  �����  �����  ������  ������      F  , ,  �k���d  �k���,  �3���,  �3���d  �k���d      F  , ,  ����d  ����,  �����,  �����d  ����d      F  , ,  �����d  �����,  �k���,  �k���d  �����d      F  , ,  �?���d  �?���,  ����,  ����d  �?���d      F  , ,  �����d  �����,  �����,  �����d  �����d      F  , ,  �k����  �k���  �3���  �3����  �k����      F  , ,  �����  ����  �����  ������  �����      F  , ,  ������  �����  �k���  �k����  ������      F  , ,  �?����  �?���  ����  �����  �?����      F  , ,  ������  �����  �����  ������  ������      F  , ,  �k���D  �k���  �3���  �3���D  �k���D      F  , ,  ����D  ����  �����  �����D  ����D      F  , ,  �����D  �����  �k���  �k���D  �����D      F  , ,  �?���D  �?���  ����  ����D  �?���D      F  , ,  �����D  �����  �����  �����D  �����D      F  , ,  �k���P  �k���  �3���  �3���P  �k���P      F  , ,  ����P  ����  �����  �����P  ����P      F  , ,  �����P  �����  �k���  �k���P  �����P      F  , ,  �?���P  �?���  ����  ����P  �?���P      F  , ,  �����P  �����  �����  �����P  �����P      F  , ,  �k���  �k���l  �3���l  �3���  �k���      F  , ,  ����  ����l  �����l  �����  ����      F  , ,  �����  �����l  �k���l  �k���  �����      F  , ,  �?���  �?���l  ����l  ����  �?���      F  , ,  �����  �����l  �����l  �����  �����      F  , ,  �k���  �k����  �3����  �3���  �k���      F  , ,  `'����  `'���  `����  `�����  `'����      F  , ,  d�����  d����  e����  e�����  d�����      F  , ,  i_����  i_���  j'���  j'����  i_����      F  , ,  m�����  m����  n����  n�����  m�����      F  , ,  r�����  r����  s_���  s_����  r�����      F  , ,  w3����  w3���  w����  w�����  w3����      F  , ,  {�����  {����  |����  |�����  {�����      F  , ,  m�����  m����  n����  n�����  m�����      F  , ,  r�����  r����  s_���  s_����  r�����      F  , ,  w3����  w3���  w����  w�����  w3����      F  , ,  {�����  {����  |����  |�����  {�����      F  , ,  w3���  w3���L  w����L  w����  w3���      F  , ,  `'���D  `'���  `����  `����D  `'���D      F  , ,  d����D  d����  e����  e����D  d����D      F  , ,  i_���D  i_���  j'���  j'���D  i_���D      F  , ,  m����D  m����  n����  n����D  m����D      F  , ,  r����D  r����  s_���  s_���D  r����D      F  , ,  w3���D  w3���  w����  w����D  w3���D      F  , ,  {����D  {����  |����  |����D  {����D      F  , ,  {����  {����L  |����L  |����  {����      F  , ,  `'���  `'���L  `����L  `����  `'���      F  , ,  d����  d����L  e����L  e����  d����      F  , ,  i_���  i_���L  j'���L  j'���  i_���      F  , ,  `'���d  `'���,  `����,  `����d  `'���d      F  , ,  `'���P  `'���  `����  `����P  `'���P      F  , ,  d����P  d����  e����  e����P  d����P      F  , ,  i_���P  i_���  j'���  j'���P  i_���P      F  , ,  m����P  m����  n����  n����P  m����P      F  , ,  r����P  r����  s_���  s_���P  r����P      F  , ,  w3���P  w3���  w����  w����P  w3���P      F  , ,  {����P  {����  |����  |����P  {����P      F  , ,  d����d  d����,  e����,  e����d  d����d      F  , ,  i_���d  i_���,  j'���,  j'���d  i_���d      F  , ,  m����d  m����,  n����,  n����d  m����d      F  , ,  r����d  r����,  s_���,  s_���d  r����d      F  , ,  w3���d  w3���,  w����,  w����d  w3���d      F  , ,  `'���  `'���l  `����l  `����  `'���      F  , ,  d����  d����l  e����l  e����  d����      F  , ,  i_���  i_���l  j'���l  j'���  i_���      F  , ,  m����  m����l  n����l  n����  m����      F  , ,  r����  r����l  s_���l  s_���  r����      F  , ,  w3���  w3���l  w����l  w����  w3���      F  , ,  {����  {����l  |����l  |����  {����      F  , ,  {����d  {����,  |����,  |����d  {����d      F  , ,  m����  m����L  n����L  n����  m����      F  , ,  r����  r����L  s_���L  s_���  r����      F  , ,  `'����  `'���  `����  `�����  `'����      F  , ,  d�����  d����  e����  e�����  d�����      F  , ,  `'���  `'����  `�����  `����  `'���      F  , ,  d����  d�����  e�����  e����  d����      F  , ,  i_���  i_����  j'����  j'���  i_���      F  , ,  m����  m�����  n�����  n����  m����      F  , ,  r����  r�����  s_����  s_���  r����      F  , ,  w3���  w3����  w�����  w����  w3���      F  , ,  {����  {�����  |�����  |����  {����      F  , ,  i_����  i_���  j'���  j'����  i_����      F  , ,  {���ؠ  {����h  |����h  |���ؠ  {���ؠ      F  , ,  `'���  `'����  `�����  `����  `'���      F  , ,  d����  d�����  e�����  e����  d����      F  , ,  i_���  i_����  j'����  j'���  i_���      F  , ,  m����  m�����  n�����  n����  m����      F  , ,  r����  r�����  s_����  s_���  r����      F  , ,  w3���  w3����  w�����  w����  w3���      F  , ,  {����  {�����  |�����  |����  {����      F  , ,  `'��Հ  `'���H  `����H  `���Հ  `'��Հ      F  , ,  d���Հ  d����H  e����H  e���Հ  d���Հ      F  , ,  i_��Հ  i_���H  j'���H  j'��Հ  i_��Հ      F  , ,  m���Հ  m����H  n����H  n���Հ  m���Հ      F  , ,  r���Հ  r����H  s_���H  s_��Հ  r���Հ      F  , ,  w3��Հ  w3���H  w����H  w���Հ  w3��Հ      F  , ,  {���Հ  {����H  |����H  |���Հ  {���Հ      F  , ,  `'����  `'��Ը  `���Ը  `�����  `'����      F  , ,  d�����  d���Ը  e���Ը  e�����  d�����      F  , ,  i_����  i_��Ը  j'��Ը  j'����  i_����      F  , ,  m�����  m���Ը  n���Ը  n�����  m�����      F  , ,  r�����  r���Ը  s_��Ը  s_����  r�����      F  , ,  w3����  w3��Ը  w���Ը  w�����  w3����      F  , ,  {�����  {���Ը  |���Ը  |�����  {�����      F  , ,  `'����  `'��܈  `���܈  `�����  `'����      F  , ,  d�����  d���܈  e���܈  e�����  d�����      F  , ,  i_����  i_��܈  j'��܈  j'����  i_����      F  , ,  m�����  m���܈  n���܈  n�����  m�����      F  , ,  r�����  r���܈  s_��܈  s_����  r�����      F  , ,  w3����  w3��܈  w���܈  w�����  w3����      F  , ,  {�����  {���܈  |���܈  |�����  {�����      F  , ,  `'���0  `'����  `�����  `����0  `'���0      F  , ,  d����0  d�����  e�����  e����0  d����0      F  , ,  i_���0  i_����  j'����  j'���0  i_���0      F  , ,  m����0  m�����  n�����  n����0  m����0      F  , ,  r����0  r�����  s_����  s_���0  r����0      F  , ,  w3���0  w3����  w�����  w����0  w3���0      F  , ,  {����0  {�����  |�����  |����0  {����0      F  , ,  `'��ؠ  `'���h  `����h  `���ؠ  `'��ؠ      F  , ,  d���ؠ  d����h  e����h  e���ؠ  d���ؠ      F  , ,  i_��ؠ  i_���h  j'���h  j'��ؠ  i_��ؠ      F  , ,  m���ؠ  m����h  n����h  n���ؠ  m���ؠ      F  , ,  r���ؠ  r����h  s_���h  s_��ؠ  r���ؠ      F  , ,  w3��ؠ  w3���h  w����h  w���ؠ  w3��ؠ      F  , ,  �?���0  �?����  �����  ����0  �?���0      F  , ,  �����0  ������  ������  �����0  �����0      F  , ,  ������  ����܈  �k��܈  �k����  ������      F  , ,  �?����  �?��܈  ���܈  �����  �?����      F  , ,  ������  ����܈  ����܈  ������  ������      F  , ,  �k����  �k��Ը  �3��Ը  �3����  �k����      F  , ,  �����  ���Ը  ����Ը  ������  �����      F  , ,  ������  ����Ը  �k��Ը  �k����  ������      F  , ,  �?����  �?��Ը  ���Ը  �����  �?����      F  , ,  ������  ����Ը  ����Ը  ������  ������      F  , ,  �'��Ś  �'���b  �����b  ����Ś  �'��Ś      F  , ,  ����Ś  �����b  �����b  ����Ś  ����Ś      F  , ,  �_��Ś  �_���b  �'���b  �'��Ś  �_��Ś      F  , ,  ����Ś  �����b  �����b  ����Ś  ����Ś      F  , ,  ����Ś  �����b  �_���b  �_��Ś  ����Ś      F  , ,  �'���
  �'����  ������  �����
  �'���
      F  , ,  �����
  ������  ������  �����
  �����
      F  , ,  �_���
  �_����  �'����  �'���
  �_���
      F  , ,  �����
  ������  ������  �����
  �����
      F  , ,  �����
  ������  �_����  �_���
  �����
      F  , ,  �'���z  �'���B  �����B  �����z  �'���z      F  , ,  �����z  �����B  �����B  �����z  �����z      F  , ,  �_���z  �_���B  �'���B  �'���z  �_���z      F  , ,  �����z  �����B  �����B  �����z  �����z      F  , ,  �����z  �����B  �_���B  �_���z  �����z      F  , ,  �'����  �'����  ������  ������  �'����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �_����  �_����  �'����  �'����  �_����      F  , ,  ������  ������  ������  ������  ������      F  , ,  ������  ������  �_����  �_����  ������      F  , ,  �k����  �k��܈  �3��܈  �3����  �k����      F  , ,  �k���  �k����  �3����  �3���  �k���      F  , ,  ����  �����  ������  �����  ����      F  , ,  �����  ������  �k����  �k���  �����      F  , ,  �?���  �?����  �����  ����  �?���      F  , ,  �����  ������  ������  �����  �����      F  , ,  �����  ���܈  ����܈  ������  �����      F  , ,  �k���0  �k����  �3����  �3���0  �k���0      F  , ,  ����0  �����  ������  �����0  ����0      F  , ,  �k��ؠ  �k���h  �3���h  �3��ؠ  �k��ؠ      F  , ,  ���ؠ  ����h  �����h  ����ؠ  ���ؠ      F  , ,  ����ؠ  �����h  �k���h  �k��ؠ  ����ؠ      F  , ,  �?��ؠ  �?���h  ����h  ���ؠ  �?��ؠ      F  , ,  �k��Հ  �k���H  �3���H  �3��Հ  �k��Հ      F  , ,  ���Հ  ����H  �����H  ����Հ  ���Հ      F  , ,  ����Հ  �����H  �k���H  �k��Հ  ����Հ      F  , ,  �?��Հ  �?���H  ����H  ���Հ  �?��Հ      F  , ,  ����Հ  �����H  �����H  ����Հ  ����Հ      F  , ,  ����ؠ  �����h  �����h  ����ؠ  ����ؠ      F  , ,  �����0  ������  �k����  �k���0  �����0      F  , ,  �k���
  �k����  �3����  �3���
  �k���
      F  , ,  �3����  �3����  ������  ������  �3����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �k����  �k����  �3����  �3����  �k����      F  , ,  �����  �����  ������  ������  �����      F  , ,  ţ����  ţ����  �k����  �k����  ţ����      F  , ,  �?����  �?����  �����  �����  �?����      F  , ,  ������  ������  ϣ����  ϣ����  ������      F  , ,  ����
  �����  ������  �����
  ����
      F  , ,  ţ���
  ţ����  �k����  �k���
  ţ���
      F  , ,  �?���
  �?����  �����  ����
  �?���
      F  , ,  �����
  ������  ϣ����  ϣ���
  �����
      F  , ,  �?��Ś  �?���b  ����b  ���Ś  �?��Ś      F  , ,  ����Ś  �����b  ϣ���b  ϣ��Ś  ����Ś      F  , ,  �3��Ś  �3���b  �����b  ����Ś  �3��Ś      F  , ,  ����Ś  �����b  �����b  ����Ś  ����Ś      F  , ,  �k��Ś  �k���b  �3���b  �3��Ś  �k��Ś      F  , ,  �3���z  �3���B  �����B  �����z  �3���z      F  , ,  �����z  �����B  �����B  �����z  �����z      F  , ,  �k���z  �k���B  �3���B  �3���z  �k���z      F  , ,  ����z  ����B  �����B  �����z  ����z      F  , ,  ţ���z  ţ���B  �k���B  �k���z  ţ���z      F  , ,  �?���z  �?���B  ����B  ����z  �?���z      F  , ,  �����z  �����B  ϣ���B  ϣ���z  �����z      F  , ,  ���Ś  ����b  �����b  ����Ś  ���Ś      F  , ,  ţ��Ś  ţ���b  �k���b  �k��Ś  ţ��Ś      F  , ,  �3���
  �3����  ������  �����
  �3���
      F  , ,  �����
  ������  ������  �����
  �����
      F  , ,  �����  �����  ������  ������  �����      F  , ,  ţ����  ţ����  �k����  �k����  ţ����      F  , ,  �?����  �?����  �����  �����  �?����      F  , ,  ������  ������  ϣ����  ϣ����  ������      F  , ,  �3���:  �3���  �����  �����:  �3���:      F  , ,  �����:  �����  �����  �����:  �����:      F  , ,  �k���:  �k���  �3���  �3���:  �k���:      F  , ,  ����:  ����  �����  �����:  ����:      F  , ,  ţ���:  ţ���  �k���  �k���:  ţ���:      F  , ,  �?���:  �?���  ����  ����:  �?���:      F  , ,  �����:  �����  ϣ���  ϣ���:  �����:      F  , ,  �3���F  �3���  �����  �����F  �3���F      F  , ,  �����F  �����  �����  �����F  �����F      F  , ,  �k���F  �k���  �3���  �3���F  �k���F      F  , ,  ����F  ����  �����  �����F  ����F      F  , ,  ţ���F  ţ���  �k���  �k���F  ţ���F      F  , ,  �?���F  �?���  ����  ����F  �?���F      F  , ,  �����F  �����  ϣ���  ϣ���F  �����F      F  , ,  �3����  �3���~  �����~  ������  �3����      F  , ,  ������  �����~  �����~  ������  ������      F  , ,  �k����  �k���~  �3���~  �3����  �k����      F  , ,  �����  ����~  �����~  ������  �����      F  , ,  ţ����  ţ���~  �k���~  �k����  ţ����      F  , ,  �?����  �?���~  ����~  �����  �?����      F  , ,  ������  �����~  ϣ���~  ϣ����  ������      F  , ,  �3���&  �3����  ������  �����&  �3���&      F  , ,  �����&  ������  ������  �����&  �����&      F  , ,  �k���&  �k����  �3����  �3���&  �k���&      F  , ,  ����&  �����  ������  �����&  ����&      F  , ,  ţ���&  ţ����  �k����  �k���&  ţ���&      F  , ,  �?���&  �?����  �����  ����&  �?���&      F  , ,  �����&  ������  ϣ����  ϣ���&  �����&      F  , ,  �3����  �3���^  �����^  ������  �3����      F  , ,  ������  �����^  �����^  ������  ������      F  , ,  �k����  �k���^  �3���^  �3����  �k����      F  , ,  �����  ����^  �����^  ������  �����      F  , ,  ţ����  ţ���^  �k���^  �k����  ţ����      F  , ,  �?����  �?���^  ����^  �����  �?����      F  , ,  ������  �����^  ϣ���^  ϣ����  ������      F  , ,  �3���  �3����  ������  �����  �3���      F  , ,  �����  ������  ������  �����  �����      F  , ,  �k���  �k����  �3����  �3���  �k���      F  , ,  ����  �����  ������  �����  ����      F  , ,  ţ���  ţ����  �k����  �k���  ţ���      F  , ,  �?���  �?����  �����  ����  �?���      F  , ,  �����  ������  ϣ����  ϣ���  �����      F  , ,  �3���v  �3���>  �����>  �����v  �3���v      F  , ,  �����v  �����>  �����>  �����v  �����v      F  , ,  �k���v  �k���>  �3���>  �3���v  �k���v      F  , ,  ����v  ����>  �����>  �����v  ����v      F  , ,  ţ���v  ţ���>  �k���>  �k���v  ţ���v      F  , ,  �?���v  �?���>  ����>  ����v  �?���v      F  , ,  �����v  �����>  ϣ���>  ϣ���v  �����v      F  , ,  �3����  �3����  ������  ������  �3����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �k����  �k����  �3����  �3����  �k����      F  , ,  �����  �����  ������  ������  �����      F  , ,  ţ����  ţ����  �k����  �k����  ţ����      F  , ,  �?����  �?����  �����  �����  �?����      F  , ,  ������  ������  ϣ����  ϣ����  ������      F  , ,  �3���Z  �3���"  �����"  �����Z  �3���Z      F  , ,  �����Z  �����"  �����"  �����Z  �����Z      F  , ,  �k���Z  �k���"  �3���"  �3���Z  �k���Z      F  , ,  ����Z  ����"  �����"  �����Z  ����Z      F  , ,  ţ���Z  ţ���"  �k���"  �k���Z  ţ���Z      F  , ,  �?���Z  �?���"  ����"  ����Z  �?���Z      F  , ,  �����Z  �����"  ϣ���"  ϣ���Z  �����Z      F  , ,  �3����  �3����  ������  ������  �3����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �k����  �k����  �3����  �3����  �k����      F  , ,  ����   �����  ������  �����   ����       F  , ,  ţ���   ţ����  �k����  �k���   ţ���       F  , ,  �?���   �?����  �����  ����   �?���       F  , ,  �����   ������  ϣ����  ϣ���   �����       F  , ,  �3���p  �3���8  �����8  �����p  �3���p      F  , ,  �����p  �����8  �����8  �����p  �����p      F  , ,  �k���p  �k���8  �3���8  �3���p  �k���p      F  , ,  ����p  ����8  �����8  �����p  ����p      F  , ,  ţ���p  ţ���8  �k���8  �k���p  ţ���p      F  , ,  �?���p  �?���8  ����8  ����p  �?���p      F  , ,  �����p  �����8  ϣ���8  ϣ���p  �����p      F  , ,  �3����  �3����  ������  ������  �3����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �k����  �k����  �3����  �3����  �k����      F  , ,  �����  �����  ������  ������  �����      F  , ,  ţ����  ţ����  �k����  �k����  ţ����      F  , ,  �?����  �?����  �����  �����  �?����      F  , ,  ������  ������  ϣ����  ϣ����  ������      F  , ,  �3���P  �3���  �����  �����P  �3���P      F  , ,  �����P  �����  �����  �����P  �����P      F  , ,  �k���P  �k���  �3���  �3���P  �k���P      F  , ,  ����P  ����  �����  �����P  ����P      F  , ,  ţ���P  ţ���  �k���  �k���P  ţ���P      F  , ,  �?���P  �?���  ����  ����P  �?���P      F  , ,  �����P  �����  ϣ���  ϣ���P  �����P      F  , ,  �3����  �3����  ������  ������  �3����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �k����  �k����  �3����  �3����  �k����      F  , ,  �����  �����  ������  ������  �����      F  , ,  ţ����  ţ����  �k����  �k����  ţ����      F  , ,  �?����  �?����  �����  �����  �?����      F  , ,  ������  ������  ϣ����  ϣ����  ������      F  , ,  �3���0  �3����  ������  �����0  �3���0      F  , ,  �����0  ������  ������  �����0  �����0      F  , ,  �k���0  �k����  �3����  �3���0  �k���0      F  , ,  ����0  �����  ������  �����0  ����0      F  , ,  ţ���0  ţ����  �k����  �k���0  ţ���0      F  , ,  �?���0  �?����  �����  ����0  �?���0      F  , ,  �����0  ������  ϣ����  ϣ���0  �����0      F  , ,  �3���<  �3���  �����  �����<  �3���<      F  , ,  �����<  �����  �����  �����<  �����<      F  , ,  �k���<  �k���  �3���  �3���<  �k���<      F  , ,  ����<  ����  �����  �����<  ����<      F  , ,  ţ���<  ţ���  �k���  �k���<  ţ���<      F  , ,  �?���<  �?���  ����  ����<  �?���<      F  , ,  �����<  �����  ϣ���  ϣ���<  �����<      F  , ,  �3����  �3���t  �����t  ������  �3����      F  , ,  ������  �����t  �����t  ������  ������      F  , ,  �k����  �k���t  �3���t  �3����  �k����      F  , ,  �����  ����t  �����t  ������  �����      F  , ,  ţ����  ţ���t  �k���t  �k����  ţ����      F  , ,  �?����  �?���t  ����t  �����  �?����      F  , ,  ������  �����t  ϣ���t  ϣ����  ������      F  , ,  �3���  �3����  ������  �����  �3���      F  , ,  �����  ������  ������  �����  �����      F  , ,  �k���  �k����  �3����  �3���  �k���      F  , ,  ����  �����  ������  �����  ����      F  , ,  ţ���  ţ����  �k����  �k���  ţ���      F  , ,  �?���  �?����  �����  ����  �?���      F  , ,  �����  ������  ϣ����  ϣ���  �����      F  , ,  �3����  �3���T  �����T  ������  �3����      F  , ,  ������  �����T  �����T  ������  ������      F  , ,  �k����  �k���T  �3���T  �3����  �k����      F  , ,  �����  ����T  �����T  ������  �����      F  , ,  ţ����  ţ���T  �k���T  �k����  ţ����      F  , ,  �?����  �?���T  ����T  �����  �?����      F  , ,  ������  �����T  ϣ���T  ϣ����  ������      F  , ,  �3����  �3����  ������  ������  �3����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �k����  �k����  �3����  �3����  �k����      F  , ,  �����  �����  ������  ������  �����      F  , ,  ţ����  ţ����  �k����  �k����  ţ����      F  , ,  �?����  �?����  �����  �����  �?����      F  , ,  ������  ������  ϣ����  ϣ����  ������      F  , ,  �3����  �3���X  �����X  ������  �3����      F  , ,  ������  �����X  �����X  ������  ������      F  , ,  �k����  �k���X  �3���X  �3����  �k����      F  , ,  �����  ����X  �����X  ������  �����      F  , ,  ţ����  ţ���X  �k���X  �k����  ţ����      F  , ,  �?����  �?���X  ����X  �����  �?����      F  , ,  ������  �����X  ϣ���X  ϣ����  ������      F  , ,  �3���   �3����  ������  �����   �3���       F  , ,  �����   ������  ������  �����   �����       F  , ,  �k���   �k����  �3����  �3���   �k���       F  , ,  ������  ������  ������  ������  ������      F  , ,  �_����  �_����  �'����  �'����  �_����      F  , ,  ������  ������  ������  ������  ������      F  , ,  ������  ������  �_����  �_����  ������      F  , ,  ������  �����^  �����^  ������  ������      F  , ,  �_����  �_���^  �'���^  �'����  �_����      F  , ,  ������  �����^  �����^  ������  ������      F  , ,  ������  �����^  �_���^  �_����  ������      F  , ,  ������  �����~  �_���~  �_����  ������      F  , ,  �_���F  �_���  �'���  �'���F  �_���F      F  , ,  �����F  �����  �����  �����F  �����F      F  , ,  �����F  �����  �_���  �_���F  �����F      F  , ,  �_���:  �_���  �'���  �'���:  �_���:      F  , ,  �����:  �����  �����  �����:  �����:      F  , ,  �����:  �����  �_���  �_���:  �����:      F  , ,  �'���  �'����  ������  �����  �'���      F  , ,  �����  ������  ������  �����  �����      F  , ,  �_���  �_����  �'����  �'���  �_���      F  , ,  �����  ������  ������  �����  �����      F  , ,  �����  ������  �_����  �_���  �����      F  , ,  �'���:  �'���  �����  �����:  �'���:      F  , ,  �'���&  �'����  ������  �����&  �'���&      F  , ,  �����&  ������  ������  �����&  �����&      F  , ,  �_���&  �_����  �'����  �'���&  �_���&      F  , ,  �����&  ������  ������  �����&  �����&      F  , ,  �����&  ������  �_����  �_���&  �����&      F  , ,  �����:  �����  �����  �����:  �����:      F  , ,  �'���v  �'���>  �����>  �����v  �'���v      F  , ,  �����v  �����>  �����>  �����v  �����v      F  , ,  �_���v  �_���>  �'���>  �'���v  �_���v      F  , ,  �����v  �����>  �����>  �����v  �����v      F  , ,  �����v  �����>  �_���>  �_���v  �����v      F  , ,  �'���F  �'���  �����  �����F  �'���F      F  , ,  �����F  �����  �����  �����F  �����F      F  , ,  �'����  �'���~  �����~  ������  �'����      F  , ,  �'���Z  �'���"  �����"  �����Z  �'���Z      F  , ,  �����Z  �����"  �����"  �����Z  �����Z      F  , ,  �_���Z  �_���"  �'���"  �'���Z  �_���Z      F  , ,  �����Z  �����"  �����"  �����Z  �����Z      F  , ,  �����Z  �����"  �_���"  �_���Z  �����Z      F  , ,  ������  �����~  �����~  ������  ������      F  , ,  �_����  �_���~  �'���~  �'����  �_����      F  , ,  ������  �����~  �����~  ������  ������      F  , ,  �'����  �'���^  �����^  ������  �'����      F  , ,  �'����  �'����  ������  ������  �'����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �_����  �_����  �'����  �'����  �_����      F  , ,  ������  ������  ������  ������  ������      F  , ,  ������  ������  �_����  �_����  ������      F  , ,  �'����  �'����  ������  ������  �'����      F  , ,  �_���0  �_����  �'����  �'���0  �_���0      F  , ,  �����0  ������  ������  �����0  �����0      F  , ,  �����0  ������  �_����  �_���0  �����0      F  , ,  �_����  �_���X  �'���X  �'����  �_����      F  , ,  �'���  �'����  ������  �����  �'���      F  , ,  �����  ������  ������  �����  �����      F  , ,  �_���  �_����  �'����  �'���  �_���      F  , ,  �����  ������  ������  �����  �����      F  , ,  �����  ������  �_����  �_���  �����      F  , ,  ������  �����X  �����X  ������  ������      F  , ,  �'���p  �'���8  �����8  �����p  �'���p      F  , ,  �����p  �����8  �����8  �����p  �����p      F  , ,  �_���p  �_���8  �'���8  �'���p  �_���p      F  , ,  �����p  �����8  �����8  �����p  �����p      F  , ,  �����p  �����8  �_���8  �_���p  �����p      F  , ,  ������  �����X  �_���X  �_����  ������      F  , ,  �'����  �'���T  �����T  ������  �'����      F  , ,  ������  �����T  �����T  ������  ������      F  , ,  �_����  �_���T  �'���T  �'����  �_����      F  , ,  ������  �����T  �����T  ������  ������      F  , ,  ������  �����T  �_���T  �_����  ������      F  , ,  �'����  �'����  ������  ������  �'����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �_����  �_����  �'����  �'����  �_����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �'���<  �'���  �����  �����<  �'���<      F  , ,  �����<  �����  �����  �����<  �����<      F  , ,  �'����  �'����  ������  ������  �'����      F  , ,  �'����  �'����  ������  ������  �'����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �_����  �_����  �'����  �'����  �_����      F  , ,  ������  ������  ������  ������  ������      F  , ,  ������  ������  �_����  �_����  ������      F  , ,  ������  ������  ������  ������  ������      F  , ,  �_����  �_����  �'����  �'����  �_����      F  , ,  ������  ������  ������  ������  ������      F  , ,  ������  ������  �_����  �_����  ������      F  , ,  �_���<  �_���  �'���  �'���<  �_���<      F  , ,  �����<  �����  �����  �����<  �����<      F  , ,  �����<  �����  �_���  �_���<  �����<      F  , ,  ������  ������  �_����  �_����  ������      F  , ,  �'����  �'���X  �����X  ������  �'����      F  , ,  ������  �����X  �����X  ������  ������      F  , ,  �'���   �'����  ������  �����   �'���       F  , ,  �����   ������  ������  �����   �����       F  , ,  �_���   �_����  �'����  �'���   �_���       F  , ,  �����   ������  ������  �����   �����       F  , ,  �'����  �'���t  �����t  ������  �'����      F  , ,  ������  �����t  �����t  ������  ������      F  , ,  �'���P  �'���  �����  �����P  �'���P      F  , ,  �����P  �����  �����  �����P  �����P      F  , ,  �_���P  �_���  �'���  �'���P  �_���P      F  , ,  �_����  �_���t  �'���t  �'����  �_����      F  , ,  ������  �����t  �����t  ������  ������      F  , ,  ������  �����t  �_���t  �_����  ������      F  , ,  �����   ������  �_����  �_���   �����       F  , ,  �'���0  �'����  ������  �����0  �'���0      F  , ,  �����P  �����  �����  �����P  �����P      F  , ,  �����P  �����  �_���  �_���P  �����P      F  , ,  �����0  ������  ������  �����0  �����0      F  , ,  �s��q�  �s��r�  �;��r�  �;��q�  �s��q�      F  , ,  ���q�  ���r�  ����r�  ����q�  ���q�      F  , ,  ����q�  ����r�  �s��r�  �s��q�  ����q�      F  , ,  �G��q�  �G��r�  ���r�  ���q�  �G��q�      F  , ,  �	��q�  �	��r�  ����r�  ����q�  �	��q�      F  , ,  ����q�  ����r�  �m��r�  �m��q�  ����q�      F  , ,  �A��q�  �A��r�  �	��r�  �	��q�  �A��q�      F  , ,  ����q�  ����r�  ����r�  ����q�  ����q�      F  , ,  �y��q�  �y��r�  �A��r�  �A��q�  �y��q�      F  , ,  �'���l  �'���4  �����4  �����l  �'���l      F  , ,  ����p1  ����p�  ����p�  ����p1  ����p1      F  , ,  �s��p1  �s��p�  �;��p�  �;��p1  �s��p1      F  , ,  ���p1  ���p�  ����p�  ����p1  ���p1      F  , ,  ����p1  ����p�  �s��p�  �s��p1  ����p1      F  , ,  �G��p1  �G��p�  ���p�  ���p1  �G��p1      F  , ,  �	��p1  �	��p�  ����p�  ����p1  �	��p1      F  , ,  ����p1  ����p�  �m��p�  �m��p1  ����p1      F  , ,  �A��p1  �A��p�  �	��p�  �	��p1  �A��p1      F  , ,  ����p1  ����p�  ����p�  ����p1  ����p1      F  , ,  �y��p1  �y��p�  �A��p�  �A��p1  �y��p1      F  , ,  �����l  �����4  �����4  �����l  �����l      F  , ,  ����n�  ����oi  ����oi  ����n�  ����n�      F  , ,  �s��n�  �s��oi  �;��oi  �;��n�  �s��n�      F  , ,  ���n�  ���oi  ����oi  ����n�  ���n�      F  , ,  ����n�  ����oi  �s��oi  �s��n�  ����n�      F  , ,  �G��n�  �G��oi  ���oi  ���n�  �G��n�      F  , ,  �	��n�  �	��oi  ����oi  ����n�  �	��n�      F  , ,  ����n�  ����oi  �m��oi  �m��n�  ����n�      F  , ,  �A��n�  �A��oi  �	��oi  �	��n�  �A��n�      F  , ,  ����n�  ����oi  ����oi  ����n�  ����n�      F  , ,  �y��n�  �y��oi  �A��oi  �A��n�  �y��n�      F  , ,  �_���l  �_���4  �'���4  �'���l  �_���l      F  , ,  ����m  ����m�  ����m�  ����m  ����m      F  , ,  �s��m  �s��m�  �;��m�  �;��m  �s��m      F  , ,  ���m  ���m�  ����m�  ����m  ���m      F  , ,  ����m  ����m�  �s��m�  �s��m  ����m      F  , ,  �G��m  �G��m�  ���m�  ���m  �G��m      F  , ,  �	��m  �	��m�  ����m�  ����m  �	��m      F  , ,  ����m  ����m�  �m��m�  �m��m  ����m      F  , ,  �A��m  �A��m�  �	��m�  �	��m  �A��m      F  , ,  ����m  ����m�  ����m�  ����m  ����m      F  , ,  �y��m  �y��m�  �A��m�  �A��m  �y��m      F  , ,  �����l  �����4  �����4  �����l  �����l      F  , ,  ����k�  ����lI  ����lI  ����k�  ����k�      F  , ,  �s��k�  �s��lI  �;��lI  �;��k�  �s��k�      F  , ,  ���k�  ���lI  ����lI  ����k�  ���k�      F  , ,  ����k�  ����lI  �s��lI  �s��k�  ����k�      F  , ,  �G��k�  �G��lI  ���lI  ���k�  �G��k�      F  , ,  �	��k�  �	��lI  ����lI  ����k�  �	��k�      F  , ,  ����k�  ����lI  �m��lI  �m��k�  ����k�      F  , ,  �A��k�  �A��lI  �	��lI  �	��k�  �A��k�      F  , ,  ����k�  ����lI  ����lI  ����k�  ����k�      F  , ,  �y��k�  �y��lI  �A��lI  �A��k�  �y��k�      F  , ,  �����l  �����4  �_���4  �_���l  �����l      F  , ,  ����i�  ����j�  ����j�  ����i�  ����i�      F  , ,  �s��i�  �s��j�  �;��j�  �;��i�  �s��i�      F  , ,  ���i�  ���j�  ����j�  ����i�  ���i�      F  , ,  ����i�  ����j�  �s��j�  �s��i�  ����i�      F  , ,  �G��i�  �G��j�  ���j�  ���i�  �G��i�      F  , ,  �	��i�  �	��j�  ����j�  ����i�  �	��i�      F  , ,  ����i�  ����j�  �m��j�  �m��i�  ����i�      F  , ,  �A��i�  �A��j�  �	��j�  �	��i�  �A��i�      F  , ,  ����i�  ����j�  ����j�  ����i�  ����i�      F  , ,  �y��i�  �y��j�  �A��j�  �A��i�  �y��i�      F  , ,  �'����  �'����  ������  ������  �'����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �_����  �_����  �'����  �'����  �_����      F  , ,  ������  ������  ������  ������  ������      F  , ,  ������  ������  �_����  �_����  ������      F  , ,  ����q�  ����r�  ����r�  ����q�  ����q�      F  , ,  y���k�  y���lI  zg��lI  zg��k�  y���k�      F  , ,  ~;��k�  ~;��lI  ��lI  ��k�  ~;��k�      F  , ,  y���n�  y���oi  zg��oi  zg��n�  y���n�      F  , ,  ~;��n�  ~;��oi  ��oi  ��n�  ~;��n�      F  , ,  ~;��p1  ~;��p�  ��p�  ��p1  ~;��p1      F  , ,  N���p�  N���q]  Ot��q]  Ot��p�  N���p�      F  , ,  u��p1  u��p�  u���p�  u���p1  u��p1      F  , ,  y���p1  y���p�  zg��p�  zg��p1  y���p1      F  , ,  u��m  u��m�  u���m�  u���m  u��m      F  , ,  y���m  y���m�  zg��m�  zg��m  y���m      F  , ,  ~;��m  ~;��m�  ��m�  ��m  ~;��m      F  , ,  u��n�  u��oi  u���oi  u���n�  u��n�      F  , ,  u��k�  u��lI  u���lI  u���k�  u��k�      F  , ,  u��i�  u��j�  u���j�  u���i�  u��i�      F  , ,  y���i�  y���j�  zg��j�  zg��i�  y���i�      F  , ,  N���y�  N���z�  Ot��z�  Ot��y�  N���y�      F  , ,  N���xe  N���y-  Ot��y-  Ot��xe  N���xe      F  , ,  N���v�  N���w�  Ot��w�  Ot��v�  N���v�      F  , ,  N���uE  N���v  Ot��v  Ot��uE  N���uE      F  , ,  N���s�  N���t}  Ot��t}  Ot��s�  N���s�      F  , ,  N���r%  N���r�  Ot��r�  Ot��r%  N���r%      F  , ,  u��q�  u��r�  u���r�  u���q�  u��q�      F  , ,  y���q�  y���r�  zg��r�  zg��q�  y���q�      F  , ,  ~;��q�  ~;��r�  ��r�  ��q�  ~;��q�      F  , ,  ~;��i�  ~;��j�  ��j�  ��i�  ~;��i�      F  , ,  y���^�  y���_o  zg��_o  zg��^�  y���^�      F  , ,  ~;��^�  ~;��_o  ��_o  ��^�  ~;��^�      F  , ,  u��]  u��]�  u���]�  u���]  u��]      F  , ,  y���]  y���]�  zg��]�  zg��]  y���]      F  , ,  ~;��]  ~;��]�  ��]�  ��]  ~;��]      F  , ,  u��[�  u��\O  u���\O  u���[�  u��[�      F  , ,  y���[�  y���\O  zg��\O  zg��[�  y���[�      F  , ,  ~;��[�  ~;��\O  ��\O  ��[�  ~;��[�      F  , ,  y���ha  y���i)  zg��i)  zg��ha  y���ha      F  , ,  u��Y�  u��Z�  u���Z�  u���Y�  u��Y�      F  , ,  y���Y�  y���Z�  zg��Z�  zg��Y�  y���Y�      F  , ,  ~;��Y�  ~;��Z�  ��Z�  ��Y�  ~;��Y�      F  , ,  ~;��ha  ~;��i)  ��i)  ��ha  ~;��ha      F  , ,  u��Xg  u��Y/  u���Y/  u���Xg  u��Xg      F  , ,  y���Xg  y���Y/  zg��Y/  zg��Xg  y���Xg      F  , ,  ~;��Xg  ~;��Y/  ��Y/  ��Xg  ~;��Xg      F  , ,  u��ha  u��i)  u���i)  u���ha  u��ha      F  , ,  u��a�  u��b�  u���b�  u���a�  u��a�      F  , ,  y���a�  y���b�  zg��b�  zg��a�  y���a�      F  , ,  ~;��a�  ~;��b�  ��b�  ��a�  ~;��a�      F  , ,  u��`7  u��`�  u���`�  u���`7  u��`7      F  , ,  y���`7  y���`�  zg��`�  zg��`7  y���`7      F  , ,  ~;��`7  ~;��`�  ��`�  ��`7  ~;��`7      F  , ,  u��^�  u��_o  u���_o  u���^�  u��^�      F  , ,  �	��`7  �	��`�  ����`�  ����`7  �	��`7      F  , ,  ����`7  ����`�  �m��`�  �m��`7  ����`7      F  , ,  �A��`7  �A��`�  �	��`�  �	��`7  �A��`7      F  , ,  ����`7  ����`�  ����`�  ����`7  ����`7      F  , ,  �y��`7  �y��`�  �A��`�  �A��`7  �y��`7      F  , ,  ����ha  ����i)  ����i)  ����ha  ����ha      F  , ,  �s��ha  �s��i)  �;��i)  �;��ha  �s��ha      F  , ,  ���ha  ���i)  ����i)  ����ha  ���ha      F  , ,  ����^�  ����_o  ����_o  ����^�  ����^�      F  , ,  �s��^�  �s��_o  �;��_o  �;��^�  �s��^�      F  , ,  ���^�  ���_o  ����_o  ����^�  ���^�      F  , ,  ����^�  ����_o  �s��_o  �s��^�  ����^�      F  , ,  �G��^�  �G��_o  ���_o  ���^�  �G��^�      F  , ,  �	��^�  �	��_o  ����_o  ����^�  �	��^�      F  , ,  ����^�  ����_o  �m��_o  �m��^�  ����^�      F  , ,  �A��^�  �A��_o  �	��_o  �	��^�  �A��^�      F  , ,  ����^�  ����_o  ����_o  ����^�  ����^�      F  , ,  �y��^�  �y��_o  �A��_o  �A��^�  �y��^�      F  , ,  ����ha  ����i)  �s��i)  �s��ha  ����ha      F  , ,  �G��ha  �G��i)  ���i)  ���ha  �G��ha      F  , ,  �	��ha  �	��i)  ����i)  ����ha  �	��ha      F  , ,  ����]  ����]�  ����]�  ����]  ����]      F  , ,  �s��]  �s��]�  �;��]�  �;��]  �s��]      F  , ,  ���]  ���]�  ����]�  ����]  ���]      F  , ,  ����]  ����]�  �s��]�  �s��]  ����]      F  , ,  �G��]  �G��]�  ���]�  ���]  �G��]      F  , ,  �	��]  �	��]�  ����]�  ����]  �	��]      F  , ,  ����]  ����]�  �m��]�  �m��]  ����]      F  , ,  �A��]  �A��]�  �	��]�  �	��]  �A��]      F  , ,  ����]  ����]�  ����]�  ����]  ����]      F  , ,  �y��]  �y��]�  �A��]�  �A��]  �y��]      F  , ,  ����ha  ����i)  �m��i)  �m��ha  ����ha      F  , ,  ����a�  ����b�  ����b�  ����a�  ����a�      F  , ,  �s��a�  �s��b�  �;��b�  �;��a�  �s��a�      F  , ,  ����[�  ����\O  ����\O  ����[�  ����[�      F  , ,  �s��[�  �s��\O  �;��\O  �;��[�  �s��[�      F  , ,  ���[�  ���\O  ����\O  ����[�  ���[�      F  , ,  ����[�  ����\O  �s��\O  �s��[�  ����[�      F  , ,  �G��[�  �G��\O  ���\O  ���[�  �G��[�      F  , ,  �	��[�  �	��\O  ����\O  ����[�  �	��[�      F  , ,  ����[�  ����\O  �m��\O  �m��[�  ����[�      F  , ,  �A��[�  �A��\O  �	��\O  �	��[�  �A��[�      F  , ,  ����[�  ����\O  ����\O  ����[�  ����[�      F  , ,  �y��[�  �y��\O  �A��\O  �A��[�  �y��[�      F  , ,  ���a�  ���b�  ����b�  ����a�  ���a�      F  , ,  ����a�  ����b�  �s��b�  �s��a�  ����a�      F  , ,  �G��a�  �G��b�  ���b�  ���a�  �G��a�      F  , ,  �	��a�  �	��b�  ����b�  ����a�  �	��a�      F  , ,  ����Y�  ����Z�  ����Z�  ����Y�  ����Y�      F  , ,  �s��Y�  �s��Z�  �;��Z�  �;��Y�  �s��Y�      F  , ,  ���Y�  ���Z�  ����Z�  ����Y�  ���Y�      F  , ,  ����Y�  ����Z�  �s��Z�  �s��Y�  ����Y�      F  , ,  �G��Y�  �G��Z�  ���Z�  ���Y�  �G��Y�      F  , ,  �	��Y�  �	��Z�  ����Z�  ����Y�  �	��Y�      F  , ,  ����Y�  ����Z�  �m��Z�  �m��Y�  ����Y�      F  , ,  �A��Y�  �A��Z�  �	��Z�  �	��Y�  �A��Y�      F  , ,  ����Y�  ����Z�  ����Z�  ����Y�  ����Y�      F  , ,  �y��Y�  �y��Z�  �A��Z�  �A��Y�  �y��Y�      F  , ,  ����a�  ����b�  �m��b�  �m��a�  ����a�      F  , ,  �A��a�  �A��b�  �	��b�  �	��a�  �A��a�      F  , ,  ����a�  ����b�  ����b�  ����a�  ����a�      F  , ,  �y��a�  �y��b�  �A��b�  �A��a�  �y��a�      F  , ,  ����Xg  ����Y/  ����Y/  ����Xg  ����Xg      F  , ,  �s��Xg  �s��Y/  �;��Y/  �;��Xg  �s��Xg      F  , ,  ���Xg  ���Y/  ����Y/  ����Xg  ���Xg      F  , ,  ����Xg  ����Y/  �s��Y/  �s��Xg  ����Xg      F  , ,  �G��Xg  �G��Y/  ���Y/  ���Xg  �G��Xg      F  , ,  �	��Xg  �	��Y/  ����Y/  ����Xg  �	��Xg      F  , ,  ����Xg  ����Y/  �m��Y/  �m��Xg  ����Xg      F  , ,  �A��Xg  �A��Y/  �	��Y/  �	��Xg  �A��Xg      F  , ,  ����Xg  ����Y/  ����Y/  ����Xg  ����Xg      F  , ,  �y��Xg  �y��Y/  �A��Y/  �A��Xg  �y��Xg      F  , ,  �A��ha  �A��i)  �	��i)  �	��ha  �A��ha      F  , ,  ����ha  ����i)  ����i)  ����ha  ����ha      F  , ,  �y��ha  �y��i)  �A��i)  �A��ha  �y��ha      F  , ,  ����`7  ����`�  ����`�  ����`7  ����`7      F  , ,  �s��`7  �s��`�  �;��`�  �;��`7  �s��`7      F  , ,  ���`7  ���`�  ����`�  ����`7  ���`7      F  , ,  ����`7  ����`�  �s��`�  �s��`7  ����`7      F  , ,  �G��`7  �G��`�  ���`�  ���`7  �G��`7      F  , ,  ����i�  ����j�  �k��j�  �k��i�  ����i�      F  , ,  �k��i�  �k��j�  �3��j�  �3��i�  �k��i�      F  , , 3��i� 3��j� ���j� ���i� 3��i�      F  , , ���i� ���j� 	���j� 	���i� ���i�      F  , , ���i� ���j� ���j� ���i� ���i�      F  , ,  ����nj  ����o2  �k��o2  �k��nj  ����nj      F  , ,  �k��nj  �k��o2  �3��o2  �3��nj  �k��nj      F  , , 3��nj 3��o2 ���o2 ���nj 3��nj      F  , , ���nj ���o2 	���o2 	���nj ���nj      F  , , ���nj ���o2 ���o2 ���nj ���nj      F  , ,  ����kJ  ����l  �k��l  �k��kJ  ����kJ      F  , ,  �k��kJ  �k��l  �3��l  �3��kJ  �k��kJ      F  , , 3��kJ 3��l ���l ���kJ 3��kJ      F  , , ���kJ ���l 	���l 	���kJ ���kJ      F  , , ���kJ ���l ���l ���kJ ���kJ      F  , ,  ����o�  ����p�  �k��p�  �k��o�  ����o�      F  , ,  �k��o�  �k��p�  �3��p�  �3��o�  �k��o�      F  , , 3��o� 3��p� ���p� ���o� 3��o�      F  , ,  ����l�  ����m�  �k��m�  �k��l�  ����l�      F  , ,  �k��l�  �k��m�  �3��m�  �3��l�  �k��l�      F  , , 3��l� 3��m� ���m� ���l� 3��l�      F  , , ���l� ���m� 	���m� 	���l� ���l�      F  , , ���l� ���m� ���m� ���l� ���l�      F  , , ���o� ���p� 	���p� 	���o� ���o�      F  , , ���o� ���p� ���p� ���o� ���o�      F  , ,  ����q�  ����rR  �k��rR  �k��q�  ����q�      F  , ,  �k��q�  �k��rR  �3��rR  �3��q�  �k��q�      F  , , 3��q� 3��rR ���rR ���q� 3��q�      F  , , ���q� ���rR 	���rR 	���q� ���q�      F  , , ���q� ���rR ���rR ���q� ���q�      F  , ,  ���k�  ���lI  ����lI  ����k�  ���k�      F  , ,  �3���l  �3���4  �����4  �����l  �3���l      F  , ,  �����l  �����4  �����4  �����l  �����l      F  , ,  �k���l  �k���4  �3���4  �3���l  �k���l      F  , ,  ���q�  ���r�  ����r�  ����q�  ���q�      F  , ,  ���p1  ���p�  ����p�  ����p1  ���p1      F  , ,  ����p1  ����p�  �y��p�  �y��p1  ����p1      F  , ,  �M��p1  �M��p�  ���p�  ���p1  �M��p1      F  , ,  ����k�  ����lI  �y��lI  �y��k�  ����k�      F  , ,  �M��k�  �M��lI  ���lI  ���k�  �M��k�      F  , ,  �k����  �k����  �3����  �3����  �k����      F  , ,  ���m  ���m�  ����m�  ����m  ���m      F  , ,  ����m  ����m�  �y��m�  �y��m  ����m      F  , ,  �M��m  �M��m�  ���m�  ���m  �M��m      F  , ,  �����  �����  ������  ������  �����      F  , ,  �?����  �?����  �����  �����  �?����      F  , ,  ������  ������  ϣ����  ϣ����  ������      F  , ,  �?���l  �?���4  ����4  ����l  �?���l      F  , ,  �����l  �����4  ϣ���4  ϣ���l  �����l      F  , ,  ���i�  ���j�  ����j�  ����i�  ���i�      F  , ,  ����i�  ����j�  �y��j�  �y��i�  ����i�      F  , ,  ����q�  ����r�  �y��r�  �y��q�  ����q�      F  , ,  �M��q�  �M��r�  ���r�  ���q�  �M��q�      F  , ,  �M��i�  �M��j�  ���j�  ���i�  �M��i�      F  , ,  ţ����  ţ����  �k����  �k����  ţ����      F  , ,  ���n�  ���oi  ����oi  ����n�  ���n�      F  , ,  ����n�  ����oi  �y��oi  �y��n�  ����n�      F  , ,  �M��n�  �M��oi  ���oi  ���n�  �M��n�      F  , ,  ����l  ����4  �����4  �����l  ����l      F  , ,  ţ���l  ţ���4  �k���4  �k���l  ţ���l      F  , ,  �3����  �3����  ������  ������  �3����      F  , ,  ������  ������  ������  ������  ������      F  , ,  �M��]  �M��]�  ���]�  ���]  �M��]      F  , ,  ���Y�  ���Z�  ����Z�  ����Y�  ���Y�      F  , ,  ����Y�  ����Z�  �y��Z�  �y��Y�  ����Y�      F  , ,  �M��Y�  �M��Z�  ���Z�  ���Y�  �M��Y�      F  , ,  �M��`7  �M��`�  ���`�  ���`7  �M��`7      F  , ,  ���`7  ���`�  ����`�  ����`7  ���`7      F  , ,  ���^�  ���_o  ����_o  ����^�  ���^�      F  , ,  ����^�  ����_o  �y��_o  �y��^�  ����^�      F  , ,  �M��^�  �M��_o  ���_o  ���^�  �M��^�      F  , ,  ����`7  ����`�  �y��`�  �y��`7  ����`7      F  , ,  ���ha  ���i)  ����i)  ����ha  ���ha      F  , ,  ����ha  ����i)  �y��i)  �y��ha  ����ha      F  , ,  �M��ha  �M��i)  ���i)  ���ha  �M��ha      F  , ,  ���Xg  ���Y/  ����Y/  ����Xg  ���Xg      F  , ,  ����Xg  ����Y/  �y��Y/  �y��Xg  ����Xg      F  , ,  �M��Xg  �M��Y/  ���Y/  ���Xg  �M��Xg      F  , ,  ���[�  ���\O  ����\O  ����[�  ���[�      F  , ,  ����[�  ����\O  �y��\O  �y��[�  ����[�      F  , ,  �M��[�  �M��\O  ���\O  ���[�  �M��[�      F  , ,  ���]  ���]�  ����]�  ����]  ���]      F  , ,  ����]  ����]�  �y��]�  �y��]  ����]      F  , ,  ���a�  ���b�  ����b�  ����a�  ���a�      F  , ,  ����a�  ����b�  �y��b�  �y��a�  ����a�      F  , ,  �M��a�  �M��b�  ���b�  ���a�  �M��a�      F  , ,  ����Yf  ����Z.  �k��Z.  �k��Yf  ����Yf      F  , ,  �k��Yf  �k��Z.  �3��Z.  �3��Yf  �k��Yf      F  , , 3��Yf 3��Z. ���Z. ���Yf 3��Yf      F  , , ���Yf ���Z. 	���Z. 	���Yf ���Yf      F  , , ���Yf ���Z. ���Z. ���Yf ���Yf      F  , ,  ����cz  ����dB  �k��dB  �k��cz  ����cz      F  , ,  �k��cz  �k��dB  �3��dB  �3��cz  �k��cz      F  , , 3��cz 3��dB ���dB ���cz 3��cz      F  , , ���cz ���dB 	���dB 	���cz ���cz      F  , , ���cz ���dB ���dB ���cz ���cz      F  , , 3��Z� 3��[� ���[� ���Z� 3��Z�      F  , , ���Z� ���[� 	���[� 	���Z� ���Z�      F  , , ���Z� ���[� ���[� ���Z� ���Z�      F  , , ���h* ���h� ���h� ���h* ���h*      F  , , ���h* ���h� 	���h� 	���h* ���h*      F  , ,  ����f�  ����gb  �k��gb  �k��f�  ����f�      F  , ,  �k��f�  �k��gb  �3��gb  �3��f�  �k��f�      F  , , 3��f� 3��gb ���gb ���f� 3��f�      F  , , ���f� ���gb 	���gb 	���f� ���f�      F  , , ���f� ���gb ���gb ���f� ���f�      F  , ,  ����h*  ����h�  �k��h�  �k��h*  ����h*      F  , ,  ����e
  ����e�  �k��e�  �k��e
  ����e
      F  , ,  ����W�  ����X�  �k��X�  �k��W�  ����W�      F  , ,  �k��W�  �k��X�  �3��X�  �3��W�  �k��W�      F  , , 3��W� 3��X� ���X� ���W� 3��W�      F  , , ���W� ���X� 	���X� 	���W� ���W�      F  , , ���W� ���X� ���X� ���W� ���W�      F  , ,  �k��e
  �k��e�  �3��e�  �3��e
  �k��e
      F  , ,  ����VF  ����W  �k��W  �k��VF  ����VF      F  , ,  �k��VF  �k��W  �3��W  �3��VF  �k��VF      F  , , 3��VF 3��W ���W ���VF 3��VF      F  , , ���VF ���W 	���W 	���VF ���VF      F  , , ���VF ���W ���W ���VF ���VF      F  , , 3��e
 3��e� ���e� ���e
 3��e
      F  , ,  ����T�  ����U~  �k��U~  �k��T�  ����T�      F  , ,  �k��T�  �k��U~  �3��U~  �3��T�  �k��T�      F  , , 3��T� 3��U~ ���U~ ���T� 3��T�      F  , , ���T� ���U~ 	���U~ 	���T� ���T�      F  , , ���T� ���U~ ���U~ ���T� ���T�      F  , , ���e
 ���e� 	���e� 	���e
 ���e
      F  , ,  ����S&  ����S�  �k��S�  �k��S&  ����S&      F  , ,  �k��S&  �k��S�  �3��S�  �3��S&  �k��S&      F  , , 3��S& 3��S� ���S� ���S& 3��S&      F  , , ���S& ���S� 	���S� 	���S& ���S&      F  , , ���S& ���S� ���S� ���S& ���S&      F  , , ���e
 ���e� ���e� ���e
 ���e
      F  , ,  ����Q�  ����R^  �k��R^  �k��Q�  ����Q�      F  , ,  �k��Q�  �k��R^  �3��R^  �3��Q�  �k��Q�      F  , , 3��Q� 3��R^ ���R^ ���Q� 3��Q�      F  , , ���Q� ���R^ 	���R^ 	���Q� ���Q�      F  , , ���Q� ���R^ ���R^ ���Q� ���Q�      F  , ,  �k��h*  �k��h�  �3��h�  �3��h*  �k��h*      F  , ,  ����P  ����P�  �k��P�  �k��P  ����P      F  , ,  �k��P  �k��P�  �3��P�  �3��P  �k��P      F  , , 3��P 3��P� ���P� ���P 3��P      F  , , ���P ���P� 	���P� 	���P ���P      F  , , ���P ���P� ���P� ���P ���P      F  , , 3��h* 3��h� ���h� ���h* 3��h*      F  , ,  ����Nv  ����O>  �k��O>  �k��Nv  ����Nv      F  , ,  �k��Nv  �k��O>  �3��O>  �3��Nv  �k��Nv      F  , , 3��Nv 3��O> ���O> ���Nv 3��Nv      F  , , ���Nv ���O> 	���O> 	���Nv ���Nv      F  , , ���Nv ���O> ���O> ���Nv ���Nv      F  , ,  ����Z�  ����[�  �k��[�  �k��Z�  ����Z�      F  , ,  ����L�  ����M�  �k��M�  �k��L�  ����L�      F  , ,  �k��L�  �k��M�  �3��M�  �3��L�  �k��L�      F  , , 3��L� 3��M� ���M� ���L� 3��L�      F  , , ���L� ���M� 	���M� 	���L� ���L�      F  , , ���L� ���M� ���M� ���L� ���L�      F  , ,  �k��Z�  �k��[�  �3��[�  �3��Z�  �k��Z�      F  , , S��i� S��j� ��j� ��i� S��i�      F  , ,  ��i�  ��j�  ���j�  ���i�  ��i�      F  , , %���i� %���j� &���j� &���i� %���i�      F  , , +���i� +���j� ,s��j� ,s��i� +���i�      F  , , 1s��i� 1s��j� 2;��j� 2;��i� 1s��i�      F  , , 7;��i� 7;��j� 8��j� 8��i� 7;��i�      F  , , =��i� =��j� =���j� =���i� =��i�      F  , , B���i� B���j� C���j� C���i� B���i�      F  , , H���i� H���j� I[��j� I[��i� H���i�      F  , , N[��i� N[��j� O#��j� O#��i� N[��i�      F  , , T#��i� T#��j� T���j� T���i� T#��i�      F  , , Y���i� Y���j� Z���j� Z���i� Y���i�      F  , , _���i� _���j� `{��j� `{��i� _���i�      F  , , e{��i� e{��j� fC��j� fC��i� e{��i�      F  , , kC��i� kC��j� l��j� l��i� kC��i�      F  , , q��i� q��j� q���j� q���i� q��i�      F  , , v���i� v���j� w���j� w���i� v���i�      F  , , _���o� _���p� `{��p� `{��o� _���o�      F  , , e{��o� e{��p� fC��p� fC��o� e{��o�      F  , , kC��o� kC��p� l��p� l��o� kC��o�      F  , , q��o� q��p� q���p� q���o� q��o�      F  , , v���o� v���p� w���p� w���o� v���o�      F  , , H���kJ H���l I[��l I[��kJ H���kJ      F  , , N[��kJ N[��l O#��l O#��kJ N[��kJ      F  , , T#��kJ T#��l T���l T���kJ T#��kJ      F  , , Y���kJ Y���l Z���l Z���kJ Y���kJ      F  , , _���kJ _���l `{��l `{��kJ _���kJ      F  , , e{��kJ e{��l fC��l fC��kJ e{��kJ      F  , , kC��kJ kC��l l��l l��kJ kC��kJ      F  , , q��kJ q��l q���l q���kJ q��kJ      F  , , v���kJ v���l w���l w���kJ v���kJ      F  , , H���q� H���rR I[��rR I[��q� H���q�      F  , , N[��q� N[��rR O#��rR O#��q� N[��q�      F  , , T#��q� T#��rR T���rR T���q� T#��q�      F  , , Y���q� Y���rR Z���rR Z���q� Y���q�      F  , , _���q� _���rR `{��rR `{��q� _���q�      F  , , e{��q� e{��rR fC��rR fC��q� e{��q�      F  , , kC��q� kC��rR l��rR l��q� kC��q�      F  , , q��q� q��rR q���rR q���q� q��q�      F  , , v���q� v���rR w���rR w���q� v���q�      F  , , H���o� H���p� I[��p� I[��o� H���o�      F  , , N[��o� N[��p� O#��p� O#��o� N[��o�      F  , , T#��o� T#��p� T���p� T���o� T#��o�      F  , , Y���o� Y���p� Z���p� Z���o� Y���o�      F  , , H���l� H���m� I[��m� I[��l� H���l�      F  , , N[��l� N[��m� O#��m� O#��l� N[��l�      F  , , T#��l� T#��m� T���m� T���l� T#��l�      F  , , Y���l� Y���m� Z���m� Z���l� Y���l�      F  , , _���l� _���m� `{��m� `{��l� _���l�      F  , , e{��l� e{��m� fC��m� fC��l� e{��l�      F  , , kC��l� kC��m� l��m� l��l� kC��l�      F  , , q��l� q��m� q���m� q���l� q��l�      F  , , v���l� v���m� w���m� w���l� v���l�      F  , , H���nj H���o2 I[��o2 I[��nj H���nj      F  , , N[��nj N[��o2 O#��o2 O#��nj N[��nj      F  , , T#��nj T#��o2 T���o2 T���nj T#��nj      F  , , Y���nj Y���o2 Z���o2 Z���nj Y���nj      F  , , _���nj _���o2 `{��o2 `{��nj _���nj      F  , , e{��nj e{��o2 fC��o2 fC��nj e{��nj      F  , , kC��nj kC��o2 l��o2 l��nj kC��nj      F  , , q��nj q��o2 q���o2 q���nj q��nj      F  , , v���nj v���o2 w���o2 w���nj v���nj      F  , , B���q� B���rR C���rR C���q� B���q�      F  , , +���o� +���p� ,s��p� ,s��o� +���o�      F  , , S��l� S��m� ��m� ��l� S��l�      F  , ,  ��l�  ��m�  ���m�  ���l�  ��l�      F  , , %���l� %���m� &���m� &���l� %���l�      F  , , +���l� +���m� ,s��m� ,s��l� +���l�      F  , , S��nj S��o2 ��o2 ��nj S��nj      F  , ,  ��nj  ��o2  ���o2  ���nj  ��nj      F  , , 1s��l� 1s��m� 2;��m� 2;��l� 1s��l�      F  , , 7;��l� 7;��m� 8��m� 8��l� 7;��l�      F  , , S��kJ S��l ��l ��kJ S��kJ      F  , ,  ��kJ  ��l  ���l  ���kJ  ��kJ      F  , , %���kJ %���l &���l &���kJ %���kJ      F  , , +���kJ +���l ,s��l ,s��kJ +���kJ      F  , , 1s��kJ 1s��l 2;��l 2;��kJ 1s��kJ      F  , , 7;��kJ 7;��l 8��l 8��kJ 7;��kJ      F  , , =��kJ =��l =���l =���kJ =��kJ      F  , , B���kJ B���l C���l C���kJ B���kJ      F  , , =��l� =��m� =���m� =���l� =��l�      F  , , B���l� B���m� C���m� C���l� B���l�      F  , , 1s��o� 1s��p� 2;��p� 2;��o� 1s��o�      F  , , 7;��o� 7;��p� 8��p� 8��o� 7;��o�      F  , , =��o� =��p� =���p� =���o� =��o�      F  , , B���o� B���p� C���p� C���o� B���o�      F  , , S��o� S��p� ��p� ��o� S��o�      F  , , %���nj %���o2 &���o2 &���nj %���nj      F  , , +���nj +���o2 ,s��o2 ,s��nj +���nj      F  , , 1s��nj 1s��o2 2;��o2 2;��nj 1s��nj      F  , , 7;��nj 7;��o2 8��o2 8��nj 7;��nj      F  , , =��nj =��o2 =���o2 =���nj =��nj      F  , , B���nj B���o2 C���o2 C���nj B���nj      F  , ,  ��o�  ��p�  ���p�  ���o�  ��o�      F  , , %���o� %���p� &���p� &���o� %���o�      F  , , S��q� S��rR ��rR ��q� S��q�      F  , ,  ��q�  ��rR  ���rR  ���q�  ��q�      F  , , %���q� %���rR &���rR &���q� %���q�      F  , , +���q� +���rR ,s��rR ,s��q� +���q�      F  , , 1s��q� 1s��rR 2;��rR 2;��q� 1s��q�      F  , , 7;��q� 7;��rR 8��rR 8��q� 7;��q�      F  , , =��q� =��rR =���rR =���q� =��q�      F  , , S��Z� S��[� ��[� ��Z� S��Z�      F  , ,  ��Z�  ��[�  ���[�  ���Z�  ��Z�      F  , , %���Z� %���[� &���[� &���Z� %���Z�      F  , , +���Z� +���[� ,s��[� ,s��Z� +���Z�      F  , , 1s��Z� 1s��[� 2;��[� 2;��Z� 1s��Z�      F  , , 7;��Z� 7;��[� 8��[� 8��Z� 7;��Z�      F  , , =��Z� =��[� =���[� =���Z� =��Z�      F  , , B���Z� B���[� C���[� C���Z� B���Z�      F  , , =��h* =��h� =���h� =���h* =��h*      F  , , B���h* B���h� C���h� C���h* B���h*      F  , , 1s��f� 1s��gb 2;��gb 2;��f� 1s��f�      F  , , 7;��f� 7;��gb 8��gb 8��f� 7;��f�      F  , , =��f� =��gb =���gb =���f� =��f�      F  , , B���f� B���gb C���gb C���f� B���f�      F  , , =��e
 =��e� =���e� =���e
 =��e
      F  , , B���e
 B���e� C���e� C���e
 B���e
      F  , , 1s��cz 1s��dB 2;��dB 2;��cz 1s��cz      F  , , 7;��cz 7;��dB 8��dB 8��cz 7;��cz      F  , , =��cz =��dB =���dB =���cz =��cz      F  , , B���cz B���dB C���dB C���cz B���cz      F  , , 1s��h* 1s��h� 2;��h� 2;��h* 1s��h*      F  , , 7;��h* 7;��h� 8��h� 8��h* 7;��h*      F  , , 1s��e
 1s��e� 2;��e� 2;��e
 1s��e
      F  , , 7;��e
 7;��e� 8��e� 8��e
 7;��e
      F  , , %���h* %���h� &���h� &���h* %���h*      F  , , +���h* +���h� ,s��h� ,s��h* +���h*      F  , , S��e
 S��e� ��e� ��e
 S��e
      F  , ,  ��e
  ��e�  ���e�  ���e
  ��e
      F  , , %���e
 %���e� &���e� &���e
 %���e
      F  , , S��f� S��gb ��gb ��f� S��f�      F  , ,  ��f�  ��gb  ���gb  ���f�  ��f�      F  , , %���f� %���gb &���gb &���f� %���f�      F  , , +���f� +���gb ,s��gb ,s��f� +���f�      F  , , S��cz S��dB ��dB ��cz S��cz      F  , ,  ��cz  ��dB  ���dB  ���cz  ��cz      F  , , %���cz %���dB &���dB &���cz %���cz      F  , , +���cz +���dB ,s��dB ,s��cz +���cz      F  , , +���e
 +���e� ,s��e� ,s��e
 +���e
      F  , , S��h* S��h� ��h� ��h* S��h*      F  , ,  ��h*  ��h�  ���h�  ���h*  ��h*      F  , , +���T� +���U~ ,s��U~ ,s��T� +���T�      F  , , S��S& S��S� ��S� ��S& S��S&      F  , ,  ��S&  ��S�  ���S�  ���S&  ��S&      F  , , %���S& %���S� &���S� &���S& %���S&      F  , , +���S& +���S� ,s��S� ,s��S& +���S&      F  , , +���W� +���X� ,s��X� ,s��W� +���W�      F  , , S��W� S��X� ��X� ��W� S��W�      F  , , S��Q� S��R^ ��R^ ��Q� S��Q�      F  , ,  ��Q�  ��R^  ���R^  ���Q�  ��Q�      F  , , %���Q� %���R^ &���R^ &���Q� %���Q�      F  , , +���Q� +���R^ ,s��R^ ,s��Q� +���Q�      F  , ,  ��W�  ��X�  ���X�  ���W�  ��W�      F  , , S��VF S��W ��W ��VF S��VF      F  , ,  ��VF  ��W  ���W  ���VF  ��VF      F  , , %���VF %���W &���W &���VF %���VF      F  , , +���VF +���W ,s��W ,s��VF +���VF      F  , , %���W� %���X� &���X� &���W� %���W�      F  , , S��P S��P� ��P� ��P S��P      F  , ,  ��P  ��P�  ���P�  ���P  ��P      F  , , %���P %���P� &���P� &���P %���P      F  , , +���P +���P� ,s��P� ,s��P +���P      F  , , S��T� S��U~ ��U~ ��T� S��T�      F  , ,  ��T�  ��U~  ���U~  ���T�  ��T�      F  , , %���T� %���U~ &���U~ &���T� %���T�      F  , , S��Yf S��Z. ��Z. ��Yf S��Yf      F  , ,  ��Yf  ��Z.  ���Z.  ���Yf  ��Yf      F  , , %���Yf %���Z. &���Z. &���Yf %���Yf      F  , , S��Nv S��O> ��O> ��Nv S��Nv      F  , ,  ��Nv  ��O>  ���O>  ���Nv  ��Nv      F  , , %���Nv %���O> &���O> &���Nv %���Nv      F  , , +���Nv +���O> ,s��O> ,s��Nv +���Nv      F  , , +���Yf +���Z. ,s��Z. ,s��Yf +���Yf      F  , , S��L� S��M� ��M� ��L� S��L�      F  , ,  ��L�  ��M�  ���M�  ���L�  ��L�      F  , , %���L� %���M� &���M� &���L� %���L�      F  , , +���L� +���M� ,s��M� ,s��L� +���L�      F  , , =��W� =��X� =���X� =���W� =��W�      F  , , 1s��T� 1s��U~ 2;��U~ 2;��T� 1s��T�      F  , , 7;��T� 7;��U~ 8��U~ 8��T� 7;��T�      F  , , =��T� =��U~ =���U~ =���T� =��T�      F  , , B���T� B���U~ C���U~ C���T� B���T�      F  , , B���W� B���X� C���X� C���W� B���W�      F  , , =��Yf =��Z. =���Z. =���Yf =��Yf      F  , , B���Yf B���Z. C���Z. C���Yf B���Yf      F  , , 1s��VF 1s��W 2;��W 2;��VF 1s��VF      F  , , 1s��P 1s��P� 2;��P� 2;��P 1s��P      F  , , 7;��P 7;��P� 8��P� 8��P 7;��P      F  , , =��P =��P� =���P� =���P =��P      F  , , B���P B���P� C���P� C���P B���P      F  , , 1s��S& 1s��S� 2;��S� 2;��S& 1s��S&      F  , , 7;��S& 7;��S� 8��S� 8��S& 7;��S&      F  , , =��S& =��S� =���S� =���S& =��S&      F  , , B���S& B���S� C���S� C���S& B���S&      F  , , 7;��VF 7;��W 8��W 8��VF 7;��VF      F  , , =��VF =��W =���W =���VF =��VF      F  , , B���VF B���W C���W C���VF B���VF      F  , , 1s��Yf 1s��Z. 2;��Z. 2;��Yf 1s��Yf      F  , , 7;��Yf 7;��Z. 8��Z. 8��Yf 7;��Yf      F  , , 1s��W� 1s��X� 2;��X� 2;��W� 1s��W�      F  , , 1s��Nv 1s��O> 2;��O> 2;��Nv 1s��Nv      F  , , 7;��Nv 7;��O> 8��O> 8��Nv 7;��Nv      F  , , =��Nv =��O> =���O> =���Nv =��Nv      F  , , B���Nv B���O> C���O> C���Nv B���Nv      F  , , 1s��Q� 1s��R^ 2;��R^ 2;��Q� 1s��Q�      F  , , 7;��Q� 7;��R^ 8��R^ 8��Q� 7;��Q�      F  , , =��Q� =��R^ =���R^ =���Q� =��Q�      F  , , B���Q� B���R^ C���R^ C���Q� B���Q�      F  , , 7;��W� 7;��X� 8��X� 8��W� 7;��W�      F  , , 1s��L� 1s��M� 2;��M� 2;��L� 1s��L�      F  , , 7;��L� 7;��M� 8��M� 8��L� 7;��L�      F  , , =��L� =��M� =���M� =���L� =��L�      F  , , B���L� B���M� C���M� C���L� B���L�      F  , , H���Z� H���[� I[��[� I[��Z� H���Z�      F  , , N[��Z� N[��[� O#��[� O#��Z� N[��Z�      F  , , T#��Z� T#��[� T���[� T���Z� T#��Z�      F  , , Y���Z� Y���[� Z���[� Z���Z� Y���Z�      F  , , _���Z� _���[� `{��[� `{��Z� _���Z�      F  , , e{��Z� e{��[� fC��[� fC��Z� e{��Z�      F  , , kC��Z� kC��[� l��[� l��Z� kC��Z�      F  , , q��Z� q��[� q���[� q���Z� q��Z�      F  , , v���Z� v���[� w���[� w���Z� v���Z�      F  , , kC��e
 kC��e� l��e� l��e
 kC��e
      F  , , q��e
 q��e� q���e� q���e
 q��e
      F  , , v���e
 v���e� w���e� w���e
 v���e
      F  , , _���f� _���gb `{��gb `{��f� _���f�      F  , , e{��f� e{��gb fC��gb fC��f� e{��f�      F  , , kC��f� kC��gb l��gb l��f� kC��f�      F  , , kC��cz kC��dB l��dB l��cz kC��cz      F  , , q��cz q��dB q���dB q���cz q��cz      F  , , v���cz v���dB w���dB w���cz v���cz      F  , , _���h* _���h� `{��h� `{��h* _���h*      F  , , e{��h* e{��h� fC��h� fC��h* e{��h*      F  , , kC��h* kC��h� l��h� l��h* kC��h*      F  , , q��h* q��h� q���h� q���h* q��h*      F  , , _���e
 _���e� `{��e� `{��e
 _���e
      F  , , e{��e
 e{��e� fC��e� fC��e
 e{��e
      F  , , q��f� q��gb q���gb q���f� q��f�      F  , , v���f� v���gb w���gb w���f� v���f�      F  , , v���h* v���h� w���h� w���h* v���h*      F  , , _���cz _���dB `{��dB `{��cz _���cz      F  , , e{��cz e{��dB fC��dB fC��cz e{��cz      F  , , Y���h* Y���h� Z���h� Z���h* Y���h*      F  , , N[��h* N[��h� O#��h� O#��h* N[��h*      F  , , H���f� H���gb I[��gb I[��f� H���f�      F  , , N[��f� N[��gb O#��gb O#��f� N[��f�      F  , , Y���f� Y���gb Z���gb Z���f� Y���f�      F  , , T#��f� T#��gb T���gb T���f� T#��f�      F  , , H���e
 H���e� I[��e� I[��e
 H���e
      F  , , N[��e
 N[��e� O#��e� O#��e
 N[��e
      F  , , T#��e
 T#��e� T���e� T���e
 T#��e
      F  , , H���h* H���h� I[��h� I[��h* H���h*      F  , , H���cz H���dB I[��dB I[��cz H���cz      F  , , N[��cz N[��dB O#��dB O#��cz N[��cz      F  , , T#��cz T#��dB T���dB T���cz T#��cz      F  , , Y���cz Y���dB Z���dB Z���cz Y���cz      F  , , Y���e
 Y���e� Z���e� Z���e
 Y���e
      F  , , T#��h* T#��h� T���h� T���h* T#��h*      F  , , Y���T� Y���U~ Z���U~ Z���T� Y���T�      F  , , T#��VF T#��W T���W T���VF T#��VF      F  , , Y���VF Y���W Z���W Z���VF Y���VF      F  , , N[��VF N[��W O#��W O#��VF N[��VF      F  , , H���Yf H���Z. I[��Z. I[��Yf H���Yf      F  , , H���W� H���X� I[��X� I[��W� H���W�      F  , , H���P H���P� I[��P� I[��P H���P      F  , , N[��P N[��P� O#��P� O#��P N[��P      F  , , T#��P T#��P� T���P� T���P T#��P      F  , , Y���P Y���P� Z���P� Z���P Y���P      F  , , N[��W� N[��X� O#��X� O#��W� N[��W�      F  , , T#��W� T#��X� T���X� T���W� T#��W�      F  , , Y���W� Y���X� Z���X� Z���W� Y���W�      F  , , N[��Yf N[��Z. O#��Z. O#��Yf N[��Yf      F  , , T#��Yf T#��Z. T���Z. T���Yf T#��Yf      F  , , H���Q� H���R^ I[��R^ I[��Q� H���Q�      F  , , N[��Q� N[��R^ O#��R^ O#��Q� N[��Q�      F  , , T#��Q� T#��R^ T���R^ T���Q� T#��Q�      F  , , Y���Q� Y���R^ Z���R^ Z���Q� Y���Q�      F  , , H���Nv H���O> I[��O> I[��Nv H���Nv      F  , , N[��Nv N[��O> O#��O> O#��Nv N[��Nv      F  , , T#��Nv T#��O> T���O> T���Nv T#��Nv      F  , , Y���Nv Y���O> Z���O> Z���Nv Y���Nv      F  , , Y���Yf Y���Z. Z���Z. Z���Yf Y���Yf      F  , , H���S& H���S� I[��S� I[��S& H���S&      F  , , N[��S& N[��S� O#��S� O#��S& N[��S&      F  , , T#��S& T#��S� T���S� T���S& T#��S&      F  , , Y���S& Y���S� Z���S� Z���S& Y���S&      F  , , H���T� H���U~ I[��U~ I[��T� H���T�      F  , , N[��T� N[��U~ O#��U~ O#��T� N[��T�      F  , , T#��T� T#��U~ T���U~ T���T� T#��T�      F  , , H���VF H���W I[��W I[��VF H���VF      F  , , H���L� H���M� I[��M� I[��L� H���L�      F  , , N[��L� N[��M� O#��M� O#��L� N[��L�      F  , , T#��L� T#��M� T���M� T���L� T#��L�      F  , , Y���L� Y���M� Z���M� Z���L� Y���L�      F  , , e{��P e{��P� fC��P� fC��P e{��P      F  , , kC��P kC��P� l��P� l��P kC��P      F  , , q��P q��P� q���P� q���P q��P      F  , , v���P v���P� w���P� w���P v���P      F  , , q��VF q��W q���W q���VF q��VF      F  , , _���T� _���U~ `{��U~ `{��T� _���T�      F  , , _���Q� _���R^ `{��R^ `{��Q� _���Q�      F  , , _���W� _���X� `{��X� `{��W� _���W�      F  , , e{��W� e{��X� fC��X� fC��W� e{��W�      F  , , kC��W� kC��X� l��X� l��W� kC��W�      F  , , q��W� q��X� q���X� q���W� q��W�      F  , , v���W� v���X� w���X� w���W� v���W�      F  , , e{��Q� e{��R^ fC��R^ fC��Q� e{��Q�      F  , , kC��Q� kC��R^ l��R^ l��Q� kC��Q�      F  , , q��Q� q��R^ q���R^ q���Q� q��Q�      F  , , v���Q� v���R^ w���R^ w���Q� v���Q�      F  , , e{��T� e{��U~ fC��U~ fC��T� e{��T�      F  , , _���S& _���S� `{��S� `{��S& _���S&      F  , , e{��S& e{��S� fC��S� fC��S& e{��S&      F  , , kC��S& kC��S� l��S� l��S& kC��S&      F  , , q��S& q��S� q���S� q���S& q��S&      F  , , v���S& v���S� w���S� w���S& v���S&      F  , , _���Nv _���O> `{��O> `{��Nv _���Nv      F  , , e{��Nv e{��O> fC��O> fC��Nv e{��Nv      F  , , kC��Nv kC��O> l��O> l��Nv kC��Nv      F  , , q��Nv q��O> q���O> q���Nv q��Nv      F  , , v���Nv v���O> w���O> w���Nv v���Nv      F  , , kC��T� kC��U~ l��U~ l��T� kC��T�      F  , , q��T� q��U~ q���U~ q���T� q��T�      F  , , v���T� v���U~ w���U~ w���T� v���T�      F  , , v���Yf v���Z. w���Z. w���Yf v���Yf      F  , , v���VF v���W w���W w���VF v���VF      F  , , _���Yf _���Z. `{��Z. `{��Yf _���Yf      F  , , e{��Yf e{��Z. fC��Z. fC��Yf e{��Yf      F  , , kC��Yf kC��Z. l��Z. l��Yf kC��Yf      F  , , q��Yf q��Z. q���Z. q���Yf q��Yf      F  , , _���VF _���W `{��W `{��VF _���VF      F  , , e{��VF e{��W fC��W fC��VF e{��VF      F  , , kC��VF kC��W l��W l��VF kC��VF      F  , , _���P _���P� `{��P� `{��P _���P      F  , , _���L� _���M� `{��M� `{��L� _���L�      F  , , e{��L� e{��M� fC��M� fC��L� e{��L�      F  , , kC��L� kC��M� l��M� l��L� kC��L�      F  , , q��L� q��M� q���M� q���L� q��L�      F  , , v���L� v���M� w���M� w���L� v���L�      F  , , |���i� |���j� }c��j� }c��i� |���i�      F  , , �c��i� �c��j� �+��j� �+��i� �c��i�      F  , , �+��i� �+��j� ����j� ����i� �+��i�      F  , , ����i� ����j� ����j� ����i� ����i�      F  , , ����i� ����j� ����j� ����i� ����i�      F  , , ����i� ����j� �K��j� �K��i� ����i�      F  , , �K��i� �K��j� ���j� ���i� �K��i�      F  , , ���i� ���j� ����j� ����i� ���i�      F  , , ����i� ����j� ����j� ����i� ����i�      F  , , ����i� ����j� �k��j� �k��i� ����i�      F  , , �k��i� �k��j� �3��j� �3��i� �k��i�      F  , , �3��i� �3��j� ����j� ����i� �3��i�      F  , , ����i� ����j� ����j� ����i� ����i�      F  , , ����i� ����j� ȋ��j� ȋ��i� ����i�      F  , , ͋��i� ͋��j� �S��j� �S��i� ͋��i�      F  , , ����l� ����m� �k��m� �k��l� ����l�      F  , , �k��l� �k��m� �3��m� �3��l� �k��l�      F  , , �3��l� �3��m� ����m� ����l� �3��l�      F  , , ����l� ����m� ����m� ����l� ����l�      F  , , ����l� ����m� ȋ��m� ȋ��l� ����l�      F  , , ͋��l� ͋��m� �S��m� �S��l� ͋��l�      F  , , ����o� ����p� ����p� ����o� ����o�      F  , , ����o� ����p� �k��p� �k��o� ����o�      F  , , �k��o� �k��p� �3��p� �3��o� �k��o�      F  , , �3��o� �3��p� ����p� ����o� �3��o�      F  , , ����o� ����p� ����p� ����o� ����o�      F  , , ����o� ����p� ȋ��p� ȋ��o� ����o�      F  , , ͋��o� ͋��p� �S��p� �S��o� ͋��o�      F  , , ����l� ����m� ����m� ����l� ����l�      F  , , ����kJ ����l ����l ����kJ ����kJ      F  , , ����kJ ����l �k��l �k��kJ ����kJ      F  , , �k��kJ �k��l �3��l �3��kJ �k��kJ      F  , , �3��kJ �3��l ����l ����kJ �3��kJ      F  , , ����kJ ����l ����l ����kJ ����kJ      F  , , ����kJ ����l ȋ��l ȋ��kJ ����kJ      F  , , ͋��kJ ͋��l �S��l �S��kJ ͋��kJ      F  , , ����q� ����rR ����rR ����q� ����q�      F  , , ����q� ����rR �k��rR �k��q� ����q�      F  , , �k��q� �k��rR �3��rR �3��q� �k��q�      F  , , �3��q� �3��rR ����rR ����q� �3��q�      F  , , ����q� ����rR ����rR ����q� ����q�      F  , , ����q� ����rR ȋ��rR ȋ��q� ����q�      F  , , ͋��q� ͋��rR �S��rR �S��q� ͋��q�      F  , , ����nj ����o2 ȋ��o2 ȋ��nj ����nj      F  , , ͋��nj ͋��o2 �S��o2 �S��nj ͋��nj      F  , , ����nj ����o2 ����o2 ����nj ����nj      F  , , ����nj ����o2 �k��o2 �k��nj ����nj      F  , , �k��nj �k��o2 �3��o2 �3��nj �k��nj      F  , , �3��nj �3��o2 ����o2 ����nj �3��nj      F  , , ����nj ����o2 ����o2 ����nj ����nj      F  , , �c��kJ �c��l �+��l �+��kJ �c��kJ      F  , , �+��kJ �+��l ����l ����kJ �+��kJ      F  , , �c��l� �c��m� �+��m� �+��l� �c��l�      F  , , �+��l� �+��m� ����m� ����l� �+��l�      F  , , ����l� ����m� ����m� ����l� ����l�      F  , , ����l� ����m� ����m� ����l� ����l�      F  , , ����kJ ����l ����l ����kJ ����kJ      F  , , ����kJ ����l ����l ����kJ ����kJ      F  , , ����kJ ����l �K��l �K��kJ ����kJ      F  , , �K��kJ �K��l ���l ���kJ �K��kJ      F  , , ���kJ ���l ����l ����kJ ���kJ      F  , , ����l� ����m� �K��m� �K��l� ����l�      F  , , �K��q� �K��rR ���rR ���q� �K��q�      F  , , ���q� ���rR ����rR ����q� ���q�      F  , , �K��l� �K��m� ���m� ���l� �K��l�      F  , , |���o� |���p� }c��p� }c��o� |���o�      F  , , �c��o� �c��p� �+��p� �+��o� �c��o�      F  , , �+��o� �+��p� ����p� ����o� �+��o�      F  , , ����o� ����p� ����p� ����o� ����o�      F  , , |���q� |���rR }c��rR }c��q� |���q�      F  , , �c��q� �c��rR �+��rR �+��q� �c��q�      F  , , �+��q� �+��rR ����rR ����q� �+��q�      F  , , ����q� ����rR ����rR ����q� ����q�      F  , , ����q� ����rR ����rR ����q� ����q�      F  , , ����q� ����rR �K��rR �K��q� ����q�      F  , , ����o� ����p� ����p� ����o� ����o�      F  , , ����o� ����p� �K��p� �K��o� ����o�      F  , , ���nj ���o2 ����o2 ����nj ���nj      F  , , �K��o� �K��p� ���p� ���o� �K��o�      F  , , ���o� ���p� ����p� ����o� ���o�      F  , , |���nj |���o2 }c��o2 }c��nj |���nj      F  , , �c��nj �c��o2 �+��o2 �+��nj �c��nj      F  , , �+��nj �+��o2 ����o2 ����nj �+��nj      F  , , ����nj ����o2 ����o2 ����nj ����nj      F  , , ����nj ����o2 ����o2 ����nj ����nj      F  , , ���l� ���m� ����m� ����l� ���l�      F  , , |���l� |���m� }c��m� }c��l� |���l�      F  , , |���kJ |���l }c��l }c��kJ |���kJ      F  , , �K��nj �K��o2 ���o2 ���nj �K��nj      F  , , ����nj ����o2 �K��o2 �K��nj ����nj      F  , , |���Z� |���[� }c��[� }c��Z� |���Z�      F  , , �c��Z� �c��[� �+��[� �+��Z� �c��Z�      F  , , �+��Z� �+��[� ����[� ����Z� �+��Z�      F  , , ����Z� ����[� ����[� ����Z� ����Z�      F  , , ����Z� ����[� ����[� ����Z� ����Z�      F  , , ����Z� ����[� �K��[� �K��Z� ����Z�      F  , , �K��Z� �K��[� ���[� ���Z� �K��Z�      F  , , ���Z� ���[� ����[� ����Z� ���Z�      F  , , ����f� ����gb ����gb ����f� ����f�      F  , , ����f� ����gb �K��gb �K��f� ����f�      F  , , �K��f� �K��gb ���gb ���f� �K��f�      F  , , ���f� ���gb ����gb ����f� ���f�      F  , , ����e
 ����e� �K��e� �K��e
 ����e
      F  , , �K��e
 �K��e� ���e� ���e
 �K��e
      F  , , ���e
 ���e� ����e� ����e
 ���e
      F  , , ����h* ����h� ����h� ����h* ����h*      F  , , ����h* ����h� �K��h� �K��h* ����h*      F  , , �K��h* �K��h� ���h� ���h* �K��h*      F  , , ���h* ���h� ����h� ����h* ���h*      F  , , ����cz ����dB ����dB ����cz ����cz      F  , , ����cz ����dB �K��dB �K��cz ����cz      F  , , �K��cz �K��dB ���dB ���cz �K��cz      F  , , ���cz ���dB ����dB ����cz ���cz      F  , , ����e
 ����e� ����e� ����e
 ����e
      F  , , ����f� ����gb ����gb ����f� ����f�      F  , , |���cz |���dB }c��dB }c��cz |���cz      F  , , |���e
 |���e� }c��e� }c��e
 |���e
      F  , , �c��e
 �c��e� �+��e� �+��e
 �c��e
      F  , , �+��e
 �+��e� ����e� ����e
 �+��e
      F  , , |���f� |���gb }c��gb }c��f� |���f�      F  , , �c��cz �c��dB �+��dB �+��cz �c��cz      F  , , �+��cz �+��dB ����dB ����cz �+��cz      F  , , ����e
 ����e� ����e� ����e
 ����e
      F  , , ����cz ����dB ����dB ����cz ����cz      F  , , �+��f� �+��gb ����gb ����f� �+��f�      F  , , �c��f� �c��gb �+��gb �+��f� �c��f�      F  , , |���h* |���h� }c��h� }c��h* |���h*      F  , , �c��h* �c��h� �+��h� �+��h* �c��h*      F  , , �+��h* �+��h� ����h� ����h* �+��h*      F  , , ����h* ����h� ����h� ����h* ����h*      F  , , �+��Q� �+��R^ ����R^ ����Q� �+��Q�      F  , , ����Q� ����R^ ����R^ ����Q� ����Q�      F  , , |���T� |���U~ }c��U~ }c��T� |���T�      F  , , �c��T� �c��U~ �+��U~ �+��T� �c��T�      F  , , �+��T� �+��U~ ����U~ ����T� �+��T�      F  , , ����S& ����S� ����S� ����S& ����S&      F  , , |���VF |���W }c��W }c��VF |���VF      F  , , �c��VF �c��W �+��W �+��VF �c��VF      F  , , �+��VF �+��W ����W ����VF �+��VF      F  , , |���P |���P� }c��P� }c��P |���P      F  , , �c��P �c��P� �+��P� �+��P �c��P      F  , , �+��P �+��P� ����P� ����P �+��P      F  , , ����P ����P� ����P� ����P ����P      F  , , ����T� ����U~ ����U~ ����T� ����T�      F  , , |���Yf |���Z. }c��Z. }c��Yf |���Yf      F  , , �c��Yf �c��Z. �+��Z. �+��Yf �c��Yf      F  , , �+��Yf �+��Z. ����Z. ����Yf �+��Yf      F  , , ����Yf ����Z. ����Z. ����Yf ����Yf      F  , , |���Nv |���O> }c��O> }c��Nv |���Nv      F  , , �c��Nv �c��O> �+��O> �+��Nv �c��Nv      F  , , �+��Nv �+��O> ����O> ����Nv �+��Nv      F  , , ����Nv ����O> ����O> ����Nv ����Nv      F  , , ����VF ����W ����W ����VF ����VF      F  , , |���W� |���X� }c��X� }c��W� |���W�      F  , , �c��W� �c��X� �+��X� �+��W� �c��W�      F  , , �+��W� �+��X� ����X� ����W� �+��W�      F  , , ����W� ����X� ����X� ����W� ����W�      F  , , |���S& |���S� }c��S� }c��S& |���S&      F  , , �c��S& �c��S� �+��S� �+��S& �c��S&      F  , , �+��S& �+��S� ����S� ����S& �+��S&      F  , , |���Q� |���R^ }c��R^ }c��Q� |���Q�      F  , , �c��Q� �c��R^ �+��R^ �+��Q� �c��Q�      F  , , |���L� |���M� }c��M� }c��L� |���L�      F  , , �c��L� �c��M� �+��M� �+��L� �c��L�      F  , , �+��L� �+��M� ����M� ����L� �+��L�      F  , , ����L� ����M� ����M� ����L� ����L�      F  , , ����S& ����S� ����S� ����S& ����S&      F  , , ����S& ����S� �K��S� �K��S& ����S&      F  , , ����Yf ����Z. ����Z. ����Yf ����Yf      F  , , ����Yf ����Z. �K��Z. �K��Yf ����Yf      F  , , �K��Yf �K��Z. ���Z. ���Yf �K��Yf      F  , , �K��S& �K��S� ���S� ���S& �K��S&      F  , , ����Q� ����R^ ����R^ ����Q� ����Q�      F  , , ����Q� ����R^ �K��R^ �K��Q� ����Q�      F  , , �K��Q� �K��R^ ���R^ ���Q� �K��Q�      F  , , ����Nv ����O> ����O> ����Nv ����Nv      F  , , ����Nv ����O> �K��O> �K��Nv ����Nv      F  , , �K��Nv �K��O> ���O> ���Nv �K��Nv      F  , , ���Nv ���O> ����O> ����Nv ���Nv      F  , , ���Yf ���Z. ����Z. ����Yf ���Yf      F  , , ���Q� ���R^ ����R^ ����Q� ���Q�      F  , , ����VF ����W �K��W �K��VF ����VF      F  , , �K��VF �K��W ���W ���VF �K��VF      F  , , ����P ����P� ����P� ����P ����P      F  , , ����P ����P� �K��P� �K��P ����P      F  , , ����W� ����X� ����X� ����W� ����W�      F  , , ����W� ����X� �K��X� �K��W� ����W�      F  , , �K��W� �K��X� ���X� ���W� �K��W�      F  , , ���W� ���X� ����X� ����W� ���W�      F  , , �K��P �K��P� ���P� ���P �K��P      F  , , ���P ���P� ����P� ����P ���P      F  , , ���VF ���W ����W ����VF ���VF      F  , , ����T� ����U~ ����U~ ����T� ����T�      F  , , ����T� ����U~ �K��U~ �K��T� ����T�      F  , , �K��T� �K��U~ ���U~ ���T� �K��T�      F  , , ���T� ���U~ ����U~ ����T� ���T�      F  , , ����VF ����W ����W ����VF ����VF      F  , , ���S& ���S� ����S� ����S& ���S&      F  , , ����L� ����M� ����M� ����L� ����L�      F  , , ����L� ����M� �K��M� �K��L� ����L�      F  , , �K��L� �K��M� ���M� ���L� �K��L�      F  , , ���L� ���M� ����M� ����L� ���L�      F  , , ����Z� ����[� ����[� ����Z� ����Z�      F  , , ����Z� ����[� �k��[� �k��Z� ����Z�      F  , , �k��Z� �k��[� �3��[� �3��Z� �k��Z�      F  , , �3��Z� �3��[� ����[� ����Z� �3��Z�      F  , , ����Z� ����[� ����[� ����Z� ����Z�      F  , , ����Z� ����[� ȋ��[� ȋ��Z� ����Z�      F  , , ͋��Z� ͋��[� �S��[� �S��Z� ͋��Z�      F  , , ͋��f� ͋��gb �S��gb �S��f� ͋��f�      F  , , ����f� ����g� ۖ��g� ۖ��f� ����f�      F  , , ����h ����iG ۖ��iG ۖ��h ����h      F  , , ����f� ����gb ȋ��gb ȋ��f� ����f�      F  , , ����[� ����\� ۖ��\� ۖ��[� ����[�      F  , , ����h* ����h� ȋ��h� ȋ��h* ����h*      F  , , ͋��h* ͋��h� �S��h� �S��h* ͋��h*      F  , , ����cz ����dB ȋ��dB ȋ��cz ����cz      F  , , ͋��cz ͋��dB �S��dB �S��cz ͋��cz      F  , , ����c� ����d� ۖ��d� ۖ��c� ����c�      F  , , ����_ ����_� ۖ��_� ۖ��_ ����_      F  , , ����`� ����aw ۖ��aw ۖ��`� ����`�      F  , , ����]� ����^W ۖ��^W ۖ��]� ����]�      F  , , ����b? ����c ۖ��c ۖ��b? ����b?      F  , , ����e
 ����e� ȋ��e� ȋ��e
 ����e
      F  , , ͋��e
 ͋��e� �S��e� �S��e
 ͋��e
      F  , , ����e_ ����f' ۖ��f' ۖ��e_ ����e_      F  , , ����cz ����dB �k��dB �k��cz ����cz      F  , , �k��cz �k��dB �3��dB �3��cz �k��cz      F  , , �3��cz �3��dB ����dB ����cz �3��cz      F  , , ����cz ����dB ����dB ����cz ����cz      F  , , ����f� ����gb ����gb ����f� ����f�      F  , , ����f� ����gb ����gb ����f� ����f�      F  , , ����e
 ����e� �k��e� �k��e
 ����e
      F  , , �k��h* �k��h� �3��h� �3��h* �k��h*      F  , , ����h* ����h� ����h� ����h* ����h*      F  , , ����e
 ����e� ����e� ����e
 ����e
      F  , , ����f� ����gb �k��gb �k��f� ����f�      F  , , �k��f� �k��gb �3��gb �3��f� �k��f�      F  , , �k��e
 �k��e� �3��e� �3��e
 �k��e
      F  , , ����h* ����h� ����h� ����h* ����h*      F  , , �3��e
 �3��e� ����e� ����e
 �3��e
      F  , , ����e
 ����e� ����e� ����e
 ����e
      F  , , ����h* ����h� �k��h� �k��h* ����h*      F  , , �3��f� �3��gb ����gb ����f� �3��f�      F  , , ����cz ����dB ����dB ����cz ����cz      F  , , �3��h* �3��h� ����h� ����h* �3��h*      F  , , ����T� ����U~ �k��U~ �k��T� ����T�      F  , , �k��T� �k��U~ �3��U~ �3��T� �k��T�      F  , , �3��T� �3��U~ ����U~ ����T� �3��T�      F  , , ����T� ����U~ ����U~ ����T� ����T�      F  , , �3��P �3��P� ����P� ����P �3��P      F  , , ����P ����P� ����P� ����P ����P      F  , , ����W� ����X� ����X� ����W� ����W�      F  , , ����W� ����X� ����X� ����W� ����W�      F  , , ����W� ����X� �k��X� �k��W� ����W�      F  , , �k��W� �k��X� �3��X� �3��W� �k��W�      F  , , ����Nv ����O> ����O> ����Nv ����Nv      F  , , ����Nv ����O> �k��O> �k��Nv ����Nv      F  , , �k��Nv �k��O> �3��O> �3��Nv �k��Nv      F  , , �3��Nv �3��O> ����O> ����Nv �3��Nv      F  , , ����Nv ����O> ����O> ����Nv ����Nv      F  , , �3��W� �3��X� ����X� ����W� �3��W�      F  , , ����S& ����S� ����S� ����S& ����S&      F  , , ����S& ����S� �k��S� �k��S& ����S&      F  , , �k��S& �k��S� �3��S� �3��S& �k��S&      F  , , ����Yf ����Z. ����Z. ����Yf ����Yf      F  , , ����Yf ����Z. �k��Z. �k��Yf ����Yf      F  , , �k��Yf �k��Z. �3��Z. �3��Yf �k��Yf      F  , , �3��Yf �3��Z. ����Z. ����Yf �3��Yf      F  , , ����Yf ����Z. ����Z. ����Yf ����Yf      F  , , �3��S& �3��S� ����S� ����S& �3��S&      F  , , ����S& ����S� ����S� ����S& ����S&      F  , , ����P ����P� ����P� ����P ����P      F  , , ����P ����P� �k��P� �k��P ����P      F  , , ����Q� ����R^ ����R^ ����Q� ����Q�      F  , , ����Q� ����R^ �k��R^ �k��Q� ����Q�      F  , , �k��Q� �k��R^ �3��R^ �3��Q� �k��Q�      F  , , �3��Q� �3��R^ ����R^ ����Q� �3��Q�      F  , , �k��P �k��P� �3��P� �3��P �k��P      F  , , ����Q� ����R^ ����R^ ����Q� ����Q�      F  , , ����VF ����W ����W ����VF ����VF      F  , , ����VF ����W �k��W �k��VF ����VF      F  , , �k��VF �k��W �3��W �3��VF �k��VF      F  , , �3��VF �3��W ����W ����VF �3��VF      F  , , ����VF ����W ����W ����VF ����VF      F  , , ����T� ����U~ ����U~ ����T� ����T�      F  , , ����L� ����M� ����M� ����L� ����L�      F  , , ����L� ����M� �k��M� �k��L� ����L�      F  , , �k��L� �k��M� �3��M� �3��L� �k��L�      F  , , �3��L� �3��M� ����M� ����L� �3��L�      F  , , ����L� ����M� ����M� ����L� ����L�      F  , , ͋��P ͋��P� �S��P� �S��P ͋��P      F  , , ����W� ����X� ȋ��X� ȋ��W� ����W�      F  , , ����Zo ����[7 ۖ��[7 ۖ��Zo ����Zo      F  , , ����T� ����U~ ȋ��U~ ȋ��T� ����T�      F  , , ����Q� ����R^ ȋ��R^ ȋ��Q� ����Q�      F  , , ͋��Q� ͋��R^ �S��R^ �S��Q� ͋��Q�      F  , , ͋��T� ͋��U~ �S��U~ �S��T� ͋��T�      F  , , ����S& ����S� ȋ��S� ȋ��S& ����S&      F  , , ͋��S& ͋��S� �S��S� �S��S& ͋��S&      F  , , ����Yf ����Z. ȋ��Z. ȋ��Yf ����Yf      F  , , ͋��Yf ͋��Z. �S��Z. �S��Yf ͋��Yf      F  , , ����Nv ����O> ȋ��O> ȋ��Nv ����Nv      F  , , ͋��Nv ͋��O> �S��O> �S��Nv ͋��Nv      F  , , ͋��W� ͋��X� �S��X� �S��W� ͋��W�      F  , , ����VF ����W ȋ��W ȋ��VF ����VF      F  , , ͋��VF ͋��W �S��W �S��VF ͋��VF      F  , , ����P ����P� ȋ��P� ȋ��P ����P      F  , , ����L� ����M� ȋ��M� ȋ��L� ����L�      F  , , ͋��L� ͋��M� �S��M� �S��L� ͋��L�      D  , , 2��_� 2��`� ���`� ���_� 2��_�      D  , , 2��^� 2��_G ���_G ���^� 2��^�      D  , , �-  &� �-  '[ ��  '[ ��  &� �-  &�      D  , , �-  %� �-  & ��  & ��  %� �-  %�      D  , , ��  2� ��  3E Ȇ  3E Ȇ  2� ��  2�      D  , , �>  2� �>  3E ��  3E ��  2� �>  2�      D  , , ̌  2� ̌  3E �"  3E �"  2� ̌  2�      D  , , ��  2� ��  3E �p  3E �p  2� ��  2�      D  , , �T  1o �T  2 ��  2 ��  1o �T  1o      D  , , Ţ  1o Ţ  2 �8  2 �8  1o Ţ  1o      D  , , ��  1o ��  2 Ȇ  2 Ȇ  1o ��  1o      D  , , �>  1o �>  2 ��  2 ��  1o �>  1o      D  , , ̌  1o ̌  2 �"  2 �"  1o ̌  1o      D  , , ��  1o ��  2 �p  2 �p  1o ��  1o      D  , , �T  0/ �T  0� ��  0� ��  0/ �T  0/      D  , , Ţ  0/ Ţ  0� �8  0� �8  0/ Ţ  0/      D  , , ��  0/ ��  0� Ȇ  0� Ȇ  0/ ��  0/      D  , , �>  0/ �>  0� ��  0� ��  0/ �>  0/      D  , , ̌  0/ ̌  0� �"  0� �"  0/ ̌  0/      D  , , ��  0/ ��  0� �p  0� �p  0/ ��  0/      D  , , �T  .� �T  /� ��  /� ��  .� �T  .�      D  , , Ţ  .� Ţ  /� �8  /� �8  .� Ţ  .�      D  , , ��  .� ��  /� Ȇ  /� Ȇ  .� ��  .�      D  , , �>  .� �>  /� ��  /� ��  .� �>  .�      D  , , ̌  .� ̌  /� �"  /� �"  .� ̌  .�      D  , , ��  .� ��  /� �p  /� �p  .� ��  .�      D  , , �T  -� �T  .E ��  .E ��  -� �T  -�      D  , , Ţ  -� Ţ  .E �8  .E �8  -� Ţ  -�      D  , , ��  -� ��  .E Ȇ  .E Ȇ  -� ��  -�      D  , , �>  -� �>  .E ��  .E ��  -� �>  -�      D  , , ̌  -� ̌  .E �"  .E �"  -� ̌  -�      D  , , ��  -� ��  .E �p  .E �p  -� ��  -�      D  , , �T  ,o �T  - ��  - ��  ,o �T  ,o      D  , , Ţ  ,o Ţ  - �8  - �8  ,o Ţ  ,o      D  , , ��  ,o ��  - Ȇ  - Ȇ  ,o ��  ,o      D  , , �>  ,o �>  - ��  - ��  ,o �>  ,o      D  , , ̌  ,o ̌  - �"  - �"  ,o ̌  ,o      D  , , ��  ,o ��  - �p  - �p  ,o ��  ,o      D  , , �T  +/ �T  +� ��  +� ��  +/ �T  +/      D  , , Ţ  +/ Ţ  +� �8  +� �8  +/ Ţ  +/      D  , , ��  +/ ��  +� Ȇ  +� Ȇ  +/ ��  +/      D  , , �>  +/ �>  +� ��  +� ��  +/ �>  +/      D  , , ̌  +/ ̌  +� �"  +� �"  +/ ̌  +/      D  , , ��  +/ ��  +� �p  +� �p  +/ ��  +/      D  , , �T  )� �T  *� ��  *� ��  )� �T  )�      D  , , Ţ  )� Ţ  *� �8  *� �8  )� Ţ  )�      D  , , ��  )� ��  *� Ȇ  *� Ȇ  )� ��  )�      D  , , �>  )� �>  *� ��  *� ��  )� �>  )�      D  , , ̌  )� ̌  *� �"  *� �"  )� ̌  )�      D  , , ��  )� ��  *� �p  *� �p  )� ��  )�      D  , , �T  2� �T  3E ��  3E ��  2� �T  2�      D  , , �{  &� �{  '[ �  '[ �  &� �{  &�      D  , , ��  &� ��  '[ �_  '[ �_  &� ��  &�      D  , , �  &� �  '[ ɭ  '[ ɭ  &� �  &�      D  , , �e  &� �e  '[ ��  '[ ��  &� �e  &�      D  , , ͳ  &� ͳ  '[ �I  '[ �I  &� ͳ  &�      D  , , Ţ  2� Ţ  3E �8  3E �8  2� Ţ  2�      D  , , �{  %� �{  & �  & �  %� �{  %�      D  , , ��  %� ��  & �_  & �_  %� ��  %�      D  , , �  %� �  & ɭ  & ɭ  %� �  %�      D  , , �e  %� �e  & ��  & ��  %� �e  %�      D  , , ͳ  %� ͳ  & �I  & �I  %� ͳ  %�      D  , , ��  1o ��  2 �  2 �  1o ��  1o      D  , , ��  -� ��  .E �  .E �  -� ��  -�      D  , , ��  ,o ��  - �  - �  ,o ��  ,o      D  , , ��  +/ ��  +� �  +� �  +/ ��  +/      D  , , ��  0/ ��  0� �  0� �  0/ ��  0/      D  , , ��  )� ��  *� �  *� �  )� ��  )�      D  , , ��  2� ��  3E �  3E �  2� ��  2�      D  , , ��  .� ��  /� �  /� �  .� ��  .�      D  , , ��  -� ��  .E �N  .E �N  -� ��  -�      D  , , �  -� �  .E ��  .E ��  -� �  -�      D  , , �  1o �  2 ��  2 ��  1o �  1o      D  , , �j  1o �j  2 �   2 �   1o �j  1o      D  , , ��  1o ��  2 �N  2 �N  1o ��  1o      D  , , �  1o �  2 ��  2 ��  1o �  1o      D  , , ��  2� ��  3E �d  3E �d  2� ��  2�      D  , , �  2� �  3E ��  3E ��  2� �  2�      D  , , ��  .� ��  /� �N  /� �N  .� ��  .�      D  , , ��  ,o ��  - �d  - �d  ,o ��  ,o      D  , , �  ,o �  - ��  - ��  ,o �  ,o      D  , , �j  ,o �j  - �   - �   ,o �j  ,o      D  , , ��  ,o ��  - �N  - �N  ,o ��  ,o      D  , , �  ,o �  - ��  - ��  ,o �  ,o      D  , , �j  2� �j  3E �   3E �   2� �j  2�      D  , , ��  2� ��  3E �N  3E �N  2� ��  2�      D  , , �  2� �  3E ��  3E ��  2� �  2�      D  , , ��  1o ��  2 �d  2 �d  1o ��  1o      D  , , �  .� �  /� ��  /� ��  .� �  .�      D  , , ��  0/ ��  0� �d  0� �d  0/ ��  0/      D  , , �  0/ �  0� ��  0� ��  0/ �  0/      D  , , ��  -� ��  .E �d  .E �d  -� ��  -�      D  , , �j  0/ �j  0� �   0� �   0/ �j  0/      D  , , ��  0/ ��  0� �N  0� �N  0/ ��  0/      D  , , �  0/ �  0� ��  0� ��  0/ �  0/      D  , , �  -� �  .E ��  .E ��  -� �  -�      D  , , �j  -� �j  .E �   .E �   -� �j  -�      D  , , ��  .� ��  /� �d  /� �d  .� ��  .�      D  , , �  .� �  /� ��  /� ��  .� �  .�      D  , , �j  .� �j  /� �   /� �   .� �j  .�      D  , , �H  1o �H  2 ��  2 ��  1o �H  1o      D  , , ��  2� ��  3E ��  3E ��  2� ��  2�      D  , , ��  0/ ��  0� ��  0� ��  0/ ��  0/      D  , , �H  0/ �H  0� ��  0� ��  0/ �H  0/      D  , , ��  ,o ��  - ��  - ��  ,o ��  ,o      D  , , ��  0/ ��  0� �,  0� �,  0/ ��  0/      D  , , ��  0/ ��  0� �z  0� �z  0/ ��  0/      D  , , �2  0/ �2  0� ��  0� ��  0/ �2  0/      D  , , �H  ,o �H  - ��  - ��  ,o �H  ,o      D  , , ��  ,o ��  - �,  - �,  ,o ��  ,o      D  , , ��  ,o ��  - �z  - �z  ,o ��  ,o      D  , , �2  ,o �2  - ��  - ��  ,o �2  ,o      D  , , ��  1o ��  2 �,  2 �,  1o ��  1o      D  , , ��  -� ��  .E ��  .E ��  -� ��  -�      D  , , �H  -� �H  .E ��  .E ��  -� �H  -�      D  , , �H  2� �H  3E ��  3E ��  2� �H  2�      D  , , ��  2� ��  3E �,  3E �,  2� ��  2�      D  , , ��  2� ��  3E �z  3E �z  2� ��  2�      D  , , �2  2� �2  3E ��  3E ��  2� �2  2�      D  , , ��  -� ��  .E �,  .E �,  -� ��  -�      D  , , ��  1o ��  2 ��  2 ��  1o ��  1o      D  , , ��  .� ��  /� ��  /� ��  .� ��  .�      D  , , �H  .� �H  /� ��  /� ��  .� �H  .�      D  , , ��  .� ��  /� �,  /� �,  .� ��  .�      D  , , ��  .� ��  /� �z  /� �z  .� ��  .�      D  , , �2  .� �2  /� ��  /� ��  .� �2  .�      D  , , ��  -� ��  .E �z  .E �z  -� ��  -�      D  , , �2  -� �2  .E ��  .E ��  -� �2  -�      D  , , ��  1o ��  2 �z  2 �z  1o ��  1o      D  , , �2  1o �2  2 ��  2 ��  1o �2  1o      D  , , ��  &� ��  '[ �S  '[ �S  &� ��  &�      D  , , �  &� �  '[ ��  '[ ��  &� �  &�      D  , , �Y  &� �Y  '[ ��  '[ ��  &� �Y  &�      D  , , ��  )� ��  *� �,  *� �,  )� ��  )�      D  , , ��  )� ��  *� �z  *� �z  )� ��  )�      D  , , �2  )� �2  *� ��  *� ��  )� �2  )�      D  , , ��  +/ ��  +� �,  +� �,  +/ ��  +/      D  , , ��  +/ ��  +� �z  +� �z  +/ ��  +/      D  , , �2  +/ �2  +� ��  +� ��  +/ �2  +/      D  , , �!  %� �!  & ��  & ��  %� �!  %�      D  , , �o  %� �o  & �  & �  %� �o  %�      D  , , ��  %� ��  & �S  & �S  %� ��  %�      D  , , �  %� �  & ��  & ��  %� �  %�      D  , , �Y  %� �Y  & ��  & ��  %� �Y  %�      D  , , ��  +/ ��  +� ��  +� ��  +/ ��  +/      D  , , �H  +/ �H  +� ��  +� ��  +/ �H  +/      D  , , ��  )� ��  *� ��  *� ��  )� ��  )�      D  , , �H  )� �H  *� ��  *� ��  )� �H  )�      D  , , �!  &� �!  '[ ��  '[ ��  &� �!  &�      D  , , �o  &� �o  '[ �  '[ �  &� �o  &�      D  , , ��  +/ ��  +� �d  +� �d  +/ ��  +/      D  , , �  +/ �  +� ��  +� ��  +/ �  +/      D  , , ��  )� ��  *� �d  *� �d  )� ��  )�      D  , , �  )� �  *� ��  *� ��  )� �  )�      D  , , �j  )� �j  *� �   *� �   )� �j  )�      D  , , ��  )� ��  *� �N  *� �N  )� ��  )�      D  , , �  )� �  *� ��  *� ��  )� �  )�      D  , , �j  +/ �j  +� �   +� �   +/ �j  +/      D  , , ��  &� ��  '[ �=  '[ �=  &� ��  &�      D  , , ��  %� ��  & �=  & �=  %� ��  %�      D  , , ��  %� ��  & ��  & ��  %� ��  %�      D  , , �C  %� �C  & ��  & ��  %� �C  %�      D  , , ��  %� ��  & �'  & �'  %� ��  %�      D  , , ��  %� ��  & �u  & �u  %� ��  %�      D  , , ��  &� ��  '[ ��  '[ ��  &� ��  &�      D  , , �C  &� �C  '[ ��  '[ ��  &� �C  &�      D  , , ��  &� ��  '[ �'  '[ �'  &� ��  &�      D  , , ��  &� ��  '[ �u  '[ �u  &� ��  &�      D  , , ��  +/ ��  +� �N  +� �N  +/ ��  +/      D  , , �  +/ �  +� ��  +� ��  +/ �  +/      D  , , ��  "[ ��  "� ��  "� ��  "[ ��  "[      D  , , �H  "[ �H  "� ��  "� ��  "[ �H  "[      D  , , ��  "[ ��  "� �,  "� �,  "[ ��  "[      D  , , ��  "[ ��  "� �z  "� �z  "[ ��  "[      D  , , �2  "[ �2  "� ��  "� ��  "[ �2  "[      D  , , ��  "[ ��  "� �  "� �  "[ ��  "[      D  , , ��  "[ ��  "� �d  "� �d  "[ ��  "[      D  , , �  "[ �  "� ��  "� ��  "[ �  "[      D  , , �j  "[ �j  "� �   "� �   "[ �j  "[      D  , , ��  "[ ��  "� �N  "� �N  "[ ��  "[      D  , , �  "[ �  "� ��  "� ��  "[ �  "[      D  , , ��  ! ��  !� ��  !� ��  ! ��  !      D  , , �H  ! �H  !� ��  !� ��  ! �H  !      D  , , ��  ! ��  !� �,  !� �,  ! ��  !      D  , , ��  ! ��  !� �z  !� �z  ! ��  !      D  , , �2  ! �2  !� ��  !� ��  ! �2  !      D  , , ��  ! ��  !� �  !� �  ! ��  !      D  , , ��  ! ��  !� �d  !� �d  ! ��  !      D  , , �  ! �  !� ��  !� ��  ! �  !      D  , , �j  ! �j  !� �   !� �   ! �j  !      D  , , ��  ! ��  !� �N  !� �N  ! ��  !      D  , , �  ! �  !� ��  !� ��  ! �  !      D  , , ��  � ��   q ��   q ��  � ��  �      D  , , �H  � �H   q ��   q ��  � �H  �      D  , , ��  � ��   q �,   q �,  � ��  �      D  , , ��  � ��   q �z   q �z  � ��  �      D  , , �2  � �2   q ��   q ��  � �2  �      D  , , ��  � ��   q �   q �  � ��  �      D  , , ��  � ��   q �d   q �d  � ��  �      D  , , �  � �   q ��   q ��  � �  �      D  , , �j  � �j   q �    q �   � �j  �      D  , , ��  � ��   q �N   q �N  � ��  �      D  , , �  � �   q ��   q ��  � �  �      D  , , ��  � ��  1 ��  1 ��  � ��  �      D  , , �H  � �H  1 ��  1 ��  � �H  �      D  , , ��  � ��  1 �,  1 �,  � ��  �      D  , , ��  � ��  1 �z  1 �z  � ��  �      D  , , �2  � �2  1 ��  1 ��  � �2  �      D  , , ��  � ��  1 �  1 �  � ��  �      D  , , ��  � ��  1 �d  1 �d  � ��  �      D  , , �  � �  1 ��  1 ��  � �  �      D  , , �j  � �j  1 �   1 �   � �j  �      D  , , ��  � ��  1 �N  1 �N  � ��  �      D  , , �  � �  1 ��  1 ��  � �  �      D  , , ��  [ ��  � ��  � ��  [ ��  [      D  , , �H  [ �H  � ��  � ��  [ �H  [      D  , , ��  [ ��  � �,  � �,  [ ��  [      D  , , ��  [ ��  � �z  � �z  [ ��  [      D  , , �2  [ �2  � ��  � ��  [ �2  [      D  , , ��  [ ��  � �  � �  [ ��  [      D  , , ��  [ ��  � �d  � �d  [ ��  [      D  , , �  [ �  � ��  � ��  [ �  [      D  , , �j  [ �j  � �   � �   [ �j  [      D  , , ��  [ ��  � �N  � �N  [ ��  [      D  , , �  [ �  � ��  � ��  [ �  [      D  , , ��   ��  � ��  � ��   ��        D  , , �H   �H  � ��  � ��   �H        D  , , ��   ��  � �,  � �,   ��        D  , , ��   ��  � �z  � �z   ��        D  , , �2   �2  � ��  � ��   �2        D  , , ��   ��  � �  � �   ��        D  , , ��   ��  � �d  � �d   ��        D  , , �   �  � ��  � ��   �        D  , , �j   �j  � �   � �    �j        D  , , ��   ��  � �N  � �N   ��        D  , , �   �  � ��  � ��   �        D  , , ��  � ��  q ��  q ��  � ��  �      D  , , �H  � �H  q ��  q ��  � �H  �      D  , , ��  � ��  q �,  q �,  � ��  �      D  , , ��  � ��  q �z  q �z  � ��  �      D  , , �2  � �2  q ��  q ��  � �2  �      D  , , ��  � ��  q �  q �  � ��  �      D  , , ��  � ��  q �d  q �d  � ��  �      D  , , �  � �  q ��  q ��  � �  �      D  , , �j  � �j  q �   q �   � �j  �      D  , , ��  � ��  q �N  q �N  � ��  �      D  , , �  � �  q ��  q ��  � �  �      D  , , ��  � ��  1 ��  1 ��  � ��  �      D  , , �H  � �H  1 ��  1 ��  � �H  �      D  , , ��  � ��  1 �,  1 �,  � ��  �      D  , , ��  � ��  1 �z  1 �z  � ��  �      D  , , �2  � �2  1 ��  1 ��  � �2  �      D  , , ��  � ��  1 �  1 �  � ��  �      D  , , ��  � ��  1 �d  1 �d  � ��  �      D  , , �  � �  1 ��  1 ��  � �  �      D  , , �j  � �j  1 �   1 �   � �j  �      D  , , ��  � ��  1 �N  1 �N  � ��  �      D  , , �  � �  1 ��  1 ��  � �  �      D  , , �T  ! �T  !� ��  !� ��  ! �T  !      D  , , Ţ  ! Ţ  !� �8  !� �8  ! Ţ  !      D  , , ��  ! ��  !� Ȇ  !� Ȇ  ! ��  !      D  , , �>  ! �>  !� ��  !� ��  ! �>  !      D  , , �T  � �T  1 ��  1 ��  � �T  �      D  , , Ţ  � Ţ  1 �8  1 �8  � Ţ  �      D  , , ��  � ��  1 Ȇ  1 Ȇ  � ��  �      D  , , �>  � �>  1 ��  1 ��  � �>  �      D  , , �T   �T  � ��  � ��   �T        D  , , Ţ   Ţ  � �8  � �8   Ţ        D  , , ��   ��  � Ȇ  � Ȇ   ��        D  , , �>   �>  � ��  � ��   �>        D  , , ̌   ̌  � �"  � �"   ̌        D  , , ��   ��  � �p  � �p   ��        D  , , ̌  � ̌  1 �"  1 �"  � ̌  �      D  , , ��  � ��  1 �p  1 �p  � ��  �      D  , , ̌  ! ̌  !� �"  !� �"  ! ̌  !      D  , , �T  � �T   q ��   q ��  � �T  �      D  , , Ţ  � Ţ   q �8   q �8  � Ţ  �      D  , , ��  � ��   q Ȇ   q Ȇ  � ��  �      D  , , �>  � �>   q ��   q ��  � �>  �      D  , , ̌  � ̌   q �"   q �"  � ̌  �      D  , , ��  � ��   q �p   q �p  � ��  �      D  , , ��  ! ��  !� �p  !� �p  ! ��  !      D  , , ��  "[ ��  "� �p  "� �p  "[ ��  "[      D  , , �T  � �T  q ��  q ��  � �T  �      D  , , Ţ  � Ţ  q �8  q �8  � Ţ  �      D  , , ��  � ��  q Ȇ  q Ȇ  � ��  �      D  , , �>  � �>  q ��  q ��  � �>  �      D  , , ̌  � ̌  q �"  q �"  � ̌  �      D  , , ��  � ��  q �p  q �p  � ��  �      D  , , �T  "[ �T  "� ��  "� ��  "[ �T  "[      D  , , Ţ  "[ Ţ  "� �8  "� �8  "[ Ţ  "[      D  , , �T  [ �T  � ��  � ��  [ �T  [      D  , , Ţ  [ Ţ  � �8  � �8  [ Ţ  [      D  , , ��  [ ��  � Ȇ  � Ȇ  [ ��  [      D  , , �>  [ �>  � ��  � ��  [ �>  [      D  , , ̌  [ ̌  � �"  � �"  [ ̌  [      D  , , ��  [ ��  � �p  � �p  [ ��  [      D  , , ��  "[ ��  "� Ȇ  "� Ȇ  "[ ��  "[      D  , , �>  "[ �>  "� ��  "� ��  "[ �>  "[      D  , , ̌  "[ ̌  "� �"  "� �"  "[ ̌  "[      D  , , �T  � �T  1 ��  1 ��  � �T  �      D  , , Ţ  � Ţ  1 �8  1 �8  � Ţ  �      D  , , ��  � ��  1 Ȇ  1 Ȇ  � ��  �      D  , , �>  � �>  1 ��  1 ��  � �>  �      D  , , ̌  � ̌  1 �"  1 �"  � ̌  �      D  , , ��  � ��  1 �p  1 �p  � ��  �      D  , , �<  .� �<  /� ��  /� ��  .� �<  .�      D  , , ��  .� ��  /� �   /� �   .� ��  .�      D  , , ��  .� ��  /� �n  /� �n  .� ��  .�      D  , , �&  .� �&  /� ��  /� ��  .� �&  .�      D  , , �t  .� �t  /� �
  /� �
  .� �t  .�      D  , , ��  .� ��  /� �X  /� �X  .� ��  .�      D  , , �  .� �  /� ��  /� ��  .� �  .�      D  , , �^  .� �^  /� ��  /� ��  .� �^  .�      D  , , �<  +/ �<  +� ��  +� ��  +/ �<  +/      D  , , ��  +/ ��  +� �   +� �   +/ ��  +/      D  , , ��  +/ ��  +� �n  +� �n  +/ ��  +/      D  , , �&  +/ �&  +� ��  +� ��  +/ �&  +/      D  , , �t  +/ �t  +� �
  +� �
  +/ �t  +/      D  , , ��  +/ ��  +� �X  +� �X  +/ ��  +/      D  , , �  +/ �  +� ��  +� ��  +/ �  +/      D  , , �^  +/ �^  +� ��  +� ��  +/ �^  +/      D  , , ��  +/ ��  +� �B  +� �B  +/ ��  +/      D  , , ��  .� ��  /� �B  /� �B  .� ��  .�      D  , , ��  2� ��  3E �B  3E �B  2� ��  2�      D  , , �<  0/ �<  0� ��  0� ��  0/ �<  0/      D  , , ��  0/ ��  0� �   0� �   0/ ��  0/      D  , , ��  0/ ��  0� �n  0� �n  0/ ��  0/      D  , , �<  )� �<  *� ��  *� ��  )� �<  )�      D  , , ��  )� ��  *� �   *� �   )� ��  )�      D  , , ��  )� ��  *� �n  *� �n  )� ��  )�      D  , , �&  )� �&  *� ��  *� ��  )� �&  )�      D  , , �t  )� �t  *� �
  *� �
  )� �t  )�      D  , , ��  )� ��  *� �X  *� �X  )� ��  )�      D  , , �  )� �  *� ��  *� ��  )� �  )�      D  , , �^  )� �^  *� ��  *� ��  )� �^  )�      D  , , ��  )� ��  *� �B  *� �B  )� ��  )�      D  , , �&  0/ �&  0� ��  0� ��  0/ �&  0/      D  , , �<  -� �<  .E ��  .E ��  -� �<  -�      D  , , ��  -� ��  .E �   .E �   -� ��  -�      D  , , ��  -� ��  .E �n  .E �n  -� ��  -�      D  , , �&  -� �&  .E ��  .E ��  -� �&  -�      D  , , �t  -� �t  .E �
  .E �
  -� �t  -�      D  , , ��  -� ��  .E �X  .E �X  -� ��  -�      D  , , �  -� �  .E ��  .E ��  -� �  -�      D  , , �^  -� �^  .E ��  .E ��  -� �^  -�      D  , , ��  -� ��  .E �B  .E �B  -� ��  -�      D  , , �t  0/ �t  0� �
  0� �
  0/ �t  0/      D  , , ��  0/ ��  0� �X  0� �X  0/ ��  0/      D  , , �  0/ �  0� ��  0� ��  0/ �  0/      D  , , �c  &� �c  '[ ��  '[ ��  &� �c  &�      D  , , ��  &� ��  '[ �G  '[ �G  &� ��  &�      D  , , ��  &� ��  '[ ��  '[ ��  &� ��  &�      D  , , �M  &� �M  '[ ��  '[ ��  &� �M  &�      D  , , ��  &� ��  '[ �1  '[ �1  &� ��  &�      D  , , ��  &� ��  '[ �  '[ �  &� ��  &�      D  , , �7  &� �7  '[ ��  '[ ��  &� �7  &�      D  , , ��  &� ��  '[ �  '[ �  &� ��  &�      D  , , ��  &� ��  '[ �i  '[ �i  &� ��  &�      D  , , �^  0/ �^  0� ��  0� ��  0/ �^  0/      D  , , ��  0/ ��  0� �B  0� �B  0/ ��  0/      D  , , �<  1o �<  2 ��  2 ��  1o �<  1o      D  , , ��  1o ��  2 �   2 �   1o ��  1o      D  , , ��  1o ��  2 �n  2 �n  1o ��  1o      D  , , �&  1o �&  2 ��  2 ��  1o �&  1o      D  , , �t  1o �t  2 �
  2 �
  1o �t  1o      D  , , ��  1o ��  2 �X  2 �X  1o ��  1o      D  , , �  1o �  2 ��  2 ��  1o �  1o      D  , , �^  1o �^  2 ��  2 ��  1o �^  1o      D  , , ��  1o ��  2 �B  2 �B  1o ��  1o      D  , , �<  2� �<  3E ��  3E ��  2� �<  2�      D  , , ��  2� ��  3E �   3E �   2� ��  2�      D  , , ��  2� ��  3E �n  3E �n  2� ��  2�      D  , , �c  %� �c  & ��  & ��  %� �c  %�      D  , , ��  %� ��  & �G  & �G  %� ��  %�      D  , , ��  %� ��  & ��  & ��  %� ��  %�      D  , , �M  %� �M  & ��  & ��  %� �M  %�      D  , , ��  %� ��  & �1  & �1  %� ��  %�      D  , , ��  %� ��  & �  & �  %� ��  %�      D  , , �7  %� �7  & ��  & ��  %� �7  %�      D  , , ��  %� ��  & �  & �  %� ��  %�      D  , , ��  %� ��  & �i  & �i  %� ��  %�      D  , , �<  ,o �<  - ��  - ��  ,o �<  ,o      D  , , ��  ,o ��  - �   - �   ,o ��  ,o      D  , , ��  ,o ��  - �n  - �n  ,o ��  ,o      D  , , �&  ,o �&  - ��  - ��  ,o �&  ,o      D  , , �t  ,o �t  - �
  - �
  ,o �t  ,o      D  , , ��  ,o ��  - �X  - �X  ,o ��  ,o      D  , , �  ,o �  - ��  - ��  ,o �  ,o      D  , , �^  ,o �^  - ��  - ��  ,o �^  ,o      D  , , ��  ,o ��  - �B  - �B  ,o ��  ,o      D  , , �&  2� �&  3E ��  3E ��  2� �&  2�      D  , , �t  2� �t  3E �
  3E �
  2� �t  2�      D  , , ��  2� ��  3E �X  3E �X  2� ��  2�      D  , , �  2� �  3E ��  3E ��  2� �  2�      D  , , �^  2� �^  3E ��  3E ��  2� �^  2�      D  , , ~S  -� ~S  .E ~�  .E ~�  -� ~S  -�      D  , , y�  1o y�  2 zM  2 zM  1o y�  1o      D  , , |  1o |  2 |�  2 |�  1o |  1o      D  , , ~S  1o ~S  2 ~�  2 ~�  1o ~S  1o      D  , , wi  0/ wi  0� w�  0� w�  0/ wi  0/      D  , , y�  0/ y�  0� zM  0� zM  0/ y�  0/      D  , , |  0/ |  0� |�  0� |�  0/ |  0/      D  , , ~S  0/ ~S  0� ~�  0� ~�  0/ ~S  0/      D  , , wi  ,o wi  - w�  - w�  ,o wi  ,o      D  , , y�  ,o y�  - zM  - zM  ,o y�  ,o      D  , , x�  %� x�  & y&  & y&  %� x�  %�      D  , , z�  %� z�  & {t  & {t  %� z�  %�      D  , , },  %� },  & }�  & }�  %� },  %�      D  , , ~S  .� ~S  /� ~�  /� ~�  .� ~S  .�      D  , , wi  +/ wi  +� w�  +� w�  +/ wi  +/      D  , , y�  +/ y�  +� zM  +� zM  +/ y�  +/      D  , , wi  )� wi  *� w�  *� w�  )� wi  )�      D  , , y�  )� y�  *� zM  *� zM  )� y�  )�      D  , , x�  &� x�  '[ y&  '[ y&  &� x�  &�      D  , , z�  &� z�  '[ {t  '[ {t  &� z�  &�      D  , , },  &� },  '[ }�  '[ }�  &� },  &�      D  , , |  )� |  *� |�  *� |�  )� |  )�      D  , , |  ,o |  - |�  - |�  ,o |  ,o      D  , , ~S  ,o ~S  - ~�  - ~�  ,o ~S  ,o      D  , , ~S  )� ~S  *� ~�  *� ~�  )� ~S  )�      D  , , |  +/ |  +� |�  +� |�  +/ |  +/      D  , , ~S  +/ ~S  +� ~�  +� ~�  +/ ~S  +/      D  , , wi  .� wi  /� w�  /� w�  .� wi  .�      D  , , y�  .� y�  /� zM  /� zM  .� y�  .�      D  , , |  .� |  /� |�  /� |�  .� |  .�      D  , , wi  2� wi  3E w�  3E w�  2� wi  2�      D  , , y�  2� y�  3E zM  3E zM  2� y�  2�      D  , , |  2� |  3E |�  3E |�  2� |  2�      D  , , ~S  2� ~S  3E ~�  3E ~�  2� ~S  2�      D  , , wi  1o wi  2 w�  2 w�  1o wi  1o      D  , , wi  -� wi  .E w�  .E w�  -� wi  -�      D  , , y�  -� y�  .E zM  .E zM  -� y�  -�      D  , , |  -� |  .E |�  .E |�  -� |  -�      D  , , ~S   ~S  � ~�  � ~�   ~S        D  , , ~S  � ~S   q ~�   q ~�  � ~S  �      D  , , y�  ! y�  !� zM  !� zM  ! y�  !      D  , , wi  � wi  1 w�  1 w�  � wi  �      D  , , y�  � y�  1 zM  1 zM  � y�  �      D  , , |  � |  1 |�  1 |�  � |  �      D  , , ~S  � ~S  1 ~�  1 ~�  � ~S  �      D  , , |  ! |  !� |�  !� |�  ! |  !      D  , , ~S  ! ~S  !� ~�  !� ~�  ! ~S  !      D  , , wi  ! wi  !� w�  !� w�  ! wi  !      D  , , wi  � wi   q w�   q w�  � wi  �      D  , , y�  � y�   q zM   q zM  � y�  �      D  , , wi  [ wi  � w�  � w�  [ wi  [      D  , , y�  [ y�  � zM  � zM  [ y�  [      D  , , |  [ |  � |�  � |�  [ |  [      D  , , wi  � wi  1 w�  1 w�  � wi  �      D  , , y�  � y�  1 zM  1 zM  � y�  �      D  , , |  � |  1 |�  1 |�  � |  �      D  , , ~S  � ~S  1 ~�  1 ~�  � ~S  �      D  , , ~S  [ ~S  � ~�  � ~�  [ ~S  [      D  , , |  � |   q |�   q |�  � |  �      D  , , wi   wi  � w�  � w�   wi        D  , , wi  � wi  q w�  q w�  � wi  �      D  , , y�  � y�  q zM  q zM  � y�  �      D  , , |  � |  q |�  q |�  � |  �      D  , , ~S  � ~S  q ~�  q ~�  � ~S  �      D  , , y�   y�  � zM  � zM   y�        D  , , |   |  � |�  � |�   |        D  , , wi  "[ wi  "� w�  "� w�  "[ wi  "[      D  , , y�  "[ y�  "� zM  "� zM  "[ y�  "[      D  , , |  "[ |  "� |�  "� |�  "[ |  "[      D  , , ~S  "[ ~S  "� ~�  "� ~�  "[ ~S  "[      D  , , ��  ! ��  !� �   !� �   ! ��  !      D  , , �<  � �<   q ��   q ��  � �<  �      D  , , ��  � ��   q �    q �   � ��  �      D  , , ��  � ��   q �n   q �n  � ��  �      D  , , �&  � �&   q ��   q ��  � �&  �      D  , , �t  � �t   q �
   q �
  � �t  �      D  , , �<  [ �<  � ��  � ��  [ �<  [      D  , , ��  [ ��  � �   � �   [ ��  [      D  , , ��  [ ��  � �n  � �n  [ ��  [      D  , , �&  [ �&  � ��  � ��  [ �&  [      D  , , �t  [ �t  � �
  � �
  [ �t  [      D  , , ��  [ ��  � �X  � �X  [ ��  [      D  , , �  [ �  � ��  � ��  [ �  [      D  , , �^  [ �^  � ��  � ��  [ �^  [      D  , , ��  [ ��  � �B  � �B  [ ��  [      D  , , ��  � ��   q �X   q �X  � ��  �      D  , , �<  � �<  q ��  q ��  � �<  �      D  , , ��  � ��  q �   q �   � ��  �      D  , , ��  � ��  q �n  q �n  � ��  �      D  , , �&  � �&  q ��  q ��  � �&  �      D  , , �t  � �t  q �
  q �
  � �t  �      D  , , ��  � ��  q �X  q �X  � ��  �      D  , , �  � �  q ��  q ��  � �  �      D  , , �^  � �^  q ��  q ��  � �^  �      D  , , ��  � ��  q �B  q �B  � ��  �      D  , , �  � �   q ��   q ��  � �  �      D  , , �<  � �<  1 ��  1 ��  � �<  �      D  , , ��  � ��  1 �   1 �   � ��  �      D  , , ��  � ��  1 �n  1 �n  � ��  �      D  , , �&  � �&  1 ��  1 ��  � �&  �      D  , , �t  � �t  1 �
  1 �
  � �t  �      D  , , ��  � ��  1 �X  1 �X  � ��  �      D  , , �  � �  1 ��  1 ��  � �  �      D  , , �^  � �^  1 ��  1 ��  � �^  �      D  , , ��  � ��  1 �B  1 �B  � ��  �      D  , , �^  � �^   q ��   q ��  � �^  �      D  , , ��  � ��   q �B   q �B  � ��  �      D  , , ��  ! ��  !� �n  !� �n  ! ��  !      D  , , �&  ! �&  !� ��  !� ��  ! �&  !      D  , , �t  ! �t  !� �
  !� �
  ! �t  !      D  , , ��  ! ��  !� �X  !� �X  ! ��  !      D  , , �  ! �  !� ��  !� ��  ! �  !      D  , , �^  ! �^  !� ��  !� ��  ! �^  !      D  , , ��  ! ��  !� �B  !� �B  ! ��  !      D  , , ��  "[ ��  "� �X  "� �X  "[ ��  "[      D  , , �<   �<  � ��  � ��   �<        D  , , �<  � �<  1 ��  1 ��  � �<  �      D  , , ��  � ��  1 �   1 �   � ��  �      D  , , ��  � ��  1 �n  1 �n  � ��  �      D  , , �&  � �&  1 ��  1 ��  � �&  �      D  , , �t  � �t  1 �
  1 �
  � �t  �      D  , , ��  � ��  1 �X  1 �X  � ��  �      D  , , �  � �  1 ��  1 ��  � �  �      D  , , �^  � �^  1 ��  1 ��  � �^  �      D  , , ��  � ��  1 �B  1 �B  � ��  �      D  , , ��   ��  � �   � �    ��        D  , , ��   ��  � �n  � �n   ��        D  , , �&   �&  � ��  � ��   �&        D  , , �t   �t  � �
  � �
   �t        D  , , ��   ��  � �X  � �X   ��        D  , , �   �  � ��  � ��   �        D  , , �^   �^  � ��  � ��   �^        D  , , ��   ��  � �B  � �B   ��        D  , , �  "[ �  "� ��  "� ��  "[ �  "[      D  , , �^  "[ �^  "� ��  "� ��  "[ �^  "[      D  , , ��  "[ ��  "� �B  "� �B  "[ ��  "[      D  , , �t  "[ �t  "� �
  "� �
  "[ �t  "[      D  , , �<  ! �<  !� ��  !� ��  ! �<  !      D  , , �<  "[ �<  "� ��  "� ��  "[ �<  "[      D  , , ��  "[ ��  "� �   "� �   "[ ��  "[      D  , , ��  "[ ��  "� �n  "� �n  "[ ��  "[      D  , , �&  "[ �&  "� ��  "� ��  "[ �&  "[      D  , , D�  2� D�  3E EK  3E EK  2� D�  2�      D  , , D�  -� D�  .E EK  .E EK  -� D�  -�      D  , , D�  "[ D�  "� EK  "� EK  "[ D�  "[      D  , , D�  0/ D�  0� EK  0� EK  0/ D�  0/      D  , , D�  ! D�  !� EK  !� EK  ! D�  !      D  , , D�  ,o D�  - EK  - EK  ,o D�  ,o      D  , , D�  � D�   q EK   q EK  � D�  �      D  , , D�  1o D�  2 EK  2 EK  1o D�  1o      D  , , D�  � D�  1 EK  1 EK  � D�  �      D  , , D�  +/ D�  +� EK  +� EK  +/ D�  +/      D  , , D�  [ D�  � EK  � EK  [ D�  [      D  , , D�  .� D�  /� EK  /� EK  .� D�  .�      D  , , D�   D�  � EK  � EK   D�        D  , , D�  )� D�  *� EK  *� EK  )� D�  )�      D  , , D�  � D�  q EK  q EK  � D�  �      D  , , D�  � D�  1 EK  1 EK  � D�  �      D  , , ^  2� ^  3E ^�  3E ^�  2� ^  2�      D  , , ^  -� ^  .E ^�  .E ^�  -� ^  -�      D  , , ^  "[ ^  "� ^�  "� ^�  "[ ^  "[      D  , , ^  0/ ^  0� ^�  0� ^�  0/ ^  0/      D  , , ^  ! ^  !� ^�  !� ^�  ! ^  !      D  , , ^  ,o ^  - ^�  - ^�  ,o ^  ,o      D  , , ^  � ^   q ^�   q ^�  � ^  �      D  , , ^  � ^  1 ^�  1 ^�  � ^  �      D  , , ^  +/ ^  +� ^�  +� ^�  +/ ^  +/      D  , , ^  [ ^  � ^�  � ^�  [ ^  [      D  , , ^  1o ^  2 ^�  2 ^�  1o ^  1o      D  , , ^   ^  � ^�  � ^�   ^        D  , , ^  )� ^  *� ^�  *� ^�  )� ^  )�      D  , , ^  � ^  q ^�  q ^�  � ^  �      D  , , ^  .� ^  /� ^�  /� ^�  .� ^  .�      D  , , ^  � ^  1 ^�  1 ^�  � ^  �      D  , , j�  &� j�  '[ kR  '[ kR  &� j�  &�      D  , , j�  %� j�  & kR  & kR  %� j�  %�      D  , , p  -� p  .E q  .E q  -� p  -�      D  , , r�  -� r�  .E sc  .E sc  -� r�  -�      D  , , u  -� u  .E u�  .E u�  -� u  -�      D  , , k�  2� k�  3E ly  3E ly  2� k�  2�      D  , , k�  -� k�  .E ly  .E ly  -� k�  -�      D  , , k�  ,o k�  - ly  - ly  ,o k�  ,o      D  , , n1  ,o n1  - n�  - n�  ,o n1  ,o      D  , , p  ,o p  - q  - q  ,o p  ,o      D  , , r�  ,o r�  - sc  - sc  ,o r�  ,o      D  , , u  ,o u  - u�  - u�  ,o u  ,o      D  , , k�  0/ k�  0� ly  0� ly  0/ k�  0/      D  , , n1  0/ n1  0� n�  0� n�  0/ n1  0/      D  , , p  0/ p  0� q  0� q  0/ p  0/      D  , , r�  0/ r�  0� sc  0� sc  0/ r�  0/      D  , , u  0/ u  0� u�  0� u�  0/ u  0/      D  , , n1  2� n1  3E n�  3E n�  2� n1  2�      D  , , p  2� p  3E q  3E q  2� p  2�      D  , , n1  -� n1  .E n�  .E n�  -� n1  -�      D  , , k�  .� k�  /� ly  /� ly  .� k�  .�      D  , , n1  .� n1  /� n�  /� n�  .� n1  .�      D  , , p  .� p  /� q  /� q  .� p  .�      D  , , r�  .� r�  /� sc  /� sc  .� r�  .�      D  , , u  .� u  /� u�  /� u�  .� u  .�      D  , , k�  1o k�  2 ly  2 ly  1o k�  1o      D  , , n1  1o n1  2 n�  2 n�  1o n1  1o      D  , , p  1o p  2 q  2 q  1o p  1o      D  , , r�  1o r�  2 sc  2 sc  1o r�  1o      D  , , u  1o u  2 u�  2 u�  1o u  1o      D  , , r�  2� r�  3E sc  3E sc  2� r�  2�      D  , , u  2� u  3E u�  3E u�  2� u  2�      D  , , d�  -� d�  .E e�  .E e�  -� d�  -�      D  , , `]  ,o `]  - `�  - `�  ,o `]  ,o      D  , , b�  ,o b�  - cA  - cA  ,o b�  ,o      D  , , d�  ,o d�  - e�  - e�  ,o d�  ,o      D  , , gG  ,o gG  - g�  - g�  ,o gG  ,o      D  , , i�  ,o i�  - j+  - j+  ,o i�  ,o      D  , , `]  1o `]  2 `�  2 `�  1o `]  1o      D  , , b�  1o b�  2 cA  2 cA  1o b�  1o      D  , , d�  1o d�  2 e�  2 e�  1o d�  1o      D  , , gG  1o gG  2 g�  2 g�  1o gG  1o      D  , , `]  -� `]  .E `�  .E `�  -� `]  -�      D  , , `]  .� `]  /� `�  /� `�  .� `]  .�      D  , , b�  .� b�  /� cA  /� cA  .� b�  .�      D  , , d�  .� d�  /� e�  /� e�  .� d�  .�      D  , , gG  .� gG  /� g�  /� g�  .� gG  .�      D  , , i�  .� i�  /� j+  /� j+  .� i�  .�      D  , , gG  -� gG  .E g�  .E g�  -� gG  -�      D  , , `]  2� `]  3E `�  3E `�  2� `]  2�      D  , , b�  2� b�  3E cA  3E cA  2� b�  2�      D  , , d�  2� d�  3E e�  3E e�  2� d�  2�      D  , , gG  2� gG  3E g�  3E g�  2� gG  2�      D  , , i�  1o i�  2 j+  2 j+  1o i�  1o      D  , , `]  0/ `]  0� `�  0� `�  0/ `]  0/      D  , , b�  0/ b�  0� cA  0� cA  0/ b�  0/      D  , , d�  0/ d�  0� e�  0� e�  0/ d�  0/      D  , , gG  0/ gG  0� g�  0� g�  0/ gG  0/      D  , , i�  0/ i�  0� j+  0� j+  0/ i�  0/      D  , , i�  2� i�  3E j+  3E j+  2� i�  2�      D  , , i�  -� i�  .E j+  .E j+  -� i�  -�      D  , , b�  -� b�  .E cA  .E cA  -� b�  -�      D  , , b�  +/ b�  +� cA  +� cA  +/ b�  +/      D  , , d�  +/ d�  +� e�  +� e�  +/ d�  +/      D  , , gG  +/ gG  +� g�  +� g�  +/ gG  +/      D  , , i�  +/ i�  +� j+  +� j+  +/ i�  +/      D  , , hn  %� hn  & i  & i  %� hn  %�      D  , , c�  %� c�  & dh  & dh  %� c�  %�      D  , , f   %� f   & f�  & f�  %� f   %�      D  , , _6  %� _6  & _�  & _�  %� _6  %�      D  , , `]  )� `]  *� `�  *� `�  )� `]  )�      D  , , b�  )� b�  *� cA  *� cA  )� b�  )�      D  , , d�  )� d�  *� e�  *� e�  )� d�  )�      D  , , gG  )� gG  *� g�  *� g�  )� gG  )�      D  , , i�  )� i�  *� j+  *� j+  )� i�  )�      D  , , hn  &� hn  '[ i  '[ i  &� hn  &�      D  , , f   &� f   '[ f�  '[ f�  &� f   &�      D  , , a�  %� a�  & b  & b  %� a�  %�      D  , , `]  +/ `]  +� `�  +� `�  +/ `]  +/      D  , , _6  &� _6  '[ _�  '[ _�  &� _6  &�      D  , , a�  &� a�  '[ b  '[ b  &� a�  &�      D  , , c�  &� c�  '[ dh  '[ dh  &� c�  &�      D  , , m
  %� m
  & m�  & m�  %� m
  %�      D  , , s�  &� s�  '[ t�  '[ t�  &� s�  &�      D  , , oX  &� oX  '[ o�  '[ o�  &� oX  &�      D  , , vB  &� vB  '[ v�  '[ v�  &� vB  &�      D  , , s�  %� s�  & t�  & t�  %� s�  %�      D  , , vB  %� vB  & v�  & v�  %� vB  %�      D  , , m
  &� m
  '[ m�  '[ m�  &� m
  &�      D  , , q�  &� q�  '[ r<  '[ r<  &� q�  &�      D  , , k�  +/ k�  +� ly  +� ly  +/ k�  +/      D  , , n1  +/ n1  +� n�  +� n�  +/ n1  +/      D  , , p  +/ p  +� q  +� q  +/ p  +/      D  , , k�  )� k�  *� ly  *� ly  )� k�  )�      D  , , r�  +/ r�  +� sc  +� sc  +/ r�  +/      D  , , n1  )� n1  *� n�  *� n�  )� n1  )�      D  , , p  )� p  *� q  *� q  )� p  )�      D  , , r�  )� r�  *� sc  *� sc  )� r�  )�      D  , , u  )� u  *� u�  *� u�  )� u  )�      D  , , u  +/ u  +� u�  +� u�  +/ u  +/      D  , , oX  %� oX  & o�  & o�  %� oX  %�      D  , , q�  %� q�  & r<  & r<  %� q�  %�      D  , , Qb  %� Qb  & Q�  & Q�  %� Qb  %�      D  , , Qb  &� Qb  '[ Q�  '[ Q�  &� Qb  &�      D  , , T�  -� T�  .E Um  .E Um  -� T�  -�      D  , , W%  -� W%  .E W�  .E W�  -� W%  -�      D  , , Ys  -� Ys  .E Z	  .E Z	  -� Ys  -�      D  , , [�  -� [�  .E \W  .E \W  -� [�  -�      D  , , R�  ,o R�  - S  - S  ,o R�  ,o      D  , , R�  1o R�  2 S  2 S  1o R�  1o      D  , , T�  1o T�  2 Um  2 Um  1o T�  1o      D  , , W%  1o W%  2 W�  2 W�  1o W%  1o      D  , , Ys  1o Ys  2 Z	  2 Z	  1o Ys  1o      D  , , [�  1o [�  2 \W  2 \W  1o [�  1o      D  , , T�  ,o T�  - Um  - Um  ,o T�  ,o      D  , , W%  ,o W%  - W�  - W�  ,o W%  ,o      D  , , Ys  ,o Ys  - Z	  - Z	  ,o Ys  ,o      D  , , [�  ,o [�  - \W  - \W  ,o [�  ,o      D  , , R�  .� R�  /� S  /� S  .� R�  .�      D  , , T�  .� T�  /� Um  /� Um  .� T�  .�      D  , , [�  2� [�  3E \W  3E \W  2� [�  2�      D  , , W%  2� W%  3E W�  3E W�  2� W%  2�      D  , , Ys  2� Ys  3E Z	  3E Z	  2� Ys  2�      D  , , R�  2� R�  3E S  3E S  2� R�  2�      D  , , Ys  0/ Ys  0� Z	  0� Z	  0/ Ys  0/      D  , , W%  .� W%  /� W�  /� W�  .� W%  .�      D  , , Ys  .� Ys  /� Z	  /� Z	  .� Ys  .�      D  , , [�  .� [�  /� \W  /� \W  .� [�  .�      D  , , R�  -� R�  .E S  .E S  -� R�  -�      D  , , R�  0/ R�  0� S  0� S  0/ R�  0/      D  , , T�  0/ T�  0� Um  0� Um  0/ T�  0/      D  , , W%  0/ W%  0� W�  0� W�  0/ W%  0/      D  , , T�  2� T�  3E Um  3E Um  2� T�  2�      D  , , [�  0/ [�  0� \W  0� \W  0/ [�  0/      D  , , G  ,o G  - G�  - G�  ,o G  ,o      D  , , IQ  ,o IQ  - I�  - I�  ,o IQ  ,o      D  , , K�  ,o K�  - L5  - L5  ,o K�  ,o      D  , , G  -� G  .E G�  .E G�  -� G  -�      D  , , M�  ,o M�  - N�  - N�  ,o M�  ,o      D  , , K�  2� K�  3E L5  3E L5  2� K�  2�      D  , , G  .� G  /� G�  /� G�  .� G  .�      D  , , IQ  .� IQ  /� I�  /� I�  .� IQ  .�      D  , , K�  .� K�  /� L5  /� L5  .� K�  .�      D  , , IQ  -� IQ  .E I�  .E I�  -� IQ  -�      D  , , K�  -� K�  .E L5  .E L5  -� K�  -�      D  , , M�  -� M�  .E N�  .E N�  -� M�  -�      D  , , P;  -� P;  .E P�  .E P�  -� P;  -�      D  , , M�  .� M�  /� N�  /� N�  .� M�  .�      D  , , G  0/ G  0� G�  0� G�  0/ G  0/      D  , , IQ  0/ IQ  0� I�  0� I�  0/ IQ  0/      D  , , K�  0/ K�  0� L5  0� L5  0/ K�  0/      D  , , M�  0/ M�  0� N�  0� N�  0/ M�  0/      D  , , P;  0/ P;  0� P�  0� P�  0/ P;  0/      D  , , P;  .� P;  /� P�  /� P�  .� P;  .�      D  , , G  1o G  2 G�  2 G�  1o G  1o      D  , , IQ  1o IQ  2 I�  2 I�  1o IQ  1o      D  , , K�  1o K�  2 L5  2 L5  1o K�  1o      D  , , M�  1o M�  2 N�  2 N�  1o M�  1o      D  , , P;  1o P;  2 P�  2 P�  1o P;  1o      D  , , P;  ,o P;  - P�  - P�  ,o P;  ,o      D  , , IQ  2� IQ  3E I�  3E I�  2� IQ  2�      D  , , M�  2� M�  3E N�  3E N�  2� M�  2�      D  , , G  2� G  3E G�  3E G�  2� G  2�      D  , , P;  2� P;  3E P�  3E P�  2� P;  2�      D  , , P;  )� P;  *� P�  *� P�  )� P;  )�      D  , , M�  +/ M�  +� N�  +� N�  +/ M�  +/      D  , , P;  +/ P;  +� P�  +� P�  +/ P;  +/      D  , , G  )� G  *� G�  *� G�  )� G  )�      D  , , IQ  )� IQ  *� I�  *� I�  )� IQ  )�      D  , , E�  %� E�  & Fr  & Fr  %� E�  %�      D  , , K�  )� K�  *� L5  *� L5  )� K�  )�      D  , , H*  %� H*  & H�  & H�  %� H*  %�      D  , , Jx  %� Jx  & K  & K  %� Jx  %�      D  , , L�  %� L�  & M\  & M\  %� L�  %�      D  , , O  %� O  & O�  & O�  %� O  %�      D  , , E�  &� E�  '[ Fr  '[ Fr  &� E�  &�      D  , , H*  &� H*  '[ H�  '[ H�  &� H*  &�      D  , , Jx  &� Jx  '[ K  '[ K  &� Jx  &�      D  , , L�  &� L�  '[ M\  '[ M\  &� L�  &�      D  , , O  &� O  '[ O�  '[ O�  &� O  &�      D  , , M�  )� M�  *� N�  *� N�  )� M�  )�      D  , , G  +/ G  +� G�  +� G�  +/ G  +/      D  , , IQ  +/ IQ  +� I�  +� I�  +/ IQ  +/      D  , , K�  +/ K�  +� L5  +� L5  +/ K�  +/      D  , , S�  %� S�  & TF  & TF  %� S�  %�      D  , , XL  %� XL  & X�  & X�  %� XL  %�      D  , , R�  +/ R�  +� S  +� S  +/ R�  +/      D  , , T�  +/ T�  +� Um  +� Um  +/ T�  +/      D  , , U�  %� U�  & V�  & V�  %� U�  %�      D  , , W%  +/ W%  +� W�  +� W�  +/ W%  +/      D  , , Ys  +/ Ys  +� Z	  +� Z	  +/ Ys  +/      D  , , [�  +/ [�  +� \W  +� \W  +/ [�  +/      D  , , R�  )� R�  *� S  *� S  )� R�  )�      D  , , T�  )� T�  *� Um  *� Um  )� T�  )�      D  , , W%  )� W%  *� W�  *� W�  )� W%  )�      D  , , Ys  )� Ys  *� Z	  *� Z	  )� Ys  )�      D  , , S�  &� S�  '[ TF  '[ TF  &� S�  &�      D  , , U�  &� U�  '[ V�  '[ V�  &� U�  &�      D  , , XL  &� XL  '[ X�  '[ X�  &� XL  &�      D  , , Z�  &� Z�  '[ [0  '[ [0  &� Z�  &�      D  , , \�  &� \�  '[ ]~  '[ ]~  &� \�  &�      D  , , [�  )� [�  *� \W  *� \W  )� [�  )�      D  , , Z�  %� Z�  & [0  & [0  %� Z�  %�      D  , , \�  %� \�  & ]~  & ]~  %� \�  %�      D  , , M�  � M�   q N�   q N�  � M�  �      D  , , P;  � P;   q P�   q P�  � P;  �      D  , , R�  � R�   q S   q S  � R�  �      D  , , T�  � T�   q Um   q Um  � T�  �      D  , , W%  � W%   q W�   q W�  � W%  �      D  , , Ys  � Ys   q Z	   q Z	  � Ys  �      D  , , [�  � [�   q \W   q \W  � [�  �      D  , , K�  "[ K�  "� L5  "� L5  "[ K�  "[      D  , , M�  "[ M�  "� N�  "� N�  "[ M�  "[      D  , , G  ! G  !� G�  !� G�  ! G  !      D  , , IQ  ! IQ  !� I�  !� I�  ! IQ  !      D  , , K�  ! K�  !� L5  !� L5  ! K�  !      D  , , M�  ! M�  !� N�  !� N�  ! M�  !      D  , , P;  ! P;  !� P�  !� P�  ! P;  !      D  , , R�  ! R�  !� S  !� S  ! R�  !      D  , , T�  ! T�  !� Um  !� Um  ! T�  !      D  , , W%  ! W%  !� W�  !� W�  ! W%  !      D  , , G  � G  q G�  q G�  � G  �      D  , , IQ  � IQ  q I�  q I�  � IQ  �      D  , , K�  � K�  q L5  q L5  � K�  �      D  , , M�  � M�  q N�  q N�  � M�  �      D  , , P;  � P;  q P�  q P�  � P;  �      D  , , R�  � R�  q S  q S  � R�  �      D  , , T�  � T�  q Um  q Um  � T�  �      D  , , W%  � W%  q W�  q W�  � W%  �      D  , , Ys  � Ys  q Z	  q Z	  � Ys  �      D  , , [�  � [�  q \W  q \W  � [�  �      D  , , G  [ G  � G�  � G�  [ G  [      D  , , IQ  [ IQ  � I�  � I�  [ IQ  [      D  , , K�  [ K�  � L5  � L5  [ K�  [      D  , , M�  [ M�  � N�  � N�  [ M�  [      D  , , P;  [ P;  � P�  � P�  [ P;  [      D  , , R�  [ R�  � S  � S  [ R�  [      D  , , T�  [ T�  � Um  � Um  [ T�  [      D  , , W%  [ W%  � W�  � W�  [ W%  [      D  , , Ys  [ Ys  � Z	  � Z	  [ Ys  [      D  , , [�  [ [�  � \W  � \W  [ [�  [      D  , , Ys  ! Ys  !� Z	  !� Z	  ! Ys  !      D  , , [�  ! [�  !� \W  !� \W  ! [�  !      D  , , P;  "[ P;  "� P�  "� P�  "[ P;  "[      D  , , R�  "[ R�  "� S  "� S  "[ R�  "[      D  , , T�  "[ T�  "� Um  "� Um  "[ T�  "[      D  , , W%  "[ W%  "� W�  "� W�  "[ W%  "[      D  , , G  � G  1 G�  1 G�  � G  �      D  , , IQ  � IQ  1 I�  1 I�  � IQ  �      D  , , K�  � K�  1 L5  1 L5  � K�  �      D  , , M�  � M�  1 N�  1 N�  � M�  �      D  , , P;  � P;  1 P�  1 P�  � P;  �      D  , , R�  � R�  1 S  1 S  � R�  �      D  , , T�  � T�  1 Um  1 Um  � T�  �      D  , , W%  � W%  1 W�  1 W�  � W%  �      D  , , Ys  � Ys  1 Z	  1 Z	  � Ys  �      D  , , [�  � [�  1 \W  1 \W  � [�  �      D  , , Ys  "[ Ys  "� Z	  "� Z	  "[ Ys  "[      D  , , [�  "[ [�  "� \W  "� \W  "[ [�  "[      D  , , G  � G  1 G�  1 G�  � G  �      D  , , IQ  � IQ  1 I�  1 I�  � IQ  �      D  , , K�  � K�  1 L5  1 L5  � K�  �      D  , , M�  � M�  1 N�  1 N�  � M�  �      D  , , P;  � P;  1 P�  1 P�  � P;  �      D  , , R�  � R�  1 S  1 S  � R�  �      D  , , T�  � T�  1 Um  1 Um  � T�  �      D  , , W%  � W%  1 W�  1 W�  � W%  �      D  , , Ys  � Ys  1 Z	  1 Z	  � Ys  �      D  , , [�  � [�  1 \W  1 \W  � [�  �      D  , , G  "[ G  "� G�  "� G�  "[ G  "[      D  , , IQ  "[ IQ  "� I�  "� I�  "[ IQ  "[      D  , , G   G  � G�  � G�   G        D  , , IQ   IQ  � I�  � I�   IQ        D  , , K�   K�  � L5  � L5   K�        D  , , M�   M�  � N�  � N�   M�        D  , , P;   P;  � P�  � P�   P;        D  , , R�   R�  � S  � S   R�        D  , , T�   T�  � Um  � Um   T�        D  , , W%   W%  � W�  � W�   W%        D  , , Ys   Ys  � Z	  � Z	   Ys        D  , , [�   [�  � \W  � \W   [�        D  , , G  � G   q G�   q G�  � G  �      D  , , IQ  � IQ   q I�   q I�  � IQ  �      D  , , K�  � K�   q L5   q L5  � K�  �      D  , , n1  � n1  1 n�  1 n�  � n1  �      D  , , p  � p  1 q  1 q  � p  �      D  , , r�  � r�  1 sc  1 sc  � r�  �      D  , , u  � u  1 u�  1 u�  � u  �      D  , , n1  � n1   q n�   q n�  � n1  �      D  , , p  � p   q q   q q  � p  �      D  , , r�  � r�   q sc   q sc  � r�  �      D  , , u  � u   q u�   q u�  � u  �      D  , , `]  � `]  q `�  q `�  � `]  �      D  , , b�  � b�  q cA  q cA  � b�  �      D  , , d�  � d�  q e�  q e�  � d�  �      D  , , gG  � gG  q g�  q g�  � gG  �      D  , , i�  � i�  q j+  q j+  � i�  �      D  , , k�  � k�  q ly  q ly  � k�  �      D  , , n1  � n1  q n�  q n�  � n1  �      D  , , p  � p  q q  q q  � p  �      D  , , r�  � r�  q sc  q sc  � r�  �      D  , , u  � u  q u�  q u�  � u  �      D  , , r�  ! r�  !� sc  !� sc  ! r�  !      D  , , u  ! u  !� u�  !� u�  ! u  !      D  , , i�  "[ i�  "� j+  "� j+  "[ i�  "[      D  , , k�  "[ k�  "� ly  "� ly  "[ k�  "[      D  , , n1  "[ n1  "� n�  "� n�  "[ n1  "[      D  , , p  "[ p  "� q  "� q  "[ p  "[      D  , , r�  "[ r�  "� sc  "� sc  "[ r�  "[      D  , , u  "[ u  "� u�  "� u�  "[ u  "[      D  , , `]  "[ `]  "� `�  "� `�  "[ `]  "[      D  , , b�  "[ b�  "� cA  "� cA  "[ b�  "[      D  , , d�  "[ d�  "� e�  "� e�  "[ d�  "[      D  , , gG  "[ gG  "� g�  "� g�  "[ gG  "[      D  , , `]  ! `]  !� `�  !� `�  ! `]  !      D  , , b�  ! b�  !� cA  !� cA  ! b�  !      D  , , d�  ! d�  !� e�  !� e�  ! d�  !      D  , , gG  ! gG  !� g�  !� g�  ! gG  !      D  , , i�  ! i�  !� j+  !� j+  ! i�  !      D  , , k�  ! k�  !� ly  !� ly  ! k�  !      D  , , n1  ! n1  !� n�  !� n�  ! n1  !      D  , , p  ! p  !� q  !� q  ! p  !      D  , , `]   `]  � `�  � `�   `]        D  , , b�   b�  � cA  � cA   b�        D  , , d�   d�  � e�  � e�   d�        D  , , gG   gG  � g�  � g�   gG        D  , , i�   i�  � j+  � j+   i�        D  , , k�   k�  � ly  � ly   k�        D  , , n1   n1  � n�  � n�   n1        D  , , p   p  � q  � q   p        D  , , r�   r�  � sc  � sc   r�        D  , , u   u  � u�  � u�   u        D  , , `]  � `]   q `�   q `�  � `]  �      D  , , b�  � b�   q cA   q cA  � b�  �      D  , , d�  � d�   q e�   q e�  � d�  �      D  , , gG  � gG   q g�   q g�  � gG  �      D  , , i�  � i�   q j+   q j+  � i�  �      D  , , k�  � k�   q ly   q ly  � k�  �      D  , , `]  � `]  1 `�  1 `�  � `]  �      D  , , b�  � b�  1 cA  1 cA  � b�  �      D  , , `]  � `]  1 `�  1 `�  � `]  �      D  , , b�  � b�  1 cA  1 cA  � b�  �      D  , , d�  � d�  1 e�  1 e�  � d�  �      D  , , gG  � gG  1 g�  1 g�  � gG  �      D  , , i�  � i�  1 j+  1 j+  � i�  �      D  , , k�  � k�  1 ly  1 ly  � k�  �      D  , , n1  � n1  1 n�  1 n�  � n1  �      D  , , p  � p  1 q  1 q  � p  �      D  , , r�  � r�  1 sc  1 sc  � r�  �      D  , , u  � u  1 u�  1 u�  � u  �      D  , , d�  � d�  1 e�  1 e�  � d�  �      D  , , gG  � gG  1 g�  1 g�  � gG  �      D  , , `]  [ `]  � `�  � `�  [ `]  [      D  , , b�  [ b�  � cA  � cA  [ b�  [      D  , , d�  [ d�  � e�  � e�  [ d�  [      D  , , gG  [ gG  � g�  � g�  [ gG  [      D  , , i�  [ i�  � j+  � j+  [ i�  [      D  , , k�  [ k�  � ly  � ly  [ k�  [      D  , , n1  [ n1  � n�  � n�  [ n1  [      D  , , p  [ p  � q  � q  [ p  [      D  , , r�  [ r�  � sc  � sc  [ r�  [      D  , , u  [ u  � u�  � u�  [ u  [      D  , , i�  � i�  1 j+  1 j+  � i�  �      D  , , k�  � k�  1 ly  1 ly  � k�  �      D  , , -�  .� -�  /� .b  /� .b  .� -�  .�      D  , , -�  1o -�  2 .b  2 .b  1o -�  1o      D  , , ,�  %� ,�  & -;  & -;  %� ,�  %�      D  , , -�  )� -�  *� .b  *� .b  )� -�  )�      D  , , -�  -� -�  .E .b  .E .b  -� -�  -�      D  , , -�  ,o -�  - .b  - .b  ,o -�  ,o      D  , , -�  2� -�  3E .b  3E .b  2� -�  2�      D  , , -�  +/ -�  +� .b  +� .b  +/ -�  +/      D  , , -�  0/ -�  0� .b  0� .b  0/ -�  0/      D  , , ,�  &� ,�  '[ -;  '[ -;  &� ,�  &�      D  , , +~  .� +~  /� ,  /� ,  .� +~  .�      D  , , �  1o �  2  �  2  �  1o �  1o      D  , , "F  1o "F  2 "�  2 "�  1o "F  1o      D  , , $�  1o $�  2 %*  2 %*  1o $�  1o      D  , , &�  1o &�  2 'x  2 'x  1o &�  1o      D  , , )0  1o )0  2 )�  2 )�  1o )0  1o      D  , , +~  1o +~  2 ,  2 ,  1o +~  1o      D  , , �  -� �  .E  �  .E  �  -� �  -�      D  , , "F  -� "F  .E "�  .E "�  -� "F  -�      D  , , $�  -� $�  .E %*  .E %*  -� $�  -�      D  , , &�  -� &�  .E 'x  .E 'x  -� &�  -�      D  , , )0  -� )0  .E )�  .E )�  -� )0  -�      D  , , +~  -� +~  .E ,  .E ,  -� +~  -�      D  , , &�  ,o &�  - 'x  - 'x  ,o &�  ,o      D  , , )0  ,o )0  - )�  - )�  ,o )0  ,o      D  , , +~  ,o +~  - ,  - ,  ,o +~  ,o      D  , , �  .� �  /�  �  /�  �  .� �  .�      D  , , +~  2� +~  3E ,  3E ,  2� +~  2�      D  , , "F  .� "F  /� "�  /� "�  .� "F  .�      D  , , �  0/ �  0�  �  0�  �  0/ �  0/      D  , , $�  .� $�  /� %*  /� %*  .� $�  .�      D  , , "F  0/ "F  0� "�  0� "�  0/ "F  0/      D  , , $�  0/ $�  0� %*  0� %*  0/ $�  0/      D  , , &�  0/ &�  0� 'x  0� 'x  0/ &�  0/      D  , , )0  0/ )0  0� )�  0� )�  0/ )0  0/      D  , , +~  0/ +~  0� ,  0� ,  0/ +~  0/      D  , , &�  .� &�  /� 'x  /� 'x  .� &�  .�      D  , , �  2� �  3E  �  3E  �  2� �  2�      D  , , �  ,o �  -  �  -  �  ,o �  ,o      D  , , "F  ,o "F  - "�  - "�  ,o "F  ,o      D  , , $�  ,o $�  - %*  - %*  ,o $�  ,o      D  , , "F  2� "F  3E "�  3E "�  2� "F  2�      D  , , $�  2� $�  3E %*  3E %*  2� $�  2�      D  , , &�  2� &�  3E 'x  3E 'x  2� &�  2�      D  , , )0  2� )0  3E )�  3E )�  2� )0  2�      D  , , )0  .� )0  /� )�  /� )�  .� )0  .�      D  , , �  0/ �  0� @  0� @  0/ �  0/      D  , , \  .� \  /� �  /� �  .� \  .�      D  , , �  -� �  .E @  .E @  -� �  -�      D  , , r  .� r  /�   /�   .� r  .�      D  , , r  1o r  2   2   1o r  1o      D  , , �  1o �  2 V  2 V  1o �  1o      D  , ,   1o   2 �  2 �  1o   1o      D  , , \  1o \  2 �  2 �  1o \  1o      D  , , �  1o �  2 @  2 @  1o �  1o      D  , , r  0/ r  0�   0�   0/ r  0/      D  , , �  0/ �  0� V  0� V  0/ �  0/      D  , ,   2�   3E �  3E �  2�   2�      D  , , \  2� \  3E �  3E �  2� \  2�      D  , , �  2� �  3E @  3E @  2� �  2�      D  , , �  .� �  /� @  /� @  .� �  .�      D  , , r  ,o r  -   -   ,o r  ,o      D  , , �  ,o �  - V  - V  ,o �  ,o      D  , ,   ,o   - �  - �  ,o   ,o      D  , , \  ,o \  - �  - �  ,o \  ,o      D  , , �  ,o �  - @  - @  ,o �  ,o      D  , , �  .� �  /� V  /� V  .� �  .�      D  , ,   .�   /� �  /� �  .�   .�      D  , , r  -� r  .E   .E   -� r  -�      D  , , �  -� �  .E V  .E V  -� �  -�      D  , ,   -�   .E �  .E �  -�   -�      D  , , \  -� \  .E �  .E �  -� \  -�      D  , ,   0/   0� �  0� �  0/   0/      D  , , \  0/ \  0� �  0� �  0/ \  0/      D  , , r  2� r  3E   3E   2� r  2�      D  , , �  2� �  3E V  3E V  2� �  2�      D  , , r  +/ r  +�   +�   +/ r  +/      D  , , �  +/ �  +� @  +� @  +/ �  +/      D  , , �  +/ �  +� V  +� V  +/ �  +/      D  , ,   +/   +� �  +� �  +/   +/      D  , , \  +/ \  +� �  +� �  +/ \  +/      D  , , r  )� r  *�   *�   )� r  )�      D  , , �  )� �  *� V  *� V  )� �  )�      D  , , K  %� K  & �  & �  %� K  %�      D  , , �  %� �  & /  & /  %� �  %�      D  , , �  %� �  &   &   %� �  %�      D  , , �  %� �  & g  & g  %� �  %�      D  , , �  %� �  & }  & }  %� �  %�      D  , , 5  %� 5  & �  & �  %� 5  %�      D  , , K  &� K  '[ �  '[ �  &� K  &�      D  , , �  &� �  '[ /  '[ /  &� �  &�      D  , , �  &� �  '[ }  '[ }  &� �  &�      D  , , 5  &� 5  '[ �  '[ �  &� 5  &�      D  , , �  &� �  '[   '[   &� �  &�      D  , , �  &� �  '[ g  '[ g  &� �  &�      D  , ,   )�   *� �  *� �  )�   )�      D  , , \  )� \  *� �  *� �  )� \  )�      D  , , �  )� �  *� @  *� @  )� �  )�      D  , , %�  %� %�  & &Q  & &Q  %� %�  %�      D  , , (	  %� (	  & (�  & (�  %� (	  %�      D  , , �  )� �  *�  �  *�  �  )� �  )�      D  , , "F  )� "F  *� "�  *� "�  )� "F  )�      D  , , $�  )� $�  *� %*  *� %*  )� $�  )�      D  , , !  %� !  & !�  & !�  %� !  %�      D  , , #m  %� #m  & $  & $  %� #m  %�      D  , , �  +/ �  +�  �  +�  �  +/ �  +/      D  , , "F  +/ "F  +� "�  +� "�  +/ "F  +/      D  , , $�  +/ $�  +� %*  +� %*  +/ $�  +/      D  , , &�  +/ &�  +� 'x  +� 'x  +/ &�  +/      D  , , )0  +/ )0  +� )�  +� )�  +/ )0  +/      D  , , +~  +/ +~  +� ,  +� ,  +/ +~  +/      D  , , &�  )� &�  *� 'x  *� 'x  )� &�  )�      D  , , !  &� !  '[ !�  '[ !�  &� !  &�      D  , , #m  &� #m  '[ $  '[ $  &� #m  &�      D  , , %�  &� %�  '[ &Q  '[ &Q  &� %�  &�      D  , , (	  &� (	  '[ (�  '[ (�  &� (	  &�      D  , , *W  &� *W  '[ *�  '[ *�  &� *W  &�      D  , , )0  )� )0  *� )�  *� )�  )� )0  )�      D  , , +~  )� +~  *� ,  *� ,  )� +~  )�      D  , , *W  %� *W  & *�  & *�  %� *W  %�      D  , , �  � �  q V  q V  � �  �      D  , ,   �   q �  q �  �   �      D  , , \  � \  q �  q �  � \  �      D  , , �  � �  q @  q @  � �  �      D  , , �  � �  q  �  q  �  � �  �      D  , , "F  � "F  q "�  q "�  � "F  �      D  , , r  "[ r  "�   "�   "[ r  "[      D  , , �  "[ �  "� V  "� V  "[ �  "[      D  , ,   "[   "� �  "� �  "[   "[      D  , , \  "[ \  "� �  "� �  "[ \  "[      D  , , r  � r   q    q   � r  �      D  , , �  � �   q V   q V  � �  �      D  , ,   �    q �   q �  �   �      D  , , \  � \   q �   q �  � \  �      D  , , �  � �   q @   q @  � �  �      D  , , �  � �   q  �   q  �  � �  �      D  , , r  [ r  �   �   [ r  [      D  , , �  [ �  � V  � V  [ �  [      D  , ,   [   � �  � �  [   [      D  , , \  [ \  � �  � �  [ \  [      D  , , �  [ �  � @  � @  [ �  [      D  , , �  [ �  �  �  �  �  [ �  [      D  , , $�  � $�  q %*  q %*  � $�  �      D  , , &�  � &�  q 'x  q 'x  � &�  �      D  , , )0  � )0  q )�  q )�  � )0  �      D  , , +~  � +~  q ,  q ,  � +~  �      D  , , r  � r  1   1   � r  �      D  , , �  � �  1 V  1 V  � �  �      D  , ,   �   1 �  1 �  �   �      D  , , \  � \  1 �  1 �  � \  �      D  , , �  � �  1 @  1 @  � �  �      D  , , �  � �  1  �  1  �  � �  �      D  , , "F  � "F  1 "�  1 "�  � "F  �      D  , , $�  � $�  1 %*  1 %*  � $�  �      D  , , &�  � &�  1 'x  1 'x  � &�  �      D  , , )0  � )0  1 )�  1 )�  � )0  �      D  , , +~  � +~  1 ,  1 ,  � +~  �      D  , , "F  [ "F  � "�  � "�  [ "F  [      D  , , $�  [ $�  � %*  � %*  [ $�  [      D  , , &�  [ &�  � 'x  � 'x  [ &�  [      D  , , )0  [ )0  � )�  � )�  [ )0  [      D  , , +~  [ +~  � ,  � ,  [ +~  [      D  , , "F  � "F   q "�   q "�  � "F  �      D  , , $�  � $�   q %*   q %*  � $�  �      D  , , &�  � &�   q 'x   q 'x  � &�  �      D  , , )0  � )0   q )�   q )�  � )0  �      D  , , +~  � +~   q ,   q ,  � +~  �      D  , , �  "[ �  "� @  "� @  "[ �  "[      D  , , �  "[ �  "�  �  "�  �  "[ �  "[      D  , , �   �  �  �  �  �   �        D  , , "F   "F  � "�  � "�   "F        D  , , $�   $�  � %*  � %*   $�        D  , , &�   &�  � 'x  � 'x   &�        D  , , )0   )0  � )�  � )�   )0        D  , , +~   +~  � ,  � ,   +~        D  , , &�  "[ &�  "� 'x  "� 'x  "[ &�  "[      D  , , )0  "[ )0  "� )�  "� )�  "[ )0  "[      D  , , �  � �  1 @  1 @  � �  �      D  , , �  � �  1  �  1  �  � �  �      D  , , "F  � "F  1 "�  1 "�  � "F  �      D  , , $�  � $�  1 %*  1 %*  � $�  �      D  , , &�  � &�  1 'x  1 'x  � &�  �      D  , , )0  � )0  1 )�  1 )�  � )0  �      D  , , +~  � +~  1 ,  1 ,  � +~  �      D  , , +~  "[ +~  "� ,  "� ,  "[ +~  "[      D  , , r   r  �   �    r        D  , , r  � r  1   1   � r  �      D  , , �  � �  1 V  1 V  � �  �      D  , ,   �   1 �  1 �  �   �      D  , , \  � \  1 �  1 �  � \  �      D  , , �   �  � V  � V   �        D  , ,      � �  � �           D  , , \   \  � �  � �   \        D  , , r  ! r  !�   !�   ! r  !      D  , , �  ! �  !� V  !� V  ! �  !      D  , ,   !   !� �  !� �  !   !      D  , , \  ! \  !� �  !� �  ! \  !      D  , , �  ! �  !� @  !� @  ! �  !      D  , , �  ! �  !�  �  !�  �  ! �  !      D  , , "F  ! "F  !� "�  !� "�  ! "F  !      D  , , $�  ! $�  !� %*  !� %*  ! $�  !      D  , , &�  ! &�  !� 'x  !� 'x  ! &�  !      D  , , )0  ! )0  !� )�  !� )�  ! )0  !      D  , , +~  ! +~  !� ,  !� ,  ! +~  !      D  , , "F  "[ "F  "� "�  "� "�  "[ "F  "[      D  , , $�  "[ $�  "� %*  "� %*  "[ $�  "[      D  , , �   �  � @  � @   �        D  , , r  � r  q   q   � r  �      D  , , -�  � -�   q .b   q .b  � -�  �      D  , , -�  [ -�  � .b  � .b  [ -�  [      D  , , -�  � -�  q .b  q .b  � -�  �      D  , , -�  ! -�  !� .b  !� .b  ! -�  !      D  , , -�   -�  � .b  � .b   -�        D  , , -�  "[ -�  "� .b  "� .b  "[ -�  "[      D  , , -�  � -�  1 .b  1 .b  � -�  �      D  , , -�  � -�  1 .b  1 .b  � -�  �      D  , ,  ��  w  ��    �2    �2  w  ��  w      D  , ,  ��  7  ��  �  �2  �  �2  7  ��  7      D  , ,  ��  �  ��  �  �2  �  �2  �  ��  �      D  , ,  ��  �  ��  M  �2  M  �2  �  ��  �      D  , ,  ��  w  ��    �2    �2  w  ��  w      D  , ,  ��  7  ��  �  �2  �  �2  7  ��  7      D  , ,  ��  �  ��  �  �2  �  �2  �  ��  �      D  , ,  ��  �  ��  M  �2  M  �2  �  ��  �      D  , ,  ��  #  ��  �  �2  �  �2  #  ��  #      D  , ,  ��  �  ��  y  �2  y  �2  �  ��  �      D  , ,  ��  �  ��  9  �2  9  �2  �  ��  �      D  , ,  ��  c  ��  �  �2  �  �2  c  ��  c      D  , ,  ��   #  ��   �  �2   �  �2   #  ��   #      D  , ,  ������  �����y  �2���y  �2����  ������      D  , ,  ������  �����9  �2���9  �2����  ������      D  , ,  �����c  ������  �2����  �2���c  �����c      D  , ,  �����m  �����  �2���  �2���m  �����m      D  , ,  �����-  ������  �2����  �2���-  �����-      D  , ,  ������  �����  �2���  �2����  ������      D  , ,  �����  �����C  �2���C  �2���  �����      D  , ,  �����m  �����  �2���  �2���m  �����m      D  , ,  �����-  ������  �2����  �2���-  �����-      D  , ,  ������  �����  �2���  �2����  ������      D  , ,  �����  �����C  �2���C  �2���  �����      D  , ,  �����  ����ݯ  �2��ݯ  �2���  �����      D  , ,  ������  �����o  �2���o  �2����  ������      D  , ,  ����ڙ  �����/  �2���/  �2��ڙ  ����ڙ      D  , ,  �����Y  ������  �2����  �2���Y  �����Y      D  , ,  �����  ����د  �2��د  �2���  �����      D  , ,  ������  �����o  �2���o  �2����  ������      D  , ,  ����ՙ  �����/  �2���/  �2��ՙ  ����ՙ      D  , ,  �����Y  ������  �2����  �2���Y  �����Y      D  , ,  �����c  ������  �F����  �F���c  �����c      D  , ,  �����#  ����Ĺ  �F��Ĺ  �F���#  �����#      D  , ,  ������  �����y  �F���y  �F����  ������      D  , ,  ������  �����9  �F���9  �F����  ������      D  , ,  �����c  ������  �F����  �F���c  �����c      D  , ,  ��  %�  ��  &  ��  &  ��  %�  ��  %�      D  , ,  ��  &�  ��  '[  ��  '[  ��  &�  ��  &�      D  , , �  1o �  2 4  2 4  1o �  1o      D  , , �  2� �  3E 4  3E 4  2� �  2�      D  , , �  )� �  *� 4  *� 4  )� �  )�      D  , , �  .� �  /� 4  /� 4  .� �  .�      D  , , �  +/ �  +� 4  +� 4  +/ �  +/      D  , , �  ,o �  - 4  - 4  ,o �  ,o      D  , , �  -� �  .E 4  .E 4  -� �  -�      D  , , �  0/ �  0� 4  0� 4  0/ �  0/      D  , , :  1o :  2 �  2 �  1o :  1o      D  , , �  1o �  2   2   1o �  1o      D  , , �  .� �  /� 	�  /� 	�  .� �  .�      D  , , :  .� :  /� �  /� �  .� :  .�      D  , , �  .� �  /�   /�   .� �  .�      D  , , �  .� �  /� l  /� l  .� �  .�      D  , , $  .� $  /� �  /� �  .� $  .�      D  , , :  2� :  3E �  3E �  2� :  2�      D  , , �  2� �  3E   3E   2� �  2�      D  , , �  2� �  3E l  3E l  2� �  2�      D  , , $  2� $  3E �  3E �  2� $  2�      D  , , �  1o �  2 l  2 l  1o �  1o      D  , , $  1o $  2 �  2 �  1o $  1o      D  , , �  ,o �  - 	�  - 	�  ,o �  ,o      D  , , :  ,o :  - �  - �  ,o :  ,o      D  , , �  ,o �  -   -   ,o �  ,o      D  , , �  ,o �  - l  - l  ,o �  ,o      D  , , $  ,o $  - �  - �  ,o $  ,o      D  , , �  1o �  2 	�  2 	�  1o �  1o      D  , , �  -� �  .E 	�  .E 	�  -� �  -�      D  , , :  -� :  .E �  .E �  -� :  -�      D  , , �  -� �  .E   .E   -� �  -�      D  , , �  -� �  .E l  .E l  -� �  -�      D  , , $  -� $  .E �  .E �  -� $  -�      D  , , �  2� �  3E 	�  3E 	�  2� �  2�      D  , , �  0/ �  0� 	�  0� 	�  0/ �  0/      D  , , :  0/ :  0� �  0� �  0/ :  0/      D  , , �  0/ �  0�   0�   0/ �  0/      D  , , �  0/ �  0� l  0� l  0/ �  0/      D  , , $  0/ $  0� �  0� �  0/ $  0/      D  , ,  ��  .�  ��  /�  J  /�  J  .�  ��  .�      D  , ,   .�   /� �  /� �  .�   .�      D  , , P  .� P  /� �  /� �  .� P  .�      D  , , P  1o P  2 �  2 �  1o P  1o      D  , ,  �  .�  �  /�  ��  /�  ��  .�  �  .�      D  , ,   1o   2 �  2 �  1o   1o      D  , ,  �f  1o  �f  2  ��  2  ��  1o  �f  1o      D  , ,  �f  .�  �f  /�  ��  /�  ��  .�  �f  .�      D  , ,  �  -�  �  .E  ��  .E  ��  -�  �  -�      D  , ,  �f  -�  �f  .E  ��  .E  ��  -�  �f  -�      D  , ,  ��  -�  ��  .E  J  .E  J  -�  ��  -�      D  , ,   -�   .E �  .E �  -�   -�      D  , ,  �  0/  �  0�  ��  0�  ��  0/  �  0/      D  , ,  �f  0/  �f  0�  ��  0�  ��  0/  �f  0/      D  , ,  ��  0/  ��  0�  J  0�  J  0/  ��  0/      D  , ,  ��  1o  ��  2  J  2  J  1o  ��  1o      D  , ,   0/   0� �  0� �  0/   0/      D  , , P  0/ P  0� �  0� �  0/ P  0/      D  , , P  -� P  .E �  .E �  -� P  -�      D  , ,  �  ,o  �  -  ��  -  ��  ,o  �  ,o      D  , ,  �f  ,o  �f  -  ��  -  ��  ,o  �f  ,o      D  , ,  ��  ,o  ��  -  J  -  J  ,o  ��  ,o      D  , ,   ,o   - �  - �  ,o   ,o      D  , , P  ,o P  - �  - �  ,o P  ,o      D  , ,  �  2�  �  3E  ��  3E  ��  2�  �  2�      D  , ,  �f  2�  �f  3E  ��  3E  ��  2�  �f  2�      D  , ,  ��  2�  ��  3E  J  3E  J  2�  ��  2�      D  , ,   2�   3E �  3E �  2�   2�      D  , , P  2� P  3E �  3E �  2� P  2�      D  , ,  �  1o  �  2  ��  2  ��  1o  �  1o      D  , ,  �f  +/  �f  +�  ��  +�  ��  +/  �f  +/      D  , ,  �?  &�  �?  '[  ��  '[  ��  &�  �?  &�      D  , ,  ��  &�  ��  '[  �#  '[  �#  &�  ��  &�      D  , ,  �  &�  �  '[ q  '[ q  &�  �  &�      D  , , )  &� )  '[ �  '[ �  &� )  &�      D  , , w  &� w  '[   '[   &� w  &�      D  , ,  ��  +/  ��  +�  J  +�  J  +/  ��  +/      D  , ,   +/   +� �  +� �  +/   +/      D  , , P  +/ P  +� �  +� �  +/ P  +/      D  , ,  �f  )�  �f  *�  ��  *�  ��  )�  �f  )�      D  , ,  ��  )�  ��  *�  J  *�  J  )�  ��  )�      D  , ,   )�   *� �  *� �  )�   )�      D  , , P  )� P  *� �  *� �  )� P  )�      D  , ,  �  )�  �  *�  ��  *�  ��  )�  �  )�      D  , ,  �?  %�  �?  &  ��  &  ��  %�  �?  %�      D  , ,  ��  %�  ��  &  �#  &  �#  %�  ��  %�      D  , ,  �  %�  �  & q  & q  %�  �  %�      D  , , )  %� )  & �  & �  %� )  %�      D  , , w  %� w  &   &   %� w  %�      D  , ,  �  +/  �  +�  ��  +�  ��  +/  �  +/      D  , , 
  %� 
  & 
�  & 
�  %� 
  %�      D  , , �  &� �  '[ [  '[ [  &� �  &�      D  , , 
  &� 
  '[ 
�  '[ 
�  &� 
  &�      D  , , a  &� a  '[ �  '[ �  &� a  &�      D  , , �  &� �  '[ E  '[ E  &� �  &�      D  , , �  &� �  '[ �  '[ �  &� �  &�      D  , , a  %� a  & �  & �  %� a  %�      D  , , �  %� �  & E  & E  %� �  %�      D  , , �  %� �  & �  & �  %� �  %�      D  , , �  )� �  *� 	�  *� 	�  )� �  )�      D  , , :  )� :  *� �  *� �  )� :  )�      D  , , �  )� �  *�   *�   )� �  )�      D  , , �  )� �  *� l  *� l  )� �  )�      D  , , $  )� $  *� �  *� �  )� $  )�      D  , , �  %� �  & [  & [  %� �  %�      D  , , �  +/ �  +� 	�  +� 	�  +/ �  +/      D  , , :  +/ :  +� �  +� �  +/ :  +/      D  , , �  +/ �  +�   +�   +/ �  +/      D  , , �  +/ �  +� l  +� l  +/ �  +/      D  , , $  +/ $  +� �  +� �  +/ $  +/      D  , ,  ��  +/  ��  +�  �`  +�  �`  +/  ��  +/      D  , ,  �|  )�  �|  *�  �  *�  �  )�  �|  )�      D  , ,  ��  )�  ��  *�  �`  *�  �`  )�  ��  )�      D  , ,  �|  .�  �|  /�  �  /�  �  .�  �|  .�      D  , ,  �U  %�  �U  &  ��  &  ��  %�  �U  %�      D  , ,  ��  %�  ��  &  �9  &  �9  %�  ��  %�      D  , ,  ��  .�  ��  /�  �`  /�  �`  .�  ��  .�      D  , ,  �.  .�  �.  /�  ��  /�  ��  .�  �.  .�      D  , ,  �.  )�  �.  *�  ��  *�  ��  )�  �.  )�      D  , ,  �.  2�  �.  3E  ��  3E  ��  2�  �.  2�      D  , ,  �|  2�  �|  3E  �  3E  �  2�  �|  2�      D  , ,  �.  0/  �.  0�  ��  0�  ��  0/  �.  0/      D  , ,  ��  -�  ��  .E  �`  .E  �`  -�  ��  -�      D  , ,  �|  0/  �|  0�  �  0�  �  0/  �|  0/      D  , ,  �.  -�  �.  .E  ��  .E  ��  -�  �.  -�      D  , ,  �|  -�  �|  .E  �  .E  �  -�  �|  -�      D  , ,  �.  +/  �.  +�  ��  +�  ��  +/  �.  +/      D  , ,  ��  0/  ��  0�  �`  0�  �`  0/  ��  0/      D  , ,  ��  2�  ��  3E  �`  3E  �`  2�  ��  2�      D  , ,  �|  +/  �|  +�  �  +�  �  +/  �|  +/      D  , ,  �.  ,o  �.  -  ��  -  ��  ,o  �.  ,o      D  , ,  �|  ,o  �|  -  �  -  �  ,o  �|  ,o      D  , ,  �U  &�  �U  '[  ��  '[  ��  &�  �U  &�      D  , ,  ��  &�  ��  '[  �9  '[  �9  &�  ��  &�      D  , ,  �.  1o  �.  2  ��  2  ��  1o  �.  1o      D  , ,  �|  1o  �|  2  �  2  �  1o  �|  1o      D  , ,  ��  1o  ��  2  �`  2  �`  1o  ��  1o      D  , ,  ��  ,o  ��  -  �`  -  �`  ,o  ��  ,o      D  , ,  �|  �  �|  1  �  1  �  �  �|  �      D  , ,  ��  �  ��  1  �`  1  �`  �  ��  �      D  , ,  �.  �  �.  1  ��  1  ��  �  �.  �      D  , ,  �|  �  �|  1  �  1  �  �  �|  �      D  , ,  ��  �  ��  1  �`  1  �`  �  ��  �      D  , ,  �|  �  �|   q  �   q  �  �  �|  �      D  , ,  ��  �  ��   q  �`   q  �`  �  ��  �      D  , ,  �|    �|  �  �  �  �    �|        D  , ,  �.  �  �.  q  ��  q  ��  �  �.  �      D  , ,  �|  �  �|  q  �  q  �  �  �|  �      D  , ,  ��  �  ��  q  �`  q  �`  �  ��  �      D  , ,  ��    ��  �  �`  �  �`    ��        D  , ,  �.    �.  �  ��  �  ��    �.        D  , ,  �.  [  �.  �  ��  �  ��  [  �.  [      D  , ,  �|  [  �|  �  �  �  �  [  �|  [      D  , ,  ��  [  ��  �  �`  �  �`  [  ��  [      D  , ,  �.  �  �.   q  ��   q  ��  �  �.  �      D  , ,  �.  "[  �.  "�  ��  "�  ��  "[  �.  "[      D  , ,  �|  "[  �|  "�  �  "�  �  "[  �|  "[      D  , ,  ��  "[  ��  "�  �`  "�  �`  "[  ��  "[      D  , ,  �.  �  �.  1  ��  1  ��  �  �.  �      D  , ,  �.  !  �.  !�  ��  !�  ��  !  �.  !      D  , ,  �|  !  �|  !�  �  !�  �  !  �|  !      D  , ,  ��  !  ��  !�  �`  !�  �`  !  ��  !      D  , , �   �  � 4  � 4   �        D  , , �   �  � 	�  � 	�   �        D  , ,  �  �  �  1  ��  1  ��  �  �  �      D  , ,  �f  �  �f  1  ��  1  ��  �  �f  �      D  , ,  ��  �  ��  1  J  1  J  �  ��  �      D  , ,   �   1 �  1 �  �   �      D  , , P  � P  1 �  1 �  � P  �      D  , , �  � �  1 4  1 4  � �  �      D  , , �  � �  1 	�  1 	�  � �  �      D  , , :  � :  1 �  1 �  � :  �      D  , , �  � �  1   1   � �  �      D  , , �  � �  1 l  1 l  � �  �      D  , , $  � $  1 �  1 �  � $  �      D  , , �  "[ �  "� 	�  "� 	�  "[ �  "[      D  , , :  "[ :  "� �  "� �  "[ :  "[      D  , , �  "[ �  "�   "�   "[ �  "[      D  , , �  "[ �  "� l  "� l  "[ �  "[      D  , , $  "[ $  "� �  "� �  "[ $  "[      D  , , :   :  � �  � �   :        D  , , �   �  �   �    �        D  , , �   �  � l  � l   �        D  , ,  �  �  �  1  ��  1  ��  �  �  �      D  , ,  �f  �  �f  1  ��  1  ��  �  �f  �      D  , ,  ��  �  ��  1  J  1  J  �  ��  �      D  , ,   �   1 �  1 �  �   �      D  , , P  � P  1 �  1 �  � P  �      D  , , �  � �  1 4  1 4  � �  �      D  , , �  � �  1 	�  1 	�  � �  �      D  , , :  � :  1 �  1 �  � :  �      D  , , �  � �  1   1   � �  �      D  , , �  � �  1 l  1 l  � �  �      D  , , $  � $  1 �  1 �  � $  �      D  , , $   $  � �  � �   $        D  , , �  ! �  !�   !�   ! �  !      D  , , �  ! �  !� l  !� l  ! �  !      D  , , $  ! $  !� �  !� �  ! $  !      D  , ,  �  �  �  q  ��  q  ��  �  �  �      D  , ,  �f  �  �f  q  ��  q  ��  �  �f  �      D  , ,  ��  �  ��  q  J  q  J  �  ��  �      D  , ,   �   q �  q �  �   �      D  , , P  � P  q �  q �  � P  �      D  , , �  � �  q 4  q 4  � �  �      D  , , �  � �  q 	�  q 	�  � �  �      D  , , :  � :  q �  q �  � :  �      D  , , �  � �  q   q   � �  �      D  , , �  � �  q l  q l  � �  �      D  , , $  � $  q �  q �  � $  �      D  , ,  �    �  �  ��  �  ��    �        D  , ,  �f    �f  �  ��  �  ��    �f        D  , ,  ��    ��  �  J  �  J    ��        D  , ,      � �  � �           D  , , P   P  � �  � �   P        D  , ,  �  �  �   q  ��   q  ��  �  �  �      D  , ,  �f  �  �f   q  ��   q  ��  �  �f  �      D  , ,  ��  �  ��   q  J   q  J  �  ��  �      D  , ,   �    q �   q �  �   �      D  , , P  � P   q �   q �  � P  �      D  , , �  � �   q 4   q 4  � �  �      D  , , �  � �   q 	�   q 	�  � �  �      D  , , :  � :   q �   q �  � :  �      D  , , �  � �   q    q   � �  �      D  , ,  �  [  �  �  ��  �  ��  [  �  [      D  , ,  �f  [  �f  �  ��  �  ��  [  �f  [      D  , ,  ��  [  ��  �  J  �  J  [  ��  [      D  , ,   [   � �  � �  [   [      D  , , P  [ P  � �  � �  [ P  [      D  , , �  [ �  � 4  � 4  [ �  [      D  , , �  [ �  � 	�  � 	�  [ �  [      D  , , :  [ :  � �  � �  [ :  [      D  , , �  [ �  �   �   [ �  [      D  , , �  [ �  � l  � l  [ �  [      D  , , $  [ $  � �  � �  [ $  [      D  , , �  � �   q l   q l  � �  �      D  , ,  �  "[  �  "�  ��  "�  ��  "[  �  "[      D  , ,  �f  "[  �f  "�  ��  "�  ��  "[  �f  "[      D  , ,  ��  "[  ��  "�  J  "�  J  "[  ��  "[      D  , ,   "[   "� �  "� �  "[   "[      D  , , P  "[ P  "� �  "� �  "[ P  "[      D  , , �  "[ �  "� 4  "� 4  "[ �  "[      D  , , $  � $   q �   q �  � $  �      D  , ,  �  !  �  !�  ��  !�  ��  !  �  !      D  , ,  �f  !  �f  !�  ��  !�  ��  !  �f  !      D  , ,  ��  !  ��  !�  J  !�  J  !  ��  !      D  , ,   !   !� �  !� �  !   !      D  , , P  ! P  !� �  !� �  ! P  !      D  , , �  ! �  !� 4  !� 4  ! �  !      D  , , �  ! �  !� 	�  !� 	�  ! �  !      D  , , :  ! :  !� �  !� �  ! :  !      D  , ,  ̜  �  ̜    �2    �2  �  ̜  �      D  , ,  �8  �  �8    ��    ��  �  �8  �      D  , ,  ��  �  ��    ��    ��  �  ��  �      D  , ,  ��  �  ��    �&    �&  �  ��  �      D  , ,  �  &�  �  'Q  ��  'Q  ��  &�  �  &�      D  , ,  �g  &�  �g  'Q  ��  'Q  ��  &�  �g  &�      D  , ,  ��  �  ��  _  �&  _  �&  �  ��  �      D  , ,  �,  �  �,  _  ��  _  ��  �  �,  �      D  , ,  ��  �  ��  _  �^  _  �^  �  ��  �      D  , ,  �d  �  �d  _  ��  _  ��  �  �d  �      D  , ,  �   �  �   _  Ȗ  _  Ȗ  �  �   �      D  , ,  ̜  �  ̜  _  �2  _  �2  �  ̜  �      D  , ,  �8  �  �8  _  ��  _  ��  �  �8  �      D  , ,  ��  &�  ��  'Q  �K  'Q  �K  &�  ��  &�      D  , ,  �  &�  �  'Q  ��  'Q  ��  &�  �  &�      D  , ,  �Q  &�  �Q  'Q  ��  'Q  ��  &�  �Q  &�      D  , ,  ��  &�  ��  'Q  �5  'Q  �5  &�  ��  &�      D  , ,  ��  &�  ��  'Q  ��  'Q  ��  &�  ��  &�      D  , ,  �;  &�  �;  'Q  ��  'Q  ��  &�  �;  &�      D  , ,  ��  &�  ��  'Q  �  'Q  �  &�  ��  &�      D  , ,  ��  &�  ��  'Q  �m  'Q  �m  &�  ��  &�      D  , ,  �%  &�  �%  'Q  ƻ  'Q  ƻ  &�  �%  &�      D  , ,  �s  &�  �s  'Q  �	  'Q  �	  &�  �s  &�      D  , ,  �,  �  �,    ��    ��  �  �,  �      D  , ,  ��  �  ��    �^    �^  �  ��  �      D  , ,  ��  	  ��  �  ��  �  ��  	  ��  	      D  , ,  ��  	  ��  �  �&  �  �&  	  ��  	      D  , ,  �,  	  �,  �  ��  �  ��  	  �,  	      D  , ,  ��  	  ��  �  �^  �  �^  	  ��  	      D  , ,  �d  	  �d  �  ��  �  ��  	  �d  	      D  , ,  �   	  �   �  Ȗ  �  Ȗ  	  �   	      D  , ,  ̜  	  ̜  �  �2  �  �2  	  ̜  	      D  , ,  �8  	  �8  �  ��  �  ��  	  �8  	      D  , ,  �d  �  �d    ��    ��  �  �d  �      D  , ,  �   �  �     Ȗ    Ȗ  �  �   �      D  , ,  ��  I  ��  �  ��  �  ��  I  ��  I      D  , ,  ��  I  ��  �  �&  �  �&  I  ��  I      D  , ,  �,  I  �,  �  ��  �  ��  I  �,  I      D  , ,  ��  I  ��  �  �^  �  �^  I  ��  I      D  , ,  �d  I  �d  �  ��  �  ��  I  �d  I      D  , ,  �   I  �   �  Ȗ  �  Ȗ  I  �   I      D  , ,  ̜  I  ̜  �  �2  �  �2  I  ̜  I      D  , ,  �8  I  �8  �  ��  �  ��  I  �8  I      D  , ,  ��  �  ��  _  ��  _  ��  �  ��  �      D  , ,  �   �  �   �  Ȗ  �  Ȗ  �  �   �      D  , ,  �   �  �   M  Ȗ  M  Ȗ  �  �   �      D  , ,  �   w  �     Ȗ    Ȗ  w  �   w      D  , ,  �   7  �   �  Ȗ  �  Ȗ  7  �   7      D  , ,  �   �  �   �  Ȗ  �  Ȗ  �  �   �      D  , ,  �   �  �   M  Ȗ  M  Ȗ  �  �   �      D  , ,  �   #  �   �  Ȗ  �  Ȗ  #  �   #      D  , ,  �   �  �   y  Ȗ  y  Ȗ  �  �   �      D  , ,  �   �  �   9  Ȗ  9  Ȗ  �  �   �      D  , ,  �   w  �     Ȗ    Ȗ  w  �   w      D  , ,  �   c  �   �  Ȗ  �  Ȗ  c  �   c      D  , ,  �    #  �    �  Ȗ   �  Ȗ   #  �    #      D  , ,  � ����  � ���y  Ȗ���y  Ȗ����  � ����      D  , ,  � ����  � ���9  Ȗ���9  Ȗ����  � ����      D  , ,  � ���c  � ����  Ȗ����  Ȗ���c  � ���c      D  , ,  �   7  �   �  Ȗ  �  Ȗ  7  �   7      D  , ,  �D  7  �D  �  ��  �  ��  7  �D  7      D  , ,  ̜  7  ̜  �  �2  �  �2  7  ̜  7      D  , ,  ��  7  ��  �  �v  �  �v  7  ��  7      D  , ,  �8  7  �8  �  ��  �  ��  7  �8  7      D  , ,  �8  �  �8  �  ��  �  ��  �  �8  �      D  , ,  �D  �  �D  �  ��  �  ��  �  �D  �      D  , ,  ̜  �  ̜  �  �2  �  �2  �  ̜  �      D  , ,  ��  �  ��  �  �v  �  �v  �  ��  �      D  , ,  �8  �  �8  �  ��  �  ��  �  �8  �      D  , ,  �D  �  �D  �  ��  �  ��  �  �D  �      D  , ,  �D  �  �D  M  ��  M  ��  �  �D  �      D  , ,  ̜  �  ̜  M  �2  M  �2  �  ̜  �      D  , ,  ��  �  ��  M  �v  M  �v  �  ��  �      D  , ,  �8  �  �8  M  ��  M  ��  �  �8  �      D  , ,  �'  	�  �'  
#  ɽ  
#  ɽ  	�  �'  	�      D  , ,  �u  	�  �u  
#  �  
#  �  	�  �u  	�      D  , ,  ��  	�  ��  
#  �Y  
#  �Y  	�  ��  	�      D  , ,  �  	�  �  
#  Ч  
#  Ч  	�  �  	�      D  , ,  �'  M  �'  �  ɽ  �  ɽ  M  �'  M      D  , ,  �u  M  �u  �  �  �  �  M  �u  M      D  , ,  ��  M  ��  �  �Y  �  �Y  M  ��  M      D  , ,  �  M  �  �  Ч  �  Ч  M  �  M      D  , ,  �D  �  �D  M  ��  M  ��  �  �D  �      D  , ,  ̜  �  ̜  M  �2  M  �2  �  ̜  �      D  , ,  ��  �  ��  M  �v  M  �v  �  ��  �      D  , ,  �8  �  �8  M  ��  M  ��  �  �8  �      D  , ,  ̜  �  ̜  �  �2  �  �2  �  ̜  �      D  , ,  �D  w  �D    ��    ��  w  �D  w      D  , ,  �D  w  �D    ��    ��  w  �D  w      D  , ,  ̜  w  ̜    �2    �2  w  ̜  w      D  , ,  ̜  w  ̜    �2    �2  w  ̜  w      D  , ,  ��  w  ��    �v    �v  w  ��  w      D  , ,  ��  w  ��    �v    �v  w  ��  w      D  , ,  �8  w  �8    ��    ��  w  �8  w      D  , ,  �8  w  �8    ��    ��  w  �8  w      D  , ,  ��  �  ��  �  �v  �  �v  �  ��  �      D  , ,  �D  7  �D  �  ��  �  ��  7  �D  7      D  , ,  ̜  7  ̜  �  �2  �  �2  7  ̜  7      D  , ,  ��  7  ��  �  �v  �  �v  7  ��  7      D  , ,  �8  7  �8  �  ��  �  ��  7  �8  7      D  , ,  �S  	�  �S  
#  ��  
#  ��  	�  �S  	�      D  , ,  �S  M  �S  �  ��  �  ��  M  �S  M      D  , ,  ��  7  ��  �  ��  �  ��  7  ��  7      D  , ,  �8  7  �8  �  ��  �  ��  7  �8  7      D  , ,  ��  7  ��  �  �&  �  �&  7  ��  7      D  , ,  ��  7  ��  �  �j  �  �j  7  ��  7      D  , ,  �,  7  �,  �  ��  �  ��  7  �,  7      D  , ,  �p  7  �p  �  �  �  �  7  �p  7      D  , ,  ��  7  ��  �  �^  �  �^  7  ��  7      D  , ,  �  7  �  �  ��  �  ��  7  �  7      D  , ,  �d  7  �d  �  ��  �  ��  7  �d  7      D  , ,  Ũ  7  Ũ  �  �>  �  �>  7  Ũ  7      D  , ,  ��  w  ��    �^    �^  w  ��  w      D  , ,  �d  �  �d  M  ��  M  ��  �  �d  �      D  , ,  �  w  �    ��    ��  w  �  w      D  , ,  �d  w  �d    ��    ��  w  �d  w      D  , ,  Ũ  w  Ũ    �>    �>  w  Ũ  w      D  , ,  �  w  �    ��    ��  w  �  w      D  , ,  �d  w  �d    ��    ��  w  �d  w      D  , ,  Ũ  w  Ũ    �>    �>  w  Ũ  w      D  , ,  �p  w  �p    �    �  w  �p  w      D  , ,  Ũ  �  Ũ  M  �>  M  �>  �  Ũ  �      D  , ,  �p  �  �p  �  �  �  �  �  �p  �      D  , ,  ��  �  ��  �  �^  �  �^  �  ��  �      D  , ,  �  �  �  �  ��  �  ��  �  �  �      D  , ,  �d  �  �d  �  ��  �  ��  �  �d  �      D  , ,  ��  w  ��    �^    �^  w  ��  w      D  , ,  Ũ  �  Ũ  �  �>  �  �>  �  Ũ  �      D  , ,  �p  7  �p  �  �  �  �  7  �p  7      D  , ,  ��  7  ��  �  �^  �  �^  7  ��  7      D  , ,  �  7  �  �  ��  �  ��  7  �  7      D  , ,  �d  7  �d  �  ��  �  ��  7  �d  7      D  , ,  Ũ  7  Ũ  �  �>  �  �>  7  Ũ  7      D  , ,  �  �  �  M  ��  M  ��  �  �  �      D  , ,  �p  w  �p    �    �  w  �p  w      D  , ,  �p  �  �p  M  �  M  �  �  �p  �      D  , ,  ��  �  ��  M  �^  M  �^  �  ��  �      D  , ,  ��  �  ��  M  ��  M  ��  �  ��  �      D  , ,  �8  w  �8    ��    ��  w  �8  w      D  , ,  �8  �  �8  M  ��  M  ��  �  �8  �      D  , ,  ��  w  ��    ��    ��  w  ��  w      D  , ,  ��  7  ��  �  ��  �  ��  7  ��  7      D  , ,  �8  7  �8  �  ��  �  ��  7  �8  7      D  , ,  ��  7  ��  �  �&  �  �&  7  ��  7      D  , ,  ��  7  ��  �  �j  �  �j  7  ��  7      D  , ,  �,  7  �,  �  ��  �  ��  7  �,  7      D  , ,  ��  w  ��    �&    �&  w  ��  w      D  , ,  ��  �  ��  M  �&  M  �&  �  ��  �      D  , ,  ��  �  ��  M  �j  M  �j  �  ��  �      D  , ,  �,  w  �,    ��    ��  w  �,  w      D  , ,  ��  w  ��    �j    �j  w  ��  w      D  , ,  ��  w  ��    �j    �j  w  ��  w      D  , ,  �,  w  �,    ��    ��  w  �,  w      D  , ,  �,  �  �,  M  ��  M  ��  �  �,  �      D  , ,  ��  w  ��    �&    �&  w  ��  w      D  , ,  ��  w  ��    ��    ��  w  ��  w      D  , ,  �8  w  �8    ��    ��  w  �8  w      D  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      D  , ,  �8  �  �8  �  ��  �  ��  �  �8  �      D  , ,  ��  �  ��  �  �&  �  �&  �  ��  �      D  , ,  ��  �  ��  �  �j  �  �j  �  ��  �      D  , ,  �,  �  �,  �  ��  �  ��  �  �,  �      D  , ,  �,  �  �,  �  ��  �  ��  �  �,  �      D  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      D  , ,  ��  	�  ��  
#  �c  
#  �c  	�  ��  	�      D  , ,  �  	�  �  
#  ��  
#  ��  	�  �  	�      D  , ,  �i  	�  �i  
#  ��  
#  ��  	�  �i  	�      D  , ,  ��  	�  ��  
#  �M  
#  �M  	�  ��  	�      D  , ,  �  	�  �  
#  ��  
#  ��  	�  �  	�      D  , ,  ��  �  ��  M  ��  M  ��  �  ��  �      D  , ,  �8  �  �8  M  ��  M  ��  �  �8  �      D  , ,  ��  �  ��  M  �&  M  �&  �  ��  �      D  , ,  ��  �  ��  M  �j  M  �j  �  ��  �      D  , ,  �,  �  �,  M  ��  M  ��  �  �,  �      D  , ,  ��  M  ��  �  �c  �  �c  M  ��  M      D  , ,  �  M  �  �  ��  �  ��  M  �  M      D  , ,  �i  M  �i  �  ��  �  ��  M  �i  M      D  , ,  ��  M  ��  �  �M  �  �M  M  ��  M      D  , ,  �  M  �  �  ��  �  ��  M  �  M      D  , ,  �8  �  �8  �  ��  �  ��  �  �8  �      D  , ,  ��  �  ��  �  �&  �  �&  �  ��  �      D  , ,  ��  �  ��  �  �j  �  �j  �  ��  �      D  , ,  �=  	�  �=  
#  ��  
#  ��  	�  �=  	�      D  , ,  ċ  	�  ċ  
#  �!  
#  �!  	�  ċ  	�      D  , ,  ��  	�  ��  
#  �o  
#  �o  	�  ��  	�      D  , ,  �  �  �  �  ��  �  ��  �  �  �      D  , ,  �d  �  �d  �  ��  �  ��  �  �d  �      D  , ,  Ũ  �  Ũ  �  �>  �  �>  �  Ũ  �      D  , ,  �p  �  �p  �  �  �  �  �  �p  �      D  , ,  �p  �  �p  M  �  M  �  �  �p  �      D  , ,  ��  �  ��  M  �^  M  �^  �  ��  �      D  , ,  �  �  �  M  ��  M  ��  �  �  �      D  , ,  �d  �  �d  M  ��  M  ��  �  �d  �      D  , ,  Ũ  �  Ũ  M  �>  M  �>  �  Ũ  �      D  , ,  ��  �  ��  �  �^  �  �^  �  ��  �      D  , ,  ��  M  ��  �  �7  �  �7  M  ��  M      D  , ,  ��  M  ��  �  ��  �  ��  M  ��  M      D  , ,  �=  M  �=  �  ��  �  ��  M  �=  M      D  , ,  ċ  M  ċ  �  �!  �  �!  M  ċ  M      D  , ,  ��  M  ��  �  �o  �  �o  M  ��  M      D  , ,  ��  	�  ��  
#  �7  
#  �7  	�  ��  	�      D  , ,  ��  	�  ��  
#  ��  
#  ��  	�  ��  	�      D  , ,  �8  c  �8  �  ��  �  ��  c  �8  c      D  , ,  ��  c  ��  �  �&  �  �&  c  ��  c      D  , ,  ��  c  ��  �  �j  �  �j  c  ��  c      D  , ,  �,  c  �,  �  ��  �  ��  c  �,  c      D  , ,  �p  c  �p  �  �  �  �  c  �p  c      D  , ,  ��  c  ��  �  �^  �  �^  c  ��  c      D  , ,  �  c  �  �  ��  �  ��  c  �  c      D  , ,  �d  c  �d  �  ��  �  ��  c  �d  c      D  , ,  Ũ  c  Ũ  �  �>  �  �>  c  Ũ  c      D  , ,  ��  #  ��  �  �^  �  �^  #  ��  #      D  , ,  �  #  �  �  ��  �  ��  #  �  #      D  , ,  ��   #  ��   �  ��   �  ��   #  ��   #      D  , ,  �8   #  �8   �  ��   �  ��   #  �8   #      D  , ,  ��   #  ��   �  �&   �  �&   #  ��   #      D  , ,  ��   #  ��   �  �j   �  �j   #  ��   #      D  , ,  �,   #  �,   �  ��   �  ��   #  �,   #      D  , ,  �p   #  �p   �  �   �  �   #  �p   #      D  , ,  ��   #  ��   �  �^   �  �^   #  ��   #      D  , ,  �   #  �   �  ��   �  ��   #  �   #      D  , ,  �d   #  �d   �  ��   �  ��   #  �d   #      D  , ,  Ũ   #  Ũ   �  �>   �  �>   #  Ũ   #      D  , ,  �d  #  �d  �  ��  �  ��  #  �d  #      D  , ,  Ũ  #  Ũ  �  �>  �  �>  #  Ũ  #      D  , ,  ������  �����y  �����y  ������  ������      D  , ,  �8����  �8���y  �����y  ������  �8����      D  , ,  ������  �����y  �&���y  �&����  ������      D  , ,  ������  �����y  �j���y  �j����  ������      D  , ,  �,����  �,���y  �����y  ������  �,����      D  , ,  �p����  �p���y  ����y  �����  �p����      D  , ,  ������  �����y  �^���y  �^����  ������      D  , ,  �����  ����y  �����y  ������  �����      D  , ,  �d����  �d���y  �����y  ������  �d����      D  , ,  Ũ����  Ũ���y  �>���y  �>����  Ũ����      D  , ,  ��  #  ��  �  ��  �  ��  #  ��  #      D  , ,  �8  #  �8  �  ��  �  ��  #  �8  #      D  , ,  ������  �����9  �����9  ������  ������      D  , ,  �8����  �8���9  �����9  ������  �8����      D  , ,  ������  �����9  �&���9  �&����  ������      D  , ,  ������  �����9  �j���9  �j����  ������      D  , ,  �,����  �,���9  �����9  ������  �,����      D  , ,  �p����  �p���9  ����9  �����  �p����      D  , ,  ������  �����9  �^���9  �^����  ������      D  , ,  �����  ����9  �����9  ������  �����      D  , ,  �d����  �d���9  �����9  ������  �d����      D  , ,  Ũ����  Ũ���9  �>���9  �>����  Ũ����      D  , ,  ��  �  ��  y  ��  y  ��  �  ��  �      D  , ,  �8  �  �8  y  ��  y  ��  �  �8  �      D  , ,  �����c  ������  ������  �����c  �����c      D  , ,  �8���c  �8����  ������  �����c  �8���c      D  , ,  �����c  ������  �&����  �&���c  �����c      D  , ,  �����c  ������  �j����  �j���c  �����c      D  , ,  �,���c  �,����  ������  �����c  �,���c      D  , ,  �p���c  �p����  �����  ����c  �p���c      D  , ,  �����c  ������  �^����  �^���c  �����c      D  , ,  ����c  �����  ������  �����c  ����c      D  , ,  �d���c  �d����  ������  �����c  �d���c      D  , ,  Ũ���c  Ũ����  �>����  �>���c  Ũ���c      D  , ,  ��  �  ��  y  �&  y  �&  �  ��  �      D  , ,  ��  �  ��  y  �j  y  �j  �  ��  �      D  , ,  �,  �  �,  y  ��  y  ��  �  �,  �      D  , ,  �p  �  �p  y  �  y  �  �  �p  �      D  , ,  ��  �  ��  y  �^  y  �^  �  ��  �      D  , ,  �  �  �  y  ��  y  ��  �  �  �      D  , ,  �d  �  �d  y  ��  y  ��  �  �d  �      D  , ,  Ũ  �  Ũ  y  �>  y  �>  �  Ũ  �      D  , ,  ��  #  ��  �  �&  �  �&  #  ��  #      D  , ,  ��  #  ��  �  �j  �  �j  #  ��  #      D  , ,  ��  �  ��  9  ��  9  ��  �  ��  �      D  , ,  �8  �  �8  9  ��  9  ��  �  �8  �      D  , ,  ��  �  ��  9  �&  9  �&  �  ��  �      D  , ,  ��  �  ��  9  �j  9  �j  �  ��  �      D  , ,  �,  �  �,  9  ��  9  ��  �  �,  �      D  , ,  �p  �  �p  9  �  9  �  �  �p  �      D  , ,  ��  �  ��  9  �^  9  �^  �  ��  �      D  , ,  �  �  �  9  ��  9  ��  �  �  �      D  , ,  �d  �  �d  9  ��  9  ��  �  �d  �      D  , ,  Ũ  �  Ũ  9  �>  9  �>  �  Ũ  �      D  , ,  �,  #  �,  �  ��  �  ��  #  �,  #      D  , ,  �p  #  �p  �  �  �  �  #  �p  #      D  , ,  ��  c  ��  �  ��  �  ��  c  ��  c      D  , ,  ��  #  ��  �  �v  �  �v  #  ��  #      D  , ,  �8  #  �8  �  ��  �  ��  #  �8  #      D  , ,  �D����  �D���y  �����y  ������  �D����      D  , ,  ̜����  ̜���y  �2���y  �2����  ̜����      D  , ,  ������  �����y  �v���y  �v����  ������      D  , ,  �8����  �8���y  �����y  ������  �8����      D  , ,  �D���c  �D����  ������  �����c  �D���c      D  , ,  ̜���c  ̜����  �2����  �2���c  ̜���c      D  , ,  �����c  ������  �v����  �v���c  �����c      D  , ,  �8���c  �8����  ������  �����c  �8���c      D  , ,  �D  �  �D  9  ��  9  ��  �  �D  �      D  , ,  ̜  �  ̜  9  �2  9  �2  �  ̜  �      D  , ,  ��  �  ��  9  �v  9  �v  �  ��  �      D  , ,  �8  �  �8  9  ��  9  ��  �  �8  �      D  , ,  �D   #  �D   �  ��   �  ��   #  �D   #      D  , ,  ̜   #  ̜   �  �2   �  �2   #  ̜   #      D  , ,  ��   #  ��   �  �v   �  �v   #  ��   #      D  , ,  �8   #  �8   �  ��   �  ��   #  �8   #      D  , ,  �D  c  �D  �  ��  �  ��  c  �D  c      D  , ,  ̜  c  ̜  �  �2  �  �2  c  ̜  c      D  , ,  ��  c  ��  �  �v  �  �v  c  ��  c      D  , ,  �8  c  �8  �  ��  �  ��  c  �8  c      D  , ,  �D����  �D���9  �����9  ������  �D����      D  , ,  ̜����  ̜���9  �2���9  �2����  ̜����      D  , ,  ������  �����9  �v���9  �v����  ������      D  , ,  �8����  �8���9  �����9  ������  �8����      D  , ,  �D  �  �D  y  ��  y  ��  �  �D  �      D  , ,  ̜  �  ̜  y  �2  y  �2  �  ̜  �      D  , ,  ��  �  ��  y  �v  y  �v  �  ��  �      D  , ,  �8  �  �8  y  ��  y  ��  �  �8  �      D  , ,  �D  #  �D  �  ��  �  ��  #  �D  #      D  , ,  ̜  #  ̜  �  �2  �  �2  #  ̜  #      D  , ,  ��  �  ��    �F    �F  �  ��  �      D  , ,  �L  �  �L    ��    ��  �  �L  �      D  , ,  ��  �  ��    �~    �~  �  ��  �      D  , ,  ~@  I  ~@  �  ~�  �  ~�  I  ~@  I      D  , ,  �)  &�  �)  'Q  ��  'Q  ��  &�  �)  &�      D  , ,  �w  &�  �w  'Q  �  'Q  �  &�  �w  &�      D  , ,  ��  &�  ��  'Q  �[  'Q  �[  &�  ��  &�      D  , ,  �  &�  �  'Q  ��  'Q  ��  &�  �  &�      D  , ,  �a  &�  �a  'Q  ��  'Q  ��  &�  �a  &�      D  , ,  ��  &�  ��  'Q  �E  'Q  �E  &�  ��  &�      D  , ,  ��  &�  ��  'Q  ��  'Q  ��  &�  ��  &�      D  , ,  �K  &�  �K  'Q  ��  'Q  ��  &�  �K  &�      D  , ,  ��  &�  ��  'Q  �/  'Q  �/  &�  ��  &�      D  , ,  ~@  �  ~@  _  ~�  _  ~�  �  ~@  �      D  , ,  ��  �  ��  _  �r  _  �r  �  ��  �      D  , ,  �x  �  �x  _  �  _  �  �  �x  �      D  , ,  �  �  �  _  ��  _  ��  �  �  �      D  , ,  ��  �  ��  _  �F  _  �F  �  ��  �      D  , ,  �L  �  �L  _  ��  _  ��  �  �L  �      D  , ,  ��  �  ��  _  �~  _  �~  �  ��  �      D  , ,  ��  �  ��  _  �  _  �  �  ��  �      D  , ,  �   �  �   _  ��  _  ��  �  �   �      D  , ,  ��  �  ��  _  �R  _  �R  �  ��  �      D  , ,  ~@  	  ~@  �  ~�  �  ~�  	  ~@  	      D  , ,  ��  	  ��  �  �r  �  �r  	  ��  	      D  , ,  �x  	  �x  �  �  �  �  	  �x  	      D  , ,  �  	  �  �  ��  �  ��  	  �  	      D  , ,  ��  	  ��  �  �F  �  �F  	  ��  	      D  , ,  �L  	  �L  �  ��  �  ��  	  �L  	      D  , ,  ��  	  ��  �  �~  �  �~  	  ��  	      D  , ,  ��  	  ��  �  �  �  �  	  ��  	      D  , ,  �   	  �   �  ��  �  ��  	  �   	      D  , ,  ��  	  ��  �  �R  �  �R  	  ��  	      D  , ,  �X  	  �X  �  ��  �  ��  	  �X  	      D  , ,  ��  I  ��  �  �r  �  �r  I  ��  I      D  , ,  �x  I  �x  �  �  �  �  I  �x  I      D  , ,  �  I  �  �  ��  �  ��  I  �  I      D  , ,  ��  I  ��  �  �F  �  �F  I  ��  I      D  , ,  �L  I  �L  �  ��  �  ��  I  �L  I      D  , ,  ��  I  ��  �  �~  �  �~  I  ��  I      D  , ,  ��  I  ��  �  �  �  �  I  ��  I      D  , ,  �   I  �   �  ��  �  ��  I  �   I      D  , ,  ��  I  ��  �  �R  �  �R  I  ��  I      D  , ,  �X  I  �X  �  ��  �  ��  I  �X  I      D  , ,  ��  &�  ��  'Q  �}  'Q  �}  &�  ��  &�      D  , ,  �5  &�  �5  'Q  ��  'Q  ��  &�  �5  &�      D  , ,  ��  &�  ��  'Q  �  'Q  �  &�  ��  &�      D  , ,  ��  &�  ��  'Q  �g  'Q  �g  &�  ��  &�      D  , ,  �  &�  �  'Q  ��  'Q  ��  &�  �  &�      D  , ,  �m  &�  �m  'Q  �  'Q  �  &�  �m  &�      D  , ,  �/  &�  �/  'Q  ��  'Q  ��  &�  �/  &�      D  , ,  �}  &�  �}  'Q  �  'Q  �  &�  �}  &�      D  , ,  ��  &�  ��  'Q  �a  'Q  �a  &�  ��  &�      D  , ,  ��  �  ��    �    �  �  ��  �      D  , ,  �   �  �     ��    ��  �  �   �      D  , ,  ��  �  ��    �R    �R  �  ��  �      D  , ,  �X  �  �X    ��    ��  �  �X  �      D  , ,  ~@  �  ~@    ~�    ~�  �  ~@  �      D  , ,  ��  �  ��    �r    �r  �  ��  �      D  , ,  �x  �  �x    �    �  �  �x  �      D  , ,  �X  �  �X  _  ��  _  ��  �  �X  �      D  , ,  �  �  �    ��    ��  �  �  �      D  , ,  u�  &�  u�  'Q  va  'Q  va  &�  u�  &�      D  , ,  x  &�  x  'Q  x�  'Q  x�  &�  x  &�      D  , ,  ]�  	  ]�  �  ^�  �  ^�  	  ]�  	      D  , ,  b�  	  b�  �  c.  �  c.  	  b�  	      D  , ,  Z#  &�  Z#  'Q  Z�  'Q  Z�  &�  Z#  &�      D  , ,  \q  &�  \q  'Q  ]  'Q  ]  &�  \q  &�      D  , ,  ^�  &�  ^�  'Q  _U  'Q  _U  &�  ^�  &�      D  , ,  a  &�  a  'Q  a�  'Q  a�  &�  a  &�      D  , ,  c[  &�  c[  'Q  c�  'Q  c�  &�  c[  &�      D  , ,  e�  &�  e�  'Q  f?  'Q  f?  &�  e�  &�      D  , ,  g�  &�  g�  'Q  h�  'Q  h�  &�  g�  &�      D  , ,  jE  &�  jE  'Q  j�  'Q  j�  &�  jE  &�      D  , ,  l�  &�  l�  'Q  m)  'Q  m)  &�  l�  &�      D  , ,  n�  &�  n�  'Q  ow  'Q  ow  &�  n�  &�      D  , ,  q/  &�  q/  'Q  q�  'Q  q�  &�  q/  &�      D  , ,  s}  &�  s}  'Q  t  'Q  t  &�  s}  &�      D  , ,  g4  	  g4  �  g�  �  g�  	  g4  	      D  , ,  k�  	  k�  �  lf  �  lf  	  k�  	      D  , ,  pl  	  pl  �  q  �  q  	  pl  	      D  , ,  u  	  u  �  u�  �  u�  	  u  	      D  , ,  y�  	  y�  �  z:  �  z:  	  y�  	      D  , ,  ]�  �  ]�  _  ^�  _  ^�  �  ]�  �      D  , ,  b�  �  b�  _  c.  _  c.  �  b�  �      D  , ,  g4  �  g4  _  g�  _  g�  �  g4  �      D  , ,  k�  �  k�  _  lf  _  lf  �  k�  �      D  , ,  pl  �  pl  _  q  _  q  �  pl  �      D  , ,  u  �  u  _  u�  _  u�  �  u  �      D  , ,  y�  �  y�  _  z:  _  z:  �  y�  �      D  , ,  zg  &�  zg  'Q  z�  'Q  z�  &�  zg  &�      D  , ,  b�  I  b�  �  c.  �  c.  I  b�  I      D  , ,  g4  I  g4  �  g�  �  g�  I  g4  I      D  , ,  ]�  �  ]�    ^�    ^�  �  ]�  �      D  , ,  b�  �  b�    c.    c.  �  b�  �      D  , ,  g4  �  g4    g�    g�  �  g4  �      D  , ,  k�  �  k�    lf    lf  �  k�  �      D  , ,  pl  �  pl    q    q  �  pl  �      D  , ,  u  �  u    u�    u�  �  u  �      D  , ,  y�  �  y�    z:    z:  �  y�  �      D  , ,  k�  I  k�  �  lf  �  lf  I  k�  I      D  , ,  pl  I  pl  �  q  �  q  I  pl  I      D  , ,  u  I  u  �  u�  �  u�  I  u  I      D  , ,  y�  I  y�  �  z:  �  z:  I  y�  I      D  , ,  ]�  I  ]�  �  ^�  �  ^�  I  ]�  I      D  , ,  c�  	�  c�  
#  dU  
#  dU  	�  c�  	�      D  , ,  c�  M  c�  �  dU  �  dU  M  c�  M      D  , ,  u  7  u  �  u�  �  u�  7  u  7      D  , ,  wL  7  wL  �  w�  �  w�  7  wL  7      D  , ,  y�  7  y�  �  z:  �  z:  7  y�  7      D  , ,  {�  7  {�  �  |~  �  |~  7  {�  7      D  , ,  pl  w  pl    q    q  w  pl  w      D  , ,  pl  7  pl  �  q  �  q  7  pl  7      D  , ,  pl  �  pl  �  q  �  q  �  pl  �      D  , ,  pl  �  pl  �  q  �  q  �  pl  �      D  , ,  d�  7  d�  �  er  �  er  7  d�  7      D  , ,  g4  7  g4  �  g�  �  g�  7  g4  7      D  , ,  ix  7  ix  �  j  �  j  7  ix  7      D  , ,  k�  7  k�  �  lf  �  lf  7  k�  7      D  , ,  n  7  n  �  n�  �  n�  7  n  7      D  , ,  pl  7  pl  �  q  �  q  7  pl  7      D  , ,  r�  7  r�  �  sF  �  sF  7  r�  7      D  , ,  pl  �  pl  M  q  M  q  �  pl  �      D  , ,  pl  �  pl  M  q  M  q  �  pl  �      D  , ,  pl  w  pl    q    q  w  pl  w      D  , ,  wL  7  wL  �  w�  �  w�  7  wL  7      D  , ,  y�  7  y�  �  z:  �  z:  7  y�  7      D  , ,  {�  7  {�  �  |~  �  |~  7  {�  7      D  , ,  {�  w  {�    |~    |~  w  {�  w      D  , ,  r�  w  r�    sF    sF  w  r�  w      D  , ,  r�  �  r�  �  sF  �  sF  �  r�  �      D  , ,  u  �  u  �  u�  �  u�  �  u  �      D  , ,  wL  �  wL  �  w�  �  w�  �  wL  �      D  , ,  y�  �  y�  �  z:  �  z:  �  y�  �      D  , ,  {�  �  {�  �  |~  �  |~  �  {�  �      D  , ,  u  w  u    u�    u�  w  u  w      D  , ,  wL  w  wL    w�    w�  w  wL  w      D  , ,  r�  w  r�    sF    sF  w  r�  w      D  , ,  u  w  u    u�    u�  w  u  w      D  , ,  wL  w  wL    w�    w�  w  wL  w      D  , ,  y�  w  y�    z:    z:  w  y�  w      D  , ,  {�  w  {�    |~    |~  w  {�  w      D  , ,  y�  w  y�    z:    z:  w  y�  w      D  , ,  r�  �  r�  M  sF  M  sF  �  r�  �      D  , ,  u  �  u  M  u�  M  u�  �  u  �      D  , ,  wL  �  wL  M  w�  M  w�  �  wL  �      D  , ,  y�  �  y�  M  z:  M  z:  �  y�  �      D  , ,  {�  �  {�  M  |~  M  |~  �  {�  �      D  , ,  r�  7  r�  �  sF  �  sF  7  r�  7      D  , ,  u  7  u  �  u�  �  u�  7  u  7      D  , ,  n  w  n    n�    n�  w  n  w      D  , ,  d�  w  d�    er    er  w  d�  w      D  , ,  d�  7  d�  �  er  �  er  7  d�  7      D  , ,  g4  7  g4  �  g�  �  g�  7  g4  7      D  , ,  d�  �  d�  �  er  �  er  �  d�  �      D  , ,  g4  �  g4  �  g�  �  g�  �  g4  �      D  , ,  ix  �  ix  �  j  �  j  �  ix  �      D  , ,  d�  w  d�    er    er  w  d�  w      D  , ,  g4  w  g4    g�    g�  w  g4  w      D  , ,  ix  w  ix    j    j  w  ix  w      D  , ,  d�  �  d�  M  er  M  er  �  d�  �      D  , ,  g4  �  g4  M  g�  M  g�  �  g4  �      D  , ,  ix  �  ix  M  j  M  j  �  ix  �      D  , ,  k�  �  k�  M  lf  M  lf  �  k�  �      D  , ,  n  �  n  M  n�  M  n�  �  n  �      D  , ,  k�  �  k�  �  lf  �  lf  �  k�  �      D  , ,  n  �  n  �  n�  �  n�  �  n  �      D  , ,  ix  7  ix  �  j  �  j  7  ix  7      D  , ,  k�  7  k�  �  lf  �  lf  7  k�  7      D  , ,  n  7  n  �  n�  �  n�  7  n  7      D  , ,  g4  w  g4    g�    g�  w  g4  w      D  , ,  k�  w  k�    lf    lf  w  k�  w      D  , ,  n  w  n    n�    n�  w  n  w      D  , ,  ix  w  ix    j    j  w  ix  w      D  , ,  k�  w  k�    lf    lf  w  k�  w      D  , ,  oE  M  oE  �  o�  �  o�  M  oE  M      D  , ,  f  	�  f  
#  f�  
#  f�  	�  f  	�      D  , ,  h[  	�  h[  
#  h�  
#  h�  	�  h[  	�      D  , ,  d�  �  d�  �  er  �  er  �  d�  �      D  , ,  g4  �  g4  �  g�  �  g�  �  g4  �      D  , ,  ix  �  ix  �  j  �  j  �  ix  �      D  , ,  k�  �  k�  �  lf  �  lf  �  k�  �      D  , ,  n  �  n  �  n�  �  n�  �  n  �      D  , ,  j�  	�  j�  
#  k?  
#  k?  	�  j�  	�      D  , ,  l�  	�  l�  
#  m�  
#  m�  	�  l�  	�      D  , ,  oE  	�  oE  
#  o�  
#  o�  	�  oE  	�      D  , ,  f  M  f  �  f�  �  f�  M  f  M      D  , ,  h[  M  h[  �  h�  �  h�  M  h[  M      D  , ,  d�  �  d�  M  er  M  er  �  d�  �      D  , ,  g4  �  g4  M  g�  M  g�  �  g4  �      D  , ,  ix  �  ix  M  j  M  j  �  ix  �      D  , ,  k�  �  k�  M  lf  M  lf  �  k�  �      D  , ,  n  �  n  M  n�  M  n�  �  n  �      D  , ,  j�  M  j�  �  k?  �  k?  M  j�  M      D  , ,  l�  M  l�  �  m�  �  m�  M  l�  M      D  , ,  u  �  u  �  u�  �  u�  �  u  �      D  , ,  wL  �  wL  �  w�  �  w�  �  wL  �      D  , ,  x}  M  x}  �  y  �  y  M  x}  M      D  , ,  z�  M  z�  �  {a  �  {a  M  z�  M      D  , ,  q�  	�  q�  
#  r)  
#  r)  	�  q�  	�      D  , ,  s�  	�  s�  
#  tw  
#  tw  	�  s�  	�      D  , ,  v/  	�  v/  
#  v�  
#  v�  	�  v/  	�      D  , ,  x}  	�  x}  
#  y  
#  y  	�  x}  	�      D  , ,  z�  	�  z�  
#  {a  
#  {a  	�  z�  	�      D  , ,  q�  M  q�  �  r)  �  r)  M  q�  M      D  , ,  s�  M  s�  �  tw  �  tw  M  s�  M      D  , ,  v/  M  v/  �  v�  �  v�  M  v/  M      D  , ,  r�  �  r�  �  sF  �  sF  �  r�  �      D  , ,  y�  �  y�  �  z:  �  z:  �  y�  �      D  , ,  r�  �  r�  M  sF  M  sF  �  r�  �      D  , ,  u  �  u  M  u�  M  u�  �  u  �      D  , ,  wL  �  wL  M  w�  M  w�  �  wL  �      D  , ,  y�  �  y�  M  z:  M  z:  �  y�  �      D  , ,  {�  �  {�  M  |~  M  |~  �  {�  �      D  , ,  {�  �  {�  �  |~  �  |~  �  {�  �      D  , ,  b�  �  b�  �  c.  �  c.  �  b�  �      D  , ,  b�  w  b�    c.    c.  w  b�  w      D  , ,  aq  M  aq  �  b  �  b  M  aq  M      D  , ,  ]�  7  ]�  �  ^�  �  ^�  7  ]�  7      D  , ,  `@  7  `@  �  `�  �  `�  7  `@  7      D  , ,  b�  7  b�  �  c.  �  c.  7  b�  7      D  , ,  aq  	�  aq  
#  b  
#  b  	�  aq  	�      D  , ,  _#  	�  _#  
#  _�  
#  _�  	�  _#  	�      D  , ,  b�  7  b�  �  c.  �  c.  7  b�  7      D  , ,  _#  M  _#  �  _�  �  _�  M  _#  M      D  , ,  ]�  w  ]�    ^�    ^�  w  ]�  w      D  , ,  ]�  �  ]�  �  ^�  �  ^�  �  ]�  �      D  , ,  `@  �  `@  �  `�  �  `�  �  `@  �      D  , ,  ]�  �  ]�  M  ^�  M  ^�  �  ]�  �      D  , ,  `@  �  `@  M  `�  M  `�  �  `@  �      D  , ,  b�  �  b�  M  c.  M  c.  �  b�  �      D  , ,  b�  �  b�  �  c.  �  c.  �  b�  �      D  , ,  `@  w  `@    `�    `�  w  `@  w      D  , ,  ]�  7  ]�  �  ^�  �  ^�  7  ]�  7      D  , ,  ]�  w  ]�    ^�    ^�  w  ]�  w      D  , ,  `@  w  `@    `�    `�  w  `@  w      D  , ,  b�  w  b�    c.    c.  w  b�  w      D  , ,  `@  7  `@  �  `�  �  `�  7  `@  7      D  , ,  ]�  �  ]�  �  ^�  �  ^�  �  ]�  �      D  , ,  `@  �  `@  �  `�  �  `�  �  `@  �      D  , ,  ]�  �  ]�  M  ^�  M  ^�  �  ]�  �      D  , ,  `@  �  `@  M  `�  M  `�  �  `@  �      D  , ,  b�  �  b�  M  c.  M  c.  �  b�  �      D  , ,  `@  c  `@  �  `�  �  `�  c  `@  c      D  , ,  b�  c  b�  �  c.  �  c.  c  b�  c      D  , ,  `@  �  `@  9  `�  9  `�  �  `@  �      D  , ,  ]����c  ]�����  ^�����  ^����c  ]����c      D  , ,  `@���c  `@����  `�����  `����c  `@���c      D  , ,  b����c  b�����  c.����  c.���c  b����c      D  , ,  b�  �  b�  9  c.  9  c.  �  b�  �      D  , ,  ]�   #  ]�   �  ^�   �  ^�   #  ]�   #      D  , ,  ]�����  ]����9  ^����9  ^�����  ]�����      D  , ,  `@����  `@���9  `����9  `�����  `@����      D  , ,  b�����  b����9  c.���9  c.����  b�����      D  , ,  `@   #  `@   �  `�   �  `�   #  `@   #      D  , ,  b�   #  b�   �  c.   �  c.   #  b�   #      D  , ,  ]�����  ]����y  ^����y  ^�����  ]�����      D  , ,  `@����  `@���y  `����y  `�����  `@����      D  , ,  b�����  b����y  c.���y  c.����  b�����      D  , ,  b�  #  b�  �  c.  �  c.  #  b�  #      D  , ,  ]�  #  ]�  �  ^�  �  ^�  #  ]�  #      D  , ,  `@  #  `@  �  `�  �  `�  #  `@  #      D  , ,  ]�  �  ]�  y  ^�  y  ^�  �  ]�  �      D  , ,  `@  �  `@  y  `�  y  `�  �  `@  �      D  , ,  b�  �  b�  y  c.  y  c.  �  b�  �      D  , ,  ]�  �  ]�  9  ^�  9  ^�  �  ]�  �      D  , ,  ]�  c  ]�  �  ^�  �  ^�  c  ]�  c      D  , ,  {�  #  {�  �  |~  �  |~  #  {�  #      D  , ,  d�  #  d�  �  er  �  er  #  d�  #      D  , ,  d�����  d����y  er���y  er����  d�����      D  , ,  g4����  g4���y  g����y  g�����  g4����      D  , ,  ix����  ix���y  j���y  j����  ix����      D  , ,  k�����  k����y  lf���y  lf����  k�����      D  , ,  n����  n���y  n����y  n�����  n����      D  , ,  pl����  pl���y  q���y  q����  pl����      D  , ,  r�����  r����y  sF���y  sF����  r�����      D  , ,  u����  u���y  u����y  u�����  u����      D  , ,  wL����  wL���y  w����y  w�����  wL����      D  , ,  y�����  y����y  z:���y  z:����  y�����      D  , ,  {�����  {����y  |~���y  |~����  {�����      D  , ,  g4  #  g4  �  g�  �  g�  #  g4  #      D  , ,  ix  #  ix  �  j  �  j  #  ix  #      D  , ,  d�  �  d�  y  er  y  er  �  d�  �      D  , ,  g4  �  g4  y  g�  y  g�  �  g4  �      D  , ,  ix  �  ix  y  j  y  j  �  ix  �      D  , ,  k�  �  k�  y  lf  y  lf  �  k�  �      D  , ,  n  �  n  y  n�  y  n�  �  n  �      D  , ,  pl  �  pl  y  q  y  q  �  pl  �      D  , ,  r�  �  r�  y  sF  y  sF  �  r�  �      D  , ,  u  �  u  y  u�  y  u�  �  u  �      D  , ,  wL  �  wL  y  w�  y  w�  �  wL  �      D  , ,  y�  �  y�  y  z:  y  z:  �  y�  �      D  , ,  {�  �  {�  y  |~  y  |~  �  {�  �      D  , ,  d�  c  d�  �  er  �  er  c  d�  c      D  , ,  g4  c  g4  �  g�  �  g�  c  g4  c      D  , ,  ix  c  ix  �  j  �  j  c  ix  c      D  , ,  d�����  d����9  er���9  er����  d�����      D  , ,  g4����  g4���9  g����9  g�����  g4����      D  , ,  ix����  ix���9  j���9  j����  ix����      D  , ,  k�����  k����9  lf���9  lf����  k�����      D  , ,  n����  n���9  n����9  n�����  n����      D  , ,  pl����  pl���9  q���9  q����  pl����      D  , ,  r�����  r����9  sF���9  sF����  r�����      D  , ,  u����  u���9  u����9  u�����  u����      D  , ,  wL����  wL���9  w����9  w�����  wL����      D  , ,  y�����  y����9  z:���9  z:����  y�����      D  , ,  {�����  {����9  |~���9  |~����  {�����      D  , ,  k�  c  k�  �  lf  �  lf  c  k�  c      D  , ,  n  c  n  �  n�  �  n�  c  n  c      D  , ,  pl  c  pl  �  q  �  q  c  pl  c      D  , ,  r�  c  r�  �  sF  �  sF  c  r�  c      D  , ,  u  c  u  �  u�  �  u�  c  u  c      D  , ,  wL  c  wL  �  w�  �  w�  c  wL  c      D  , ,  y�  c  y�  �  z:  �  z:  c  y�  c      D  , ,  {�  c  {�  �  |~  �  |~  c  {�  c      D  , ,  k�  #  k�  �  lf  �  lf  #  k�  #      D  , ,  n  #  n  �  n�  �  n�  #  n  #      D  , ,  pl  #  pl  �  q  �  q  #  pl  #      D  , ,  d�  �  d�  9  er  9  er  �  d�  �      D  , ,  g4  �  g4  9  g�  9  g�  �  g4  �      D  , ,  ix  �  ix  9  j  9  j  �  ix  �      D  , ,  k�  �  k�  9  lf  9  lf  �  k�  �      D  , ,  n  �  n  9  n�  9  n�  �  n  �      D  , ,  pl  �  pl  9  q  9  q  �  pl  �      D  , ,  r�  �  r�  9  sF  9  sF  �  r�  �      D  , ,  u  �  u  9  u�  9  u�  �  u  �      D  , ,  d����c  d�����  er����  er���c  d����c      D  , ,  g4���c  g4����  g�����  g����c  g4���c      D  , ,  ix���c  ix����  j����  j���c  ix���c      D  , ,  k����c  k�����  lf����  lf���c  k����c      D  , ,  n���c  n����  n�����  n����c  n���c      D  , ,  pl���c  pl����  q����  q���c  pl���c      D  , ,  r����c  r�����  sF����  sF���c  r����c      D  , ,  u���c  u����  u�����  u����c  u���c      D  , ,  wL���c  wL����  w�����  w����c  wL���c      D  , ,  y����c  y�����  z:����  z:���c  y����c      D  , ,  {����c  {�����  |~����  |~���c  {����c      D  , ,  wL  �  wL  9  w�  9  w�  �  wL  �      D  , ,  y�  �  y�  9  z:  9  z:  �  y�  �      D  , ,  {�  �  {�  9  |~  9  |~  �  {�  �      D  , ,  r�  #  r�  �  sF  �  sF  #  r�  #      D  , ,  u  #  u  �  u�  �  u�  #  u  #      D  , ,  wL  #  wL  �  w�  �  w�  #  wL  #      D  , ,  d�   #  d�   �  er   �  er   #  d�   #      D  , ,  g4   #  g4   �  g�   �  g�   #  g4   #      D  , ,  ix   #  ix   �  j   �  j   #  ix   #      D  , ,  k�   #  k�   �  lf   �  lf   #  k�   #      D  , ,  n   #  n   �  n�   �  n�   #  n   #      D  , ,  pl   #  pl   �  q   �  q   #  pl   #      D  , ,  r�   #  r�   �  sF   �  sF   #  r�   #      D  , ,  u   #  u   �  u�   �  u�   #  u   #      D  , ,  wL   #  wL   �  w�   �  w�   #  wL   #      D  , ,  y�   #  y�   �  z:   �  z:   #  y�   #      D  , ,  {�   #  {�   �  |~   �  |~   #  {�   #      D  , ,  y�  #  y�  �  z:  �  z:  #  y�  #      D  , ,  ��  7  ��  �  �&  �  �&  7  ��  7      D  , ,  ��  7  ��  �  �~  �  �~  7  ��  7      D  , ,  �,  7  �,  �  ��  �  ��  7  �,  7      D  , ,  ��  7  ��  �  �  �  �  7  ��  7      D  , ,  ��  7  ��  �  �^  �  �^  7  ��  7      D  , ,  �   7  �   �  ��  �  ��  7  �   7      D  , ,  �d  7  �d  �  ��  �  ��  7  �d  7      D  , ,  ��  7  ��  �  �R  �  �R  7  ��  7      D  , ,  �   7  �   �  ��  �  ��  7  �   7      D  , ,  �X  7  �X  �  ��  �  ��  7  �X  7      D  , ,  �   �  �   �  ��  �  ��  �  �   �      D  , ,  �d  �  �d  �  ��  �  ��  �  �d  �      D  , ,  �   7  �   �  ��  �  ��  7  �   7      D  , ,  ��  �  ��  �  �R  �  �R  �  ��  �      D  , ,  �   �  �   �  ��  �  ��  �  �   �      D  , ,  �X  �  �X  �  ��  �  ��  �  �X  �      D  , ,  �d  7  �d  �  ��  �  ��  7  �d  7      D  , ,  ��  7  ��  �  �R  �  �R  7  ��  7      D  , ,  �   7  �   �  ��  �  ��  7  �   7      D  , ,  �X  7  �X  �  ��  �  ��  7  �X  7      D  , ,  �   w  �     ��    ��  w  �   w      D  , ,  �d  w  �d    ��    ��  w  �d  w      D  , ,  ��  w  ��    �R    �R  w  ��  w      D  , ,  �   w  �     ��    ��  w  �   w      D  , ,  �X  w  �X    ��    ��  w  �X  w      D  , ,  �   w  �     ��    ��  w  �   w      D  , ,  �d  w  �d    ��    ��  w  �d  w      D  , ,  ��  w  ��    �R    �R  w  ��  w      D  , ,  �   w  �     ��    ��  w  �   w      D  , ,  �X  w  �X    ��    ��  w  �X  w      D  , ,  �   �  �   M  ��  M  ��  �  �   �      D  , ,  �d  �  �d  M  ��  M  ��  �  �d  �      D  , ,  ��  �  ��  M  �R  M  �R  �  ��  �      D  , ,  �   �  �   M  ��  M  ��  �  �   �      D  , ,  �X  �  �X  M  ��  M  ��  �  �X  �      D  , ,  ��  �  ��  �  �&  �  �&  �  ��  �      D  , ,  ��  �  ��  �  �~  �  �~  �  ��  �      D  , ,  �,  �  �,  �  ��  �  ��  �  �,  �      D  , ,  ��  �  ��  �  �  �  �  �  ��  �      D  , ,  ��  �  ��  �  �^  �  �^  �  ��  �      D  , ,  ��  w  ��    �&    �&  w  ��  w      D  , ,  ��  w  ��    �~    �~  w  ��  w      D  , ,  �,  w  �,    ��    ��  w  �,  w      D  , ,  ��  w  ��    �    �  w  ��  w      D  , ,  ��  w  ��    �^    �^  w  ��  w      D  , ,  ��  w  ��    �&    �&  w  ��  w      D  , ,  ��  w  ��    �~    �~  w  ��  w      D  , ,  �,  w  �,    ��    ��  w  �,  w      D  , ,  ��  w  ��    �    �  w  ��  w      D  , ,  ��  w  ��    �^    �^  w  ��  w      D  , ,  ��  �  ��  M  �&  M  �&  �  ��  �      D  , ,  ��  �  ��  M  �~  M  �~  �  ��  �      D  , ,  �,  �  �,  M  ��  M  ��  �  �,  �      D  , ,  ��  �  ��  M  �  M  �  �  ��  �      D  , ,  ��  �  ��  M  �^  M  �^  �  ��  �      D  , ,  ��  7  ��  �  �&  �  �&  7  ��  7      D  , ,  ��  7  ��  �  �~  �  �~  7  ��  7      D  , ,  �,  7  �,  �  ��  �  ��  7  �,  7      D  , ,  ��  7  ��  �  �  �  �  7  ��  7      D  , ,  ��  7  ��  �  �^  �  �^  7  ��  7      D  , ,  ��  	�  ��  
#  �A  
#  �A  	�  ��  	�      D  , ,  ��  	�  ��  
#  ��  
#  ��  	�  ��  	�      D  , ,  �s  M  �s  �  �	  �  �	  M  �s  M      D  , ,  ��  M  ��  �  �W  �  �W  M  ��  M      D  , ,  ��  �  ��  M  �  M  �  �  ��  �      D  , ,  ��  �  ��  �  �&  �  �&  �  ��  �      D  , ,  ��  �  ��  �  �~  �  �~  �  ��  �      D  , ,  �  M  �  �  ��  �  ��  M  �  M      D  , ,  �]  M  �]  �  ��  �  ��  M  �]  M      D  , ,  ��  M  ��  �  �A  �  �A  M  ��  M      D  , ,  ��  M  ��  �  ��  �  ��  M  ��  M      D  , ,  �,  �  �,  �  ��  �  ��  �  �,  �      D  , ,  ��  �  ��  �  �  �  �  �  ��  �      D  , ,  ��  �  ��  �  �^  �  �^  �  ��  �      D  , ,  ��  �  ��  M  �^  M  �^  �  ��  �      D  , ,  �,  �  �,  M  ��  M  ��  �  �,  �      D  , ,  �s  	�  �s  
#  �	  
#  �	  	�  �s  	�      D  , ,  ��  	�  ��  
#  �W  
#  �W  	�  ��  	�      D  , ,  �  	�  �  
#  ��  
#  ��  	�  �  	�      D  , ,  �]  	�  �]  
#  ��  
#  ��  	�  �]  	�      D  , ,  ��  �  ��  M  �&  M  �&  �  ��  �      D  , ,  ��  �  ��  M  �~  M  �~  �  ��  �      D  , ,  �   �  �   �  ��  �  ��  �  �   �      D  , ,  �X  �  �X  �  ��  �  ��  �  �X  �      D  , ,  �G  	�  �G  
#  ��  
#  ��  	�  �G  	�      D  , ,  ��  	�  ��  
#  �+  
#  �+  	�  ��  	�      D  , ,  �G  M  �G  �  ��  �  ��  M  �G  M      D  , ,  ��  M  ��  �  �+  �  �+  M  ��  M      D  , ,  ��  M  ��  �  �y  �  �y  M  ��  M      D  , ,  �1  M  �1  �  ��  �  ��  M  �1  M      D  , ,  �  M  �  �  �  �  �  M  �  M      D  , ,  ��  	�  ��  
#  �y  
#  �y  	�  ��  	�      D  , ,  �1  	�  �1  
#  ��  
#  ��  	�  �1  	�      D  , ,  �  	�  �  
#  �  
#  �  	�  �  	�      D  , ,  �d  �  �d  M  ��  M  ��  �  �d  �      D  , ,  ��  �  ��  M  �R  M  �R  �  ��  �      D  , ,  �   �  �   M  ��  M  ��  �  �   �      D  , ,  �X  �  �X  M  ��  M  ��  �  �X  �      D  , ,  �   �  �   M  ��  M  ��  �  �   �      D  , ,  �   �  �   �  ��  �  ��  �  �   �      D  , ,  �d  �  �d  �  ��  �  ��  �  �d  �      D  , ,  ��  �  ��  �  �R  �  �R  �  ��  �      D  , ,  ��  7  ��  �  ��  �  ��  7  ��  7      D  , ,  �L  7  �L  �  ��  �  ��  7  �L  7      D  , ,  ~@  7  ~@  �  ~�  �  ~�  7  ~@  7      D  , ,  ��  7  ��  �  �  �  �  7  ��  7      D  , ,  ��  7  ��  �  �r  �  �r  7  ��  7      D  , ,  �   7  �   �  ��  �  ��  7  �   7      D  , ,  �x  7  �x  �  �  �  �  7  �x  7      D  , ,  ��  7  ��  �  �R  �  �R  7  ��  7      D  , ,  �  7  �  �  ��  �  ��  7  �  7      D  , ,  �X  7  �X  �  ��  �  ��  7  �X  7      D  , ,  ��  7  ��  �  �F  �  �F  7  ��  7      D  , ,  �X  w  �X    ��    ��  w  �X  w      D  , ,  ��  w  ��    �F    �F  w  ��  w      D  , ,  ��  �  ��  �  �R  �  �R  �  ��  �      D  , ,  �  �  �  �  ��  �  ��  �  �  �      D  , ,  �X  �  �X  �  ��  �  ��  �  �X  �      D  , ,  ��  7  ��  �  �R  �  �R  7  ��  7      D  , ,  �  7  �  �  ��  �  ��  7  �  7      D  , ,  �X  7  �X  �  ��  �  ��  7  �X  7      D  , ,  �L  w  �L    ��    ��  w  �L  w      D  , ,  ��  7  ��  �  �F  �  �F  7  ��  7      D  , ,  ��  w  ��    ��    ��  w  ��  w      D  , ,  �L  w  �L    ��    ��  w  �L  w      D  , ,  ��  w  ��    �R    �R  w  ��  w      D  , ,  �  w  �    ��    ��  w  �  w      D  , ,  �X  w  �X    ��    ��  w  �X  w      D  , ,  ��  w  ��    �F    �F  w  ��  w      D  , ,  ��  w  ��    �R    �R  w  ��  w      D  , ,  ��  �  ��  M  �R  M  �R  �  ��  �      D  , ,  �  �  �  M  ��  M  ��  �  �  �      D  , ,  �X  �  �X  M  ��  M  ��  �  �X  �      D  , ,  ��  �  ��  M  �F  M  �F  �  ��  �      D  , ,  ��  �  ��  M  ��  M  ��  �  ��  �      D  , ,  �L  �  �L  M  ��  M  ��  �  �L  �      D  , ,  ��  w  ��    ��    ��  w  ��  w      D  , ,  ��  �  ��  �  �F  �  �F  �  ��  �      D  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      D  , ,  �L  �  �L  �  ��  �  ��  �  �L  �      D  , ,  ��  7  ��  �  ��  �  ��  7  ��  7      D  , ,  �L  7  �L  �  ��  �  ��  7  �L  7      D  , ,  �  w  �    ��    ��  w  �  w      D  , ,  �x  w  �x    �    �  w  �x  w      D  , ,  �   �  �   �  ��  �  ��  �  �   �      D  , ,  ~@  �  ~@  M  ~�  M  ~�  �  ~@  �      D  , ,  ��  �  ��  M  �  M  �  �  ��  �      D  , ,  ��  �  ��  M  �r  M  �r  �  ��  �      D  , ,  �   �  �   M  ��  M  ��  �  �   �      D  , ,  �x  �  �x  M  �  M  �  �  �x  �      D  , ,  �x  �  �x  �  �  �  �  �  �x  �      D  , ,  �   w  �     ��    ��  w  �   w      D  , ,  �x  w  �x    �    �  w  �x  w      D  , ,  ��  �  ��  �  �r  �  �r  �  ��  �      D  , ,  ~@  w  ~@    ~�    ~�  w  ~@  w      D  , ,  ��  w  ��    �    �  w  ��  w      D  , ,  ��  w  ��    �r    �r  w  ��  w      D  , ,  ~@  �  ~@  �  ~�  �  ~�  �  ~@  �      D  , ,  ��  �  ��  �  �  �  �  �  ��  �      D  , ,  ~@  w  ~@    ~�    ~�  w  ~@  w      D  , ,  ��  w  ��    �    �  w  ��  w      D  , ,  ��  w  ��    �r    �r  w  ��  w      D  , ,  �   w  �     ��    ��  w  �   w      D  , ,  ~@  7  ~@  �  ~�  �  ~�  7  ~@  7      D  , ,  ��  7  ��  �  �  �  �  7  ��  7      D  , ,  ��  7  ��  �  �r  �  �r  7  ��  7      D  , ,  �   7  �   �  ��  �  ��  7  �   7      D  , ,  �x  7  �x  �  �  �  �  7  �x  7      D  , ,  ��  M  ��  �  �5  �  �5  M  ��  M      D  , ,  �Q  	�  �Q  
#  ��  
#  ��  	�  �Q  	�      D  , ,  ��  	�  ��  
#  �5  
#  �5  	�  ��  	�      D  , ,  �   �  �   �  ��  �  ��  �  �   �      D  , ,  �x  �  �x  �  �  �  �  �  �x  �      D  , ,  }  	�  }  
#  }�  
#  }�  	�  }  	�      D  , ,  g  	�  g  
#  �  
#  �  	�  g  	�      D  , ,  ~@  �  ~@  M  ~�  M  ~�  �  ~@  �      D  , ,  ��  �  ��  M  �  M  �  �  ��  �      D  , ,  ��  	�  ��  
#  �K  
#  �K  	�  ��  	�      D  , ,  �  	�  �  
#  ��  
#  ��  	�  �  	�      D  , ,  ~@  �  ~@  �  ~�  �  ~�  �  ~@  �      D  , ,  ��  �  ��  M  �r  M  �r  �  ��  �      D  , ,  �   �  �   M  ��  M  ��  �  �   �      D  , ,  �x  �  �x  M  �  M  �  �  �x  �      D  , ,  ��  �  ��  �  �  �  �  �  ��  �      D  , ,  ��  �  ��  �  �r  �  �r  �  ��  �      D  , ,  }  M  }  �  }�  �  }�  M  }  M      D  , ,  g  M  g  �  �  �  �  M  g  M      D  , ,  ��  M  ��  �  �K  �  �K  M  ��  M      D  , ,  �  M  �  �  ��  �  ��  M  �  M      D  , ,  �Q  M  �Q  �  ��  �  ��  M  �Q  M      D  , ,  ��  	�  ��  
#  �  
#  �  	�  ��  	�      D  , ,  ��  	�  ��  
#  �m  
#  �m  	�  ��  	�      D  , ,  �%  	�  �%  
#  ��  
#  ��  	�  �%  	�      D  , ,  �X  �  �X  �  ��  �  ��  �  �X  �      D  , ,  ��  �  ��  �  �F  �  �F  �  ��  �      D  , ,  ��  M  ��  �  ��  �  ��  M  ��  M      D  , ,  �;  M  �;  �  ��  �  ��  M  �;  M      D  , ,  ��  M  ��  �  �  �  �  M  ��  M      D  , ,  ��  M  ��  �  �m  �  �m  M  ��  M      D  , ,  ��  �  ��  M  �R  M  �R  �  ��  �      D  , ,  �  �  �  M  ��  M  ��  �  �  �      D  , ,  �X  �  �X  M  ��  M  ��  �  �X  �      D  , ,  ��  �  ��  M  �F  M  �F  �  ��  �      D  , ,  ��  �  ��  M  ��  M  ��  �  ��  �      D  , ,  �L  �  �L  M  ��  M  ��  �  �L  �      D  , ,  �%  M  �%  �  ��  �  ��  M  �%  M      D  , ,  ��  �  ��  �  �R  �  �R  �  ��  �      D  , ,  �  �  �  �  ��  �  ��  �  �  �      D  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      D  , ,  �L  �  �L  �  ��  �  ��  �  �L  �      D  , ,  ��  	�  ��  
#  ��  
#  ��  	�  ��  	�      D  , ,  �;  	�  �;  
#  ��  
#  ��  	�  �;  	�      D  , ,  �   �  �   9  ��  9  ��  �  �   �      D  , ,  �x  �  �x  9  �  9  �  �  �x  �      D  , ,  ��  �  ��  9  �R  9  �R  �  ��  �      D  , ,  �  �  �  9  ��  9  ��  �  �  �      D  , ,  �X  �  �X  9  ��  9  ��  �  �X  �      D  , ,  ��  �  ��  9  �F  9  �F  �  ��  �      D  , ,  ��  �  ��  9  ��  9  ��  �  ��  �      D  , ,  ~@����  ~@���9  ~����9  ~�����  ~@����      D  , ,  ������  �����9  ����9  �����  ������      D  , ,  ������  �����9  �r���9  �r����  ������      D  , ,  � ����  � ���9  �����9  ������  � ����      D  , ,  �x����  �x���9  ����9  �����  �x����      D  , ,  ������  �����9  �R���9  �R����  ������      D  , ,  �����  ����9  �����9  ������  �����      D  , ,  �X����  �X���9  �����9  ������  �X����      D  , ,  ������  �����9  �F���9  �F����  ������      D  , ,  ������  �����9  �����9  ������  ������      D  , ,  �L����  �L���9  �����9  ������  �L����      D  , ,  �L  �  �L  9  ��  9  ��  �  �L  �      D  , ,  ��  �  ��  y  �F  y  �F  �  ��  �      D  , ,  ��  �  ��  y  ��  y  ��  �  ��  �      D  , ,  �L  �  �L  y  ��  y  ��  �  �L  �      D  , ,  ~@  �  ~@  y  ~�  y  ~�  �  ~@  �      D  , ,  ��  �  ��  y  �  y  �  �  ��  �      D  , ,  ��  �  ��  y  �r  y  �r  �  ��  �      D  , ,  �   �  �   y  ��  y  ��  �  �   �      D  , ,  �x  �  �x  y  �  y  �  �  �x  �      D  , ,  ~@  c  ~@  �  ~�  �  ~�  c  ~@  c      D  , ,  ��  c  ��  �  �  �  �  c  ��  c      D  , ,  ~@  #  ~@  �  ~�  �  ~�  #  ~@  #      D  , ,  ��  #  ��  �  �  �  �  #  ��  #      D  , ,  ��  #  ��  �  �r  �  �r  #  ��  #      D  , ,  �   #  �   �  ��  �  ��  #  �   #      D  , ,  �x  #  �x  �  �  �  �  #  �x  #      D  , ,  ��  #  ��  �  �R  �  �R  #  ��  #      D  , ,  �  #  �  �  ��  �  ��  #  �  #      D  , ,  �X  #  �X  �  ��  �  ��  #  �X  #      D  , ,  ��  #  ��  �  �F  �  �F  #  ��  #      D  , ,  ��  #  ��  �  ��  �  ��  #  ��  #      D  , ,  �L  #  �L  �  ��  �  ��  #  �L  #      D  , ,  ~@���c  ~@����  ~�����  ~����c  ~@���c      D  , ,  �����c  ������  �����  ����c  �����c      D  , ,  �����c  ������  �r����  �r���c  �����c      D  , ,  � ���c  � ����  ������  �����c  � ���c      D  , ,  �x���c  �x����  �����  ����c  �x���c      D  , ,  �����c  ������  �R����  �R���c  �����c      D  , ,  ����c  �����  ������  �����c  ����c      D  , ,  �X���c  �X����  ������  �����c  �X���c      D  , ,  �����c  ������  �F����  �F���c  �����c      D  , ,  �����c  ������  ������  �����c  �����c      D  , ,  �L���c  �L����  ������  �����c  �L���c      D  , ,  ��  c  ��  �  �r  �  �r  c  ��  c      D  , ,  �   c  �   �  ��  �  ��  c  �   c      D  , ,  �x  c  �x  �  �  �  �  c  �x  c      D  , ,  ~@����  ~@���y  ~����y  ~�����  ~@����      D  , ,  ������  �����y  ����y  �����  ������      D  , ,  ������  �����y  �r���y  �r����  ������      D  , ,  � ����  � ���y  �����y  ������  � ����      D  , ,  �x����  �x���y  ����y  �����  �x����      D  , ,  ������  �����y  �R���y  �R����  ������      D  , ,  �����  ����y  �����y  ������  �����      D  , ,  �X����  �X���y  �����y  ������  �X����      D  , ,  ������  �����y  �F���y  �F����  ������      D  , ,  ������  �����y  �����y  ������  ������      D  , ,  �L����  �L���y  �����y  ������  �L����      D  , ,  ��  c  ��  �  �R  �  �R  c  ��  c      D  , ,  �  c  �  �  ��  �  ��  c  �  c      D  , ,  �X  c  �X  �  ��  �  ��  c  �X  c      D  , ,  ~@   #  ~@   �  ~�   �  ~�   #  ~@   #      D  , ,  ��   #  ��   �  �   �  �   #  ��   #      D  , ,  ��   #  ��   �  �r   �  �r   #  ��   #      D  , ,  �    #  �    �  ��   �  ��   #  �    #      D  , ,  �x   #  �x   �  �   �  �   #  �x   #      D  , ,  ��   #  ��   �  �R   �  �R   #  ��   #      D  , ,  �   #  �   �  ��   �  ��   #  �   #      D  , ,  �X   #  �X   �  ��   �  ��   #  �X   #      D  , ,  ��   #  ��   �  �F   �  �F   #  ��   #      D  , ,  ��   #  ��   �  ��   �  ��   #  ��   #      D  , ,  �L   #  �L   �  ��   �  ��   #  �L   #      D  , ,  ��  c  ��  �  �F  �  �F  c  ��  c      D  , ,  ��  c  ��  �  ��  �  ��  c  ��  c      D  , ,  �L  c  �L  �  ��  �  ��  c  �L  c      D  , ,  ��  �  ��  y  �R  y  �R  �  ��  �      D  , ,  �  �  �  y  ��  y  ��  �  �  �      D  , ,  �X  �  �X  y  ��  y  ��  �  �X  �      D  , ,  ~@  �  ~@  9  ~�  9  ~�  �  ~@  �      D  , ,  ��  �  ��  9  �  9  �  �  ��  �      D  , ,  ��  �  ��  9  �r  9  �r  �  ��  �      D  , ,  ��  �  ��  9  �^  9  �^  �  ��  �      D  , ,  �   �  �   9  ��  9  ��  �  �   �      D  , ,  �d  �  �d  9  ��  9  ��  �  �d  �      D  , ,  ��  �  ��  9  �R  9  �R  �  ��  �      D  , ,  �   �  �   9  ��  9  ��  �  �   �      D  , ,  �X  �  �X  9  ��  9  ��  �  �X  �      D  , ,  ��  �  ��  y  �~  y  �~  �  ��  �      D  , ,  ��  c  ��  �  �&  �  �&  c  ��  c      D  , ,  ��  c  ��  �  �~  �  �~  c  ��  c      D  , ,  �,  c  �,  �  ��  �  ��  c  �,  c      D  , ,  ��  c  ��  �  �  �  �  c  ��  c      D  , ,  ��  c  ��  �  �^  �  �^  c  ��  c      D  , ,  ��  #  ��  �  �&  �  �&  #  ��  #      D  , ,  ��  #  ��  �  �~  �  �~  #  ��  #      D  , ,  �,  #  �,  �  ��  �  ��  #  �,  #      D  , ,  ��  #  ��  �  �  �  �  #  ��  #      D  , ,  ��  #  ��  �  �^  �  �^  #  ��  #      D  , ,  �   #  �   �  ��  �  ��  #  �   #      D  , ,  �d  #  �d  �  ��  �  ��  #  �d  #      D  , ,  ��  #  ��  �  �R  �  �R  #  ��  #      D  , ,  �   c  �   �  ��  �  ��  c  �   c      D  , ,  �d  c  �d  �  ��  �  ��  c  �d  c      D  , ,  ��  c  ��  �  �R  �  �R  c  ��  c      D  , ,  �   c  �   �  ��  �  ��  c  �   c      D  , ,  �X  c  �X  �  ��  �  ��  c  �X  c      D  , ,  �,  �  �,  y  ��  y  ��  �  �,  �      D  , ,  ��  �  ��  y  �  y  �  �  ��  �      D  , ,  ��  �  ��  y  �^  y  �^  �  ��  �      D  , ,  �   �  �   y  ��  y  ��  �  �   �      D  , ,  �d  �  �d  y  ��  y  ��  �  �d  �      D  , ,  ��  �  ��  y  �R  y  �R  �  ��  �      D  , ,  �����c  ������  �&����  �&���c  �����c      D  , ,  �����c  ������  �~����  �~���c  �����c      D  , ,  �,���c  �,����  ������  �����c  �,���c      D  , ,  �����c  ������  �����  ����c  �����c      D  , ,  �����c  ������  �^����  �^���c  �����c      D  , ,  � ���c  � ����  ������  �����c  � ���c      D  , ,  �d���c  �d����  ������  �����c  �d���c      D  , ,  �����c  ������  �R����  �R���c  �����c      D  , ,  � ���c  � ����  ������  �����c  � ���c      D  , ,  �X���c  �X����  ������  �����c  �X���c      D  , ,  �   #  �   �  ��  �  ��  #  �   #      D  , ,  �   �  �   y  ��  y  ��  �  �   �      D  , ,  �X  �  �X  y  ��  y  ��  �  �X  �      D  , ,  ��  �  ��  y  �&  y  �&  �  ��  �      D  , ,  ��  �  ��  9  �&  9  �&  �  ��  �      D  , ,  ��  �  ��  9  �~  9  �~  �  ��  �      D  , ,  ��   #  ��   �  �&   �  �&   #  ��   #      D  , ,  ��   #  ��   �  �~   �  �~   #  ��   #      D  , ,  �,   #  �,   �  ��   �  ��   #  �,   #      D  , ,  ��   #  ��   �  �   �  �   #  ��   #      D  , ,  ��   #  ��   �  �^   �  �^   #  ��   #      D  , ,  �    #  �    �  ��   �  ��   #  �    #      D  , ,  �d   #  �d   �  ��   �  ��   #  �d   #      D  , ,  ��   #  ��   �  �R   �  �R   #  ��   #      D  , ,  �    #  �    �  ��   �  ��   #  �    #      D  , ,  �X   #  �X   �  ��   �  ��   #  �X   #      D  , ,  �,  �  �,  9  ��  9  ��  �  �,  �      D  , ,  ������  �����y  �&���y  �&����  ������      D  , ,  ������  �����9  �&���9  �&����  ������      D  , ,  ������  �����9  �~���9  �~����  ������      D  , ,  �,����  �,���9  �����9  ������  �,����      D  , ,  ������  �����9  ����9  �����  ������      D  , ,  �X  #  �X  �  ��  �  ��  #  �X  #      D  , ,  ������  �����9  �^���9  �^����  ������      D  , ,  � ����  � ���9  �����9  ������  � ����      D  , ,  �d����  �d���9  �����9  ������  �d����      D  , ,  ������  �����9  �R���9  �R����  ������      D  , ,  � ����  � ���9  �����9  ������  � ����      D  , ,  �X����  �X���9  �����9  ������  �X����      D  , ,  ������  �����y  �~���y  �~����  ������      D  , ,  �,����  �,���y  �����y  ������  �,����      D  , ,  ������  �����y  ����y  �����  ������      D  , ,  ������  �����y  �^���y  �^����  ������      D  , ,  � ����  � ���y  �����y  ������  � ����      D  , ,  �d����  �d���y  �����y  ������  �d����      D  , ,  ������  �����y  �R���y  �R����  ������      D  , ,  � ����  � ���y  �����y  ������  � ����      D  , ,  �X����  �X���y  �����y  ������  �X����      D  , ,  ��  �  ��  9  �  9  �  �  ��  �      D  , ,  ~@����  ~@���  ~����  ~�����  ~@����      D  , ,  ������  �����  ����  �����  ������      D  , ,  ������  �����  �r���  �r����  ������      D  , ,  � ����  � ���  �����  ������  � ����      D  , ,  �x����  �x���  ����  �����  �x����      D  , ,  ������  �����  �R���  �R����  ������      D  , ,  �����  ����  �����  ������  �����      D  , ,  �X����  �X���  �����  ������  �X����      D  , ,  ������  �����  �F���  �F����  ������      D  , ,  ������  �����  �����  ������  ������      D  , ,  �L����  �L���  �����  ������  �L����      D  , ,  ������  �����  �&���  �&����  ������      D  , ,  ������  �����  �~���  �~����  ������      D  , ,  �,����  �,���  �����  ������  �,����      D  , ,  ������  �����  ����  �����  ������      D  , ,  ������  �����  �^���  �^����  ������      D  , ,  � ����  � ���  �����  ������  � ����      D  , ,  �d����  �d���  �����  ������  �d����      D  , ,  ������  �����  �R���  �R����  ������      D  , ,  � ����  � ���  �����  ������  � ����      D  , ,  �X����  �X���  �����  ������  �X����      D  , ,  �d���m  �d���  �����  �����m  �d���m      D  , ,  �����m  �����  �R���  �R���m  �����m      D  , ,  � ���m  � ���  �����  �����m  � ���m      D  , ,  �X���m  �X���  �����  �����m  �X���m      D  , ,  �����-  ������  �&����  �&���-  �����-      D  , ,  �����-  ������  �~����  �~���-  �����-      D  , ,  �,���-  �,����  ������  �����-  �,���-      D  , ,  �����-  ������  �����  ����-  �����-      D  , ,  �����-  ������  �^����  �^���-  �����-      D  , ,  � ���-  � ����  ������  �����-  � ���-      D  , ,  �d���-  �d����  ������  �����-  �d���-      D  , ,  �����-  ������  �R����  �R���-  �����-      D  , ,  � ���-  � ����  ������  �����-  � ���-      D  , ,  �X���-  �X����  ������  �����-  �X���-      D  , ,  ������  �����'  �~���'  �~����  ������      D  , ,  ������  �����'  ����'  �����  ������      D  , ,  � ����  � ���'  �����'  ������  � ����      D  , ,  ������  �����'  �R���'  �R����  ������      D  , ,  �X����  �X���'  �����'  ������  �X����      D  , ,  �����Q  ������  �~����  �~���Q  �����Q      D  , ,  �����Q  ������  �����  ����Q  �����Q      D  , ,  � ���Q  � ����  ������  �����Q  � ���Q      D  , ,  �����Q  ������  �R����  �R���Q  �����Q      D  , ,  �X���Q  �X����  ������  �����Q  �X���Q      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �����  ������  �����  ����  �����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �����  ������  �R����  �R���  �����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  �����m  �����  �&���  �&���m  �����m      D  , ,  �����m  �����  �~���  �~���m  �����m      D  , ,  �,���m  �,���  �����  �����m  �,���m      D  , ,  �����m  �����  ����  ����m  �����m      D  , ,  �����m  �����  �^���  �^���m  �����m      D  , ,  � ���m  � ���  �����  �����m  � ���m      D  , ,  ������  �����g  �~���g  �~����  ������      D  , ,  ������  �����g  ����g  �����  ������      D  , ,  � ����  � ���g  �����g  ������  � ����      D  , ,  ������  �����g  �R���g  �R����  ������      D  , ,  �X����  �X���g  �����g  ������  �X����      D  , ,  �X���-  �X����  ������  �����-  �X���-      D  , ,  �����-  ������  �F����  �F���-  �����-      D  , ,  �����-  ������  ������  �����-  �����-      D  , ,  �L���-  �L����  ������  �����-  �L���-      D  , ,  ����  �����  ������  �����  ����      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  ������  �����'  �F���'  �F����  ������      D  , ,  ~@���Q  ~@����  ~�����  ~����Q  ~@���Q      D  , ,  �����Q  ������  �r����  �r���Q  �����Q      D  , ,  �x���Q  �x����  �����  ����Q  �x���Q      D  , ,  ����Q  �����  ������  �����Q  ����Q      D  , ,  ~@���m  ~@���  ~����  ~����m  ~@���m      D  , ,  �����m  �����  ����  ����m  �����m      D  , ,  �����m  �����  �r���  �r���m  �����m      D  , ,  � ���m  � ���  �����  �����m  � ���m      D  , ,  �x���m  �x���  ����  ����m  �x���m      D  , ,  �����m  �����  �R���  �R���m  �����m      D  , ,  ����m  ����  �����  �����m  ����m      D  , ,  �X���m  �X���  �����  �����m  �X���m      D  , ,  �����m  �����  �F���  �F���m  �����m      D  , ,  �����m  �����  �����  �����m  �����m      D  , ,  �L���m  �L���  �����  �����m  �L���m      D  , ,  �����Q  ������  �F����  �F���Q  �����Q      D  , ,  �L���Q  �L����  ������  �����Q  �L���Q      D  , ,  �L����  �L���'  �����'  ������  �L����      D  , ,  ~@����  ~@���'  ~����'  ~�����  ~@����      D  , ,  ������  �����'  �r���'  �r����  ������      D  , ,  �x����  �x���'  ����'  �����  �x����      D  , ,  �����  ����'  �����'  ������  �����      D  , ,  ~@���  ~@����  ~�����  ~����  ~@���      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  ~@���-  ~@����  ~�����  ~����-  ~@���-      D  , ,  �����-  ������  �����  ����-  �����-      D  , ,  ~@����  ~@���g  ~����g  ~�����  ~@����      D  , ,  ������  �����g  �r���g  �r����  ������      D  , ,  �x����  �x���g  ����g  �����  �x����      D  , ,  �����  ����g  �����g  ������  �����      D  , ,  ������  �����g  �F���g  �F����  ������      D  , ,  �L����  �L���g  �����g  ������  �L����      D  , ,  �����-  ������  �r����  �r���-  �����-      D  , ,  � ���-  � ����  ������  �����-  � ���-      D  , ,  �x���-  �x����  �����  ����-  �x���-      D  , ,  �����-  ������  �R����  �R���-  �����-      D  , ,  ����-  �����  ������  �����-  ����-      D  , ,  ~@���m  ~@���  ~����  ~����m  ~@���m      D  , ,  �����m  �����  ����  ����m  �����m      D  , ,  �����m  �����  �r���  �r���m  �����m      D  , ,  � ���m  � ���  �����  �����m  � ���m      D  , ,  �x���m  �x���  ����  ����m  �x���m      D  , ,  �����m  �����  �R���  �R���m  �����m      D  , ,  ����m  ����  �����  �����m  ����m      D  , ,  �X���m  �X���  �����  �����m  �X���m      D  , ,  �����m  �����  �F���  �F���m  �����m      D  , ,  �����m  �����  �����  �����m  �����m      D  , ,  �L���m  �L���  �����  �����m  �L���m      D  , ,  ~@���-  ~@����  ~�����  ~����-  ~@���-      D  , ,  �����-  ������  �����  ����-  �����-      D  , ,  �����-  ������  �r����  �r���-  �����-      D  , ,  � ���-  � ����  ������  �����-  � ���-      D  , ,  �x���-  �x����  �����  ����-  �x���-      D  , ,  �����-  ������  �R����  �R���-  �����-      D  , ,  ����-  �����  ������  �����-  ����-      D  , ,  �X���-  �X����  ������  �����-  �X���-      D  , ,  �����-  ������  �F����  �F���-  �����-      D  , ,  �����-  ������  ������  �����-  �����-      D  , ,  �L���-  �L����  ������  �����-  �L���-      D  , ,  ~@����  ~@���  ~����  ~�����  ~@����      D  , ,  ������  �����  ����  �����  ������      D  , ,  ������  �����  �r���  �r����  ������      D  , ,  � ����  � ���  �����  ������  � ����      D  , ,  �x����  �x���  ����  �����  �x����      D  , ,  ������  �����  �R���  �R����  ������      D  , ,  �����  ����  �����  ������  �����      D  , ,  �X����  �X���  �����  ������  �X����      D  , ,  ������  �����  �F���  �F����  ������      D  , ,  ������  �����  �����  ������  ������      D  , ,  �L����  �L���  �����  ������  �L����      D  , ,  ~@���  ~@���C  ~����C  ~����  ~@���      D  , ,  �����  �����C  ����C  ����  �����      D  , ,  �����  �����C  �r���C  �r���  �����      D  , ,  � ���  � ���C  �����C  �����  � ���      D  , ,  �x���  �x���C  ����C  ����  �x���      D  , ,  �����  �����C  �R���C  �R���  �����      D  , ,  ����  ����C  �����C  �����  ����      D  , ,  �X���  �X���C  �����C  �����  �X���      D  , ,  �����  �����C  �F���C  �F���  �����      D  , ,  �����  �����C  �����C  �����  �����      D  , ,  �L���  �L���C  �����C  �����  �L���      D  , ,  ~@���  ~@���C  ~����C  ~����  ~@���      D  , ,  }���  }���  }����  }����  }���      D  , ,  g���  g���  ����  ����  g���      D  , ,  �����  �����  �K���  �K���  �����      D  , ,  ����  ����  �����  �����  ����      D  , ,  �Q���  �Q���  �����  �����  �Q���      D  , ,  �����  �����  �5���  �5���  �����      D  , ,  �����  �����  �����  �����  �����      D  , ,  �;���  �;���  �����  �����  �;���      D  , ,  �����  �����  ����  ����  �����      D  , ,  �����  �����  �m���  �m���  �����      D  , ,  �%���  �%���  �����  �����  �%���      D  , ,  }���C  }����  }�����  }����C  }���C      D  , ,  g���C  g����  �����  ����C  g���C      D  , ,  �����C  ������  �K����  �K���C  �����C      D  , ,  ����C  �����  ������  �����C  ����C      D  , ,  �Q���C  �Q����  ������  �����C  �Q���C      D  , ,  �����C  ������  �5����  �5���C  �����C      D  , ,  �����C  ������  ������  �����C  �����C      D  , ,  �;���C  �;����  ������  �����C  �;���C      D  , ,  �����C  ������  �����  ����C  �����C      D  , ,  �����C  ������  �m����  �m���C  �����C      D  , ,  �%���C  �%����  ������  �����C  �%���C      D  , ,  ~@���  ~@��ݯ  ~���ݯ  ~����  ~@���      D  , ,  �����  ����ݯ  ���ݯ  ����  �����      D  , ,  �����  ����ݯ  �r��ݯ  �r���  �����      D  , ,  � ���  � ��ݯ  ����ݯ  �����  � ���      D  , ,  �x���  �x��ݯ  ���ݯ  ����  �x���      D  , ,  �����  ����ݯ  �R��ݯ  �R���  �����      D  , ,  ����  ���ݯ  ����ݯ  �����  ����      D  , ,  �X���  �X��ݯ  ����ݯ  �����  �X���      D  , ,  �����  ����ݯ  �F��ݯ  �F���  �����      D  , ,  �����  ����ݯ  ����ݯ  �����  �����      D  , ,  �L���  �L��ݯ  ����ݯ  �����  �L���      D  , ,  �����  �����C  ����C  ����  �����      D  , ,  �����  �����C  �r���C  �r���  �����      D  , ,  � ���  � ���C  �����C  �����  � ���      D  , ,  �x���  �x���C  ����C  ����  �x���      D  , ,  �����  �����C  �R���C  �R���  �����      D  , ,  ����  ����C  �����C  �����  ����      D  , ,  �X���  �X���C  �����C  �����  �X���      D  , ,  �����  �����C  �F���C  �F���  �����      D  , ,  �����  �����C  �����C  �����  �����      D  , ,  �L���  �L���C  �����C  �����  �L���      D  , ,  �����  �����C  �^���C  �^���  �����      D  , ,  � ���  � ���C  �����C  �����  � ���      D  , ,  �d���  �d���C  �����C  �����  �d���      D  , ,  �����  �����C  �R���C  �R���  �����      D  , ,  � ���  � ���C  �����C  �����  � ���      D  , ,  �X���  �X���C  �����C  �����  �X���      D  , ,  �,���-  �,����  ������  �����-  �,���-      D  , ,  �����-  ������  �����  ����-  �����-      D  , ,  �����-  ������  �^����  �^���-  �����-      D  , ,  � ���-  � ����  ������  �����-  � ���-      D  , ,  �d���-  �d����  ������  �����-  �d���-      D  , ,  �����-  ������  �R����  �R���-  �����-      D  , ,  � ���-  � ����  ������  �����-  � ���-      D  , ,  �X���-  �X����  ������  �����-  �X���-      D  , ,  �����m  �����  �~���  �~���m  �����m      D  , ,  �,���m  �,���  �����  �����m  �,���m      D  , ,  �����m  �����  ����  ����m  �����m      D  , ,  �����m  �����  �^���  �^���m  �����m      D  , ,  �s���  �s���  �	���  �	���  �s���      D  , ,  �����  �����  �W���  �W���  �����      D  , ,  ����  ����  �����  �����  ����      D  , ,  �]���  �]���  �����  �����  �]���      D  , ,  �����  �����  �A���  �A���  �����      D  , ,  �����  �����  �����  �����  �����      D  , ,  �G���  �G���  �����  �����  �G���      D  , ,  �����  �����  �+���  �+���  �����      D  , ,  �����  �����  �y���  �y���  �����      D  , ,  �1���  �1���  �����  �����  �1���      D  , ,  ����  ����  ����  ����  ����      D  , ,  � ���m  � ���  �����  �����m  � ���m      D  , ,  �d���m  �d���  �����  �����m  �d���m      D  , ,  �����m  �����  �R���  �R���m  �����m      D  , ,  � ���m  � ���  �����  �����m  � ���m      D  , ,  �X���m  �X���  �����  �����m  �X���m      D  , ,  �����  �����C  �~���C  �~���  �����      D  , ,  �,���  �,���C  �����C  �����  �,���      D  , ,  ������  �����  �&���  �&����  ������      D  , ,  ������  �����  �~���  �~����  ������      D  , ,  �,����  �,���  �����  ������  �,����      D  , ,  ������  �����  ����  �����  ������      D  , ,  �s���C  �s����  �	����  �	���C  �s���C      D  , ,  �����C  ������  �W����  �W���C  �����C      D  , ,  ����C  �����  ������  �����C  ����C      D  , ,  �]���C  �]����  ������  �����C  �]���C      D  , ,  �����C  ������  �A����  �A���C  �����C      D  , ,  �����C  ������  ������  �����C  �����C      D  , ,  �G���C  �G����  ������  �����C  �G���C      D  , ,  �����C  ������  �+����  �+���C  �����C      D  , ,  �����C  ������  �y����  �y���C  �����C      D  , ,  �1���C  �1����  ������  �����C  �1���C      D  , ,  ����C  �����  �����  ����C  ����C      D  , ,  ������  �����  �^���  �^����  ������      D  , ,  � ����  � ���  �����  ������  � ����      D  , ,  �d����  �d���  �����  ������  �d����      D  , ,  ������  �����  �R���  �R����  ������      D  , ,  � ����  � ���  �����  ������  � ����      D  , ,  �X����  �X���  �����  ������  �X����      D  , ,  �����  �����C  ����C  ����  �����      D  , ,  �����  �����C  �^���C  �^���  �����      D  , ,  � ���  � ���C  �����C  �����  � ���      D  , ,  �d���  �d���C  �����C  �����  �d���      D  , ,  �����  �����C  �R���C  �R���  �����      D  , ,  �����  ����ݯ  �&��ݯ  �&���  �����      D  , ,  �����  ����ݯ  �~��ݯ  �~���  �����      D  , ,  �,���  �,��ݯ  ����ݯ  �����  �,���      D  , ,  �����  ����ݯ  ���ݯ  ����  �����      D  , ,  �����  ����ݯ  �^��ݯ  �^���  �����      D  , ,  � ���  � ��ݯ  ����ݯ  �����  � ���      D  , ,  �d���  �d��ݯ  ����ݯ  �����  �d���      D  , ,  �����  ����ݯ  �R��ݯ  �R���  �����      D  , ,  � ���  � ��ݯ  ����ݯ  �����  � ���      D  , ,  �X���  �X��ݯ  ����ݯ  �����  �X���      D  , ,  � ���  � ���C  �����C  �����  � ���      D  , ,  �X���  �X���C  �����C  �����  �X���      D  , ,  �����  �����C  �&���C  �&���  �����      D  , ,  �����m  �����  �&���  �&���m  �����m      D  , ,  �����-  ������  �&����  �&���-  �����-      D  , ,  �����-  ������  �~����  �~���-  �����-      D  , ,  �����  �����C  �&���C  �&���  �����      D  , ,  �����  �����C  �~���C  �~���  �����      D  , ,  �,���  �,���C  �����C  �����  �,���      D  , ,  �����  �����C  ����C  ����  �����      D  , ,  c����  c����  dU���  dU���  c����      D  , ,  ]�����  ]����  ^����  ^�����  ]�����      D  , ,  `@����  `@���  `����  `�����  `@����      D  , ,  b�����  b����  c.���  c.����  b�����      D  , ,  d�����  d����  er���  er����  d�����      D  , ,  g4����  g4���  g����  g�����  g4����      D  , ,  ix����  ix���  j���  j����  ix����      D  , ,  k�����  k����  lf���  lf����  k�����      D  , ,  n����  n���  n����  n�����  n����      D  , ,  pl����  pl���  q���  q����  pl����      D  , ,  r�����  r����  sF���  sF����  r�����      D  , ,  u����  u���  u����  u�����  u����      D  , ,  wL����  wL���  w����  w�����  wL����      D  , ,  y�����  y����  z:���  z:����  y�����      D  , ,  c����C  c�����  dU����  dU���C  c����C      D  , ,  {�����  {����  |~���  |~����  {�����      D  , ,  u���  u����  u�����  u����  u���      D  , ,  y����  y�����  z:����  z:���  y����      D  , ,  g4���Q  g4����  g�����  g����Q  g4���Q      D  , ,  k����Q  k�����  lf����  lf���Q  k����Q      D  , ,  k�����  k����g  lf���g  lf����  k�����      D  , ,  wL���-  wL����  w�����  w����-  wL���-      D  , ,  pl���Q  pl����  q����  q���Q  pl���Q      D  , ,  u���Q  u����  u�����  u����Q  u���Q      D  , ,  y����Q  y�����  z:����  z:���Q  y����Q      D  , ,  y����-  y�����  z:����  z:���-  y����-      D  , ,  {����-  {�����  |~����  |~���-  {����-      D  , ,  ix���m  ix���  j���  j���m  ix���m      D  , ,  k����m  k����  lf���  lf���m  k����m      D  , ,  n���m  n���  n����  n����m  n���m      D  , ,  pl���m  pl���  q���  q���m  pl���m      D  , ,  r����m  r����  sF���  sF���m  r����m      D  , ,  u���m  u���  u����  u����m  u���m      D  , ,  y�����  y����g  z:���g  z:����  y�����      D  , ,  wL���m  wL���  w����  w����m  wL���m      D  , ,  y����m  y����  z:���  z:���m  y����m      D  , ,  {����m  {����  |~���  |~���m  {����m      D  , ,  g4���  g4����  g�����  g����  g4���      D  , ,  k����  k�����  lf����  lf���  k����      D  , ,  pl���  pl����  q����  q���  pl���      D  , ,  y�����  y����'  z:���'  z:����  y�����      D  , ,  u����  u���'  u����'  u�����  u����      D  , ,  pl����  pl���g  q���g  q����  pl����      D  , ,  d����m  d����  er���  er���m  d����m      D  , ,  g4���m  g4���  g����  g����m  g4���m      D  , ,  d����-  d�����  er����  er���-  d����-      D  , ,  g4���-  g4����  g�����  g����-  g4���-      D  , ,  ix���-  ix����  j����  j���-  ix���-      D  , ,  k����-  k�����  lf����  lf���-  k����-      D  , ,  n���-  n����  n�����  n����-  n���-      D  , ,  pl���-  pl����  q����  q���-  pl���-      D  , ,  r����-  r�����  sF����  sF���-  r����-      D  , ,  u���-  u����  u�����  u����-  u���-      D  , ,  g4����  g4���g  g����g  g�����  g4����      D  , ,  u����  u���g  u����g  u�����  u����      D  , ,  g4����  g4���'  g����'  g�����  g4����      D  , ,  k�����  k����'  lf���'  lf����  k�����      D  , ,  pl����  pl���'  q���'  q����  pl����      D  , ,  b�����  b����g  c.���g  c.����  b�����      D  , ,  b����  b�����  c.����  c.���  b����      D  , ,  ]����m  ]����  ^����  ^����m  ]����m      D  , ,  `@���m  `@���  `����  `����m  `@���m      D  , ,  b����m  b����  c.���  c.���m  b����m      D  , ,  b����Q  b�����  c.����  c.���Q  b����Q      D  , ,  ]����Q  ]�����  ^�����  ^����Q  ]����Q      D  , ,  ]�����  ]����g  ^����g  ^�����  ]�����      D  , ,  ]����-  ]�����  ^�����  ^����-  ]����-      D  , ,  ]�����  ]����'  ^����'  ^�����  ]�����      D  , ,  b�����  b����'  c.���'  c.����  b�����      D  , ,  `@���-  `@����  `�����  `����-  `@���-      D  , ,  b����-  b�����  c.����  c.���-  b����-      D  , ,  ]����  ]�����  ^�����  ^����  ]����      D  , ,  b����  b����C  c.���C  c.���  b����      D  , ,  ]����m  ]����  ^����  ^����m  ]����m      D  , ,  `@���m  `@���  `����  `����m  `@���m      D  , ,  ]����-  ]�����  ^�����  ^����-  ]����-      D  , ,  `@���-  `@����  `�����  `����-  `@���-      D  , ,  b����-  b�����  c.����  c.���-  b����-      D  , ,  b����m  b����  c.���  c.���m  b����m      D  , ,  _#���  _#���  _����  _����  _#���      D  , ,  aq���  aq���  b���  b���  aq���      D  , ,  ]����  ]���ݯ  ^���ݯ  ^����  ]����      D  , ,  `@���  `@��ݯ  `���ݯ  `����  `@���      D  , ,  ]����  ]����C  ^����C  ^����  ]����      D  , ,  `@���  `@���C  `����C  `����  `@���      D  , ,  b����  b���ݯ  c.��ݯ  c.���  b����      D  , ,  ]�����  ]����  ^����  ^�����  ]�����      D  , ,  `@����  `@���  `����  `�����  `@����      D  , ,  b�����  b����  c.���  c.����  b�����      D  , ,  _#���C  _#����  _�����  _����C  _#���C      D  , ,  aq���C  aq����  b����  b���C  aq���C      D  , ,  ]����  ]����C  ^����C  ^����  ]����      D  , ,  `@���  `@���C  `����C  `����  `@���      D  , ,  b����  b����C  c.���C  c.���  b����      D  , ,  y����  y����C  z:���C  z:���  y����      D  , ,  {����  {����C  |~���C  |~���  {����      D  , ,  d����  d����C  er���C  er���  d����      D  , ,  g4���  g4���C  g����C  g����  g4���      D  , ,  f���C  f����  f�����  f����C  f���C      D  , ,  h[���C  h[����  h�����  h����C  h[���C      D  , ,  j����C  j�����  k?����  k?���C  j����C      D  , ,  l����C  l�����  m�����  m����C  l����C      D  , ,  oE���C  oE����  o�����  o����C  oE���C      D  , ,  q����C  q�����  r)����  r)���C  q����C      D  , ,  s����C  s�����  tw����  tw���C  s����C      D  , ,  v/���C  v/����  v�����  v����C  v/���C      D  , ,  x}���C  x}����  y����  y���C  x}���C      D  , ,  z����C  z�����  {a����  {a���C  z����C      D  , ,  ix���  ix���C  j���C  j���  ix���      D  , ,  d����m  d����  er���  er���m  d����m      D  , ,  g4���m  g4���  g����  g����m  g4���m      D  , ,  ix���m  ix���  j���  j���m  ix���m      D  , ,  k����m  k����  lf���  lf���m  k����m      D  , ,  n���m  n���  n����  n����m  n���m      D  , ,  pl���m  pl���  q���  q���m  pl���m      D  , ,  k����  k����C  lf���C  lf���  k����      D  , ,  d����-  d�����  er����  er���-  d����-      D  , ,  g4���-  g4����  g�����  g����-  g4���-      D  , ,  ix���-  ix����  j����  j���-  ix���-      D  , ,  k����-  k�����  lf����  lf���-  k����-      D  , ,  n���-  n����  n�����  n����-  n���-      D  , ,  pl���-  pl����  q����  q���-  pl���-      D  , ,  r����-  r�����  sF����  sF���-  r����-      D  , ,  u���-  u����  u�����  u����-  u���-      D  , ,  wL���-  wL����  w�����  w����-  wL���-      D  , ,  y����-  y�����  z:����  z:���-  y����-      D  , ,  {����-  {�����  |~����  |~���-  {����-      D  , ,  n���  n���C  n����C  n����  n���      D  , ,  pl���  pl���C  q���C  q���  pl���      D  , ,  f���  f���  f����  f����  f���      D  , ,  h[���  h[���  h����  h����  h[���      D  , ,  j����  j����  k?���  k?���  j����      D  , ,  l����  l����  m����  m����  l����      D  , ,  d����  d���ݯ  er��ݯ  er���  d����      D  , ,  g4���  g4��ݯ  g���ݯ  g����  g4���      D  , ,  ix���  ix��ݯ  j��ݯ  j���  ix���      D  , ,  k����  k���ݯ  lf��ݯ  lf���  k����      D  , ,  n���  n��ݯ  n���ݯ  n����  n���      D  , ,  pl���  pl��ݯ  q��ݯ  q���  pl���      D  , ,  r����  r���ݯ  sF��ݯ  sF���  r����      D  , ,  u���  u��ݯ  u���ݯ  u����  u���      D  , ,  wL���  wL��ݯ  w���ݯ  w����  wL���      D  , ,  y����  y���ݯ  z:��ݯ  z:���  y����      D  , ,  {����  {���ݯ  |~��ݯ  |~���  {����      D  , ,  oE���  oE���  o����  o����  oE���      D  , ,  q����  q����  r)���  r)���  q����      D  , ,  s����  s����  tw���  tw���  s����      D  , ,  v/���  v/���  v����  v����  v/���      D  , ,  x}���  x}���  y���  y���  x}���      D  , ,  z����  z����  {a���  {a���  z����      D  , ,  r����m  r����  sF���  sF���m  r����m      D  , ,  u���m  u���  u����  u����m  u���m      D  , ,  wL���m  wL���  w����  w����m  wL���m      D  , ,  y����m  y����  z:���  z:���m  y����m      D  , ,  {����m  {����  |~���  |~���m  {����m      D  , ,  r����  r����C  sF���C  sF���  r����      D  , ,  u���  u���C  u����C  u����  u���      D  , ,  wL���  wL���C  w����C  w����  wL���      D  , ,  y����  y����C  z:���C  z:���  y����      D  , ,  {����  {����C  |~���C  |~���  {����      D  , ,  {�����  {����  |~���  |~����  {�����      D  , ,  y�����  y����  z:���  z:����  y�����      D  , ,  d����  d����C  er���C  er���  d����      D  , ,  g4���  g4���C  g����C  g����  g4���      D  , ,  ix���  ix���C  j���C  j���  ix���      D  , ,  k����  k����C  lf���C  lf���  k����      D  , ,  d�����  d����  er���  er����  d�����      D  , ,  g4����  g4���  g����  g�����  g4����      D  , ,  ix����  ix���  j���  j����  ix����      D  , ,  k�����  k����  lf���  lf����  k�����      D  , ,  n����  n���  n����  n�����  n����      D  , ,  pl����  pl���  q���  q����  pl����      D  , ,  r�����  r����  sF���  sF����  r�����      D  , ,  u����  u���  u����  u�����  u����      D  , ,  wL����  wL���  w����  w�����  wL����      D  , ,  n���  n���C  n����C  n����  n���      D  , ,  pl���  pl���C  q���C  q���  pl���      D  , ,  r����  r����C  sF���C  sF���  r����      D  , ,  u���  u���C  u����C  u����  u���      D  , ,  wL���  wL���C  w����C  w����  wL���      D  , ,  d���ڙ  d����/  er���/  er��ڙ  d���ڙ      D  , ,  g4��ڙ  g4���/  g����/  g���ڙ  g4��ڙ      D  , ,  ix��ڙ  ix���/  j���/  j��ڙ  ix��ڙ      D  , ,  k���ڙ  k����/  lf���/  lf��ڙ  k���ڙ      D  , ,  n��ڙ  n���/  n����/  n���ڙ  n��ڙ      D  , ,  pl��ڙ  pl���/  q���/  q��ڙ  pl��ڙ      D  , ,  r���ڙ  r����/  sF���/  sF��ڙ  r���ڙ      D  , ,  u��ڙ  u���/  u����/  u���ڙ  u��ڙ      D  , ,  wL��ڙ  wL���/  w����/  w���ڙ  wL��ڙ      D  , ,  y���ڙ  y����/  z:���/  z:��ڙ  y���ڙ      D  , ,  {���ڙ  {����/  |~���/  |~��ڙ  {���ڙ      D  , ,  d����Y  d�����  er����  er���Y  d����Y      D  , ,  g4���Y  g4����  g�����  g����Y  g4���Y      D  , ,  ix���Y  ix����  j����  j���Y  ix���Y      D  , ,  k����Y  k�����  lf����  lf���Y  k����Y      D  , ,  n���Y  n����  n�����  n����Y  n���Y      D  , ,  pl���Y  pl����  q����  q���Y  pl���Y      D  , ,  r����Y  r�����  sF����  sF���Y  r����Y      D  , ,  u���Y  u����  u�����  u����Y  u���Y      D  , ,  wL���Y  wL����  w�����  w����Y  wL���Y      D  , ,  y����Y  y�����  z:����  z:���Y  y����Y      D  , ,  {����Y  {�����  |~����  |~���Y  {����Y      D  , ,  d����  d���د  er��د  er���  d����      D  , ,  g4���  g4��د  g���د  g����  g4���      D  , ,  ix���  ix��د  j��د  j���  ix���      D  , ,  k����  k���د  lf��د  lf���  k����      D  , ,  n���  n��د  n���د  n����  n���      D  , ,  pl���  pl��د  q��د  q���  pl���      D  , ,  r����  r���د  sF��د  sF���  r����      D  , ,  u���  u��د  u���د  u����  u���      D  , ,  wL���  wL��د  w���د  w����  wL���      D  , ,  y����  y���د  z:��د  z:���  y����      D  , ,  {����  {���د  |~��د  |~���  {����      D  , ,  d�����  d����o  er���o  er����  d�����      D  , ,  d�����  d����o  er���o  er����  d�����      D  , ,  g4����  g4���o  g����o  g�����  g4����      D  , ,  ix����  ix���o  j���o  j����  ix����      D  , ,  k�����  k����o  lf���o  lf����  k�����      D  , ,  n����  n���o  n����o  n�����  n����      D  , ,  pl����  pl���o  q���o  q����  pl����      D  , ,  r�����  r����o  sF���o  sF����  r�����      D  , ,  u����  u���o  u����o  u�����  u����      D  , ,  wL����  wL���o  w����o  w�����  wL����      D  , ,  y�����  y����o  z:���o  z:����  y�����      D  , ,  {�����  {����o  |~���o  |~����  {�����      D  , ,  g4����  g4���o  g����o  g�����  g4����      D  , ,  d���ՙ  d����/  er���/  er��ՙ  d���ՙ      D  , ,  g4��ՙ  g4���/  g����/  g���ՙ  g4��ՙ      D  , ,  ix��ՙ  ix���/  j���/  j��ՙ  ix��ՙ      D  , ,  k���ՙ  k����/  lf���/  lf��ՙ  k���ՙ      D  , ,  n��ՙ  n���/  n����/  n���ՙ  n��ՙ      D  , ,  pl��ՙ  pl���/  q���/  q��ՙ  pl��ՙ      D  , ,  r���ՙ  r����/  sF���/  sF��ՙ  r���ՙ      D  , ,  u��ՙ  u���/  u����/  u���ՙ  u��ՙ      D  , ,  wL��ՙ  wL���/  w����/  w���ՙ  wL��ՙ      D  , ,  y���ՙ  y����/  z:���/  z:��ՙ  y���ՙ      D  , ,  {���ՙ  {����/  |~���/  |~��ՙ  {���ՙ      D  , ,  ix����  ix���o  j���o  j����  ix����      D  , ,  d����Y  d�����  er����  er���Y  d����Y      D  , ,  g4���Y  g4����  g�����  g����Y  g4���Y      D  , ,  ix���Y  ix����  j����  j���Y  ix���Y      D  , ,  k����Y  k�����  lf����  lf���Y  k����Y      D  , ,  n���Y  n����  n�����  n����Y  n���Y      D  , ,  pl���Y  pl����  q����  q���Y  pl���Y      D  , ,  r����Y  r�����  sF����  sF���Y  r����Y      D  , ,  u���Y  u����  u�����  u����Y  u���Y      D  , ,  wL���Y  wL����  w�����  w����Y  wL���Y      D  , ,  y����Y  y�����  z:����  z:���Y  y����Y      D  , ,  {����Y  {�����  |~����  |~���Y  {����Y      D  , ,  k�����  k����o  lf���o  lf����  k�����      D  , ,  g4����  g4���]  g����]  g�����  g4����      D  , ,  k�����  k����]  lf���]  lf����  k�����      D  , ,  pl����  pl���]  q���]  q����  pl����      D  , ,  u����  u���]  u����]  u�����  u����      D  , ,  y�����  y����]  z:���]  z:����  y�����      D  , ,  g4��·  g4���  g����  g���·  g4��·      D  , ,  k���·  k����  lf���  lf��·  k���·      D  , ,  pl��·  pl���  q���  q��·  pl��·      D  , ,  u��·  u���  u����  u���·  u��·      D  , ,  y���·  y����  z:���  z:��·  y���·      D  , ,  n����  n���o  n����o  n�����  n����      D  , ,  pl����  pl���o  q���o  q����  pl����      D  , ,  r�����  r����o  sF���o  sF����  r�����      D  , ,  u����  u���o  u����o  u�����  u����      D  , ,  wL����  wL���o  w����o  w�����  wL����      D  , ,  y�����  y����o  z:���o  z:����  y�����      D  , ,  {�����  {����o  |~���o  |~����  {�����      D  , ,  b�����  b����o  c.���o  c.����  b�����      D  , ,  `@��ڙ  `@���/  `����/  `���ڙ  `@��ڙ      D  , ,  `@����  `@���o  `����o  `�����  `@����      D  , ,  ]����Y  ]�����  ^�����  ^����Y  ]����Y      D  , ,  ]�����  ]����]  ^����]  ^�����  ]�����      D  , ,  b�����  b����]  c.���]  c.����  b�����      D  , ,  `@���Y  `@����  `�����  `����Y  `@���Y      D  , ,  b����Y  b�����  c.����  c.���Y  b����Y      D  , ,  b���ڙ  b����/  c.���/  c.��ڙ  b���ڙ      D  , ,  ]�����  ]����o  ^����o  ^�����  ]�����      D  , ,  ]���ڙ  ]����/  ^����/  ^���ڙ  ]���ڙ      D  , ,  ]���·  ]����  ^����  ^���·  ]���·      D  , ,  b���·  b����  c.���  c.��·  b���·      D  , ,  b�����  b����o  c.���o  c.����  b�����      D  , ,  ]����Y  ]�����  ^�����  ^����Y  ]����Y      D  , ,  `@���Y  `@����  `�����  `����Y  `@���Y      D  , ,  b����Y  b�����  c.����  c.���Y  b����Y      D  , ,  ]����  ]���د  ^���د  ^����  ]����      D  , ,  `@���  `@��د  `���د  `����  `@���      D  , ,  b����  b���د  c.��د  c.���  b����      D  , ,  ]���ՙ  ]����/  ^����/  ^���ՙ  ]���ՙ      D  , ,  `@��ՙ  `@���/  `����/  `���ՙ  `@��ՙ      D  , ,  b���ՙ  b����/  c.���/  c.��ՙ  b���ՙ      D  , ,  ]�����  ]����o  ^����o  ^�����  ]�����      D  , ,  `@����  `@���o  `����o  `�����  `@����      D  , ,  ]����G  ]�����  ^�����  ^����G  ]����G      D  , ,  ]����#  ]���Ĺ  ^���Ĺ  ^����#  ]����#      D  , ,  `T���#  `T��Ĺ  `���Ĺ  `����#  `T���#      D  , ,  b����#  b���Ĺ  c.��Ĺ  c.���#  b����#      D  , ,  b����G  b�����  c.����  c.���G  b����G      D  , ,  ]�����  ]����y  ^����y  ^�����  ]�����      D  , ,  `T����  `T���y  `����y  `�����  `T����      D  , ,  b�����  b����y  c.���y  c.����  b�����      D  , ,  ]����  ]���̝  ^���̝  ^����  ]����      D  , ,  ]�����  ]����9  ^����9  ^�����  ]�����      D  , ,  `T����  `T���9  `����9  `�����  `T����      D  , ,  b�����  b����9  c.���9  c.����  b�����      D  , ,  b����  b���̝  c.��̝  c.���  b����      D  , ,  ]����c  ]�����  ^�����  ^����c  ]����c      D  , ,  `T���c  `T����  `�����  `����c  `T���c      D  , ,  b����c  b�����  c.����  c.���c  b����c      D  , ,  ]����c  ]�����  ^�����  ^����c  ]����c      D  , ,  `T���c  `T����  `�����  `����c  `T���c      D  , ,  b����c  b�����  c.����  c.���c  b����c      D  , ,  y����c  y�����  z:����  z:���c  y����c      D  , ,  {����c  {�����  |�����  |����c  {����c      D  , ,  g4���G  g4����  g�����  g����G  g4���G      D  , ,  k����G  k�����  lf����  lf���G  k����G      D  , ,  g4���  g4��̝  g���̝  g����  g4���      D  , ,  k����  k���̝  lf��̝  lf���  k����      D  , ,  d����#  d���Ĺ  e���Ĺ  e����#  d����#      D  , ,  g4���#  g4��Ĺ  g���Ĺ  g����#  g4���#      D  , ,  i����#  i���Ĺ  j"��Ĺ  j"���#  i����#      D  , ,  k����#  k���Ĺ  lf��Ĺ  lf���#  k����#      D  , ,  n(���#  n(��Ĺ  n���Ĺ  n����#  n(���#      D  , ,  pl���#  pl��Ĺ  q��Ĺ  q���#  pl���#      D  , ,  r����#  r���Ĺ  sZ��Ĺ  sZ���#  r����#      D  , ,  u���#  u��Ĺ  u���Ĺ  u����#  u���#      D  , ,  w`���#  w`��Ĺ  w���Ĺ  w����#  w`���#      D  , ,  y����#  y���Ĺ  z:��Ĺ  z:���#  y����#      D  , ,  {����#  {���Ĺ  |���Ĺ  |����#  {����#      D  , ,  pl���  pl��̝  q��̝  q���  pl���      D  , ,  u���  u��̝  u���̝  u����  u���      D  , ,  y����  y���̝  z:��̝  z:���  y����      D  , ,  pl���G  pl����  q����  q���G  pl���G      D  , ,  d�����  d����y  e����y  e�����  d�����      D  , ,  g4����  g4���y  g����y  g�����  g4����      D  , ,  i�����  i����y  j"���y  j"����  i�����      D  , ,  k�����  k����y  lf���y  lf����  k�����      D  , ,  n(����  n(���y  n����y  n�����  n(����      D  , ,  pl����  pl���y  q���y  q����  pl����      D  , ,  r�����  r����y  sZ���y  sZ����  r�����      D  , ,  u����  u���y  u����y  u�����  u����      D  , ,  w`����  w`���y  w����y  w�����  w`����      D  , ,  y�����  y����y  z:���y  z:����  y�����      D  , ,  {�����  {����y  |����y  |�����  {�����      D  , ,  u���G  u����  u�����  u����G  u���G      D  , ,  y����G  y�����  z:����  z:���G  y����G      D  , ,  d����c  d�����  e�����  e����c  d����c      D  , ,  g4���c  g4����  g�����  g����c  g4���c      D  , ,  d�����  d����9  e����9  e�����  d�����      D  , ,  g4����  g4���9  g����9  g�����  g4����      D  , ,  i�����  i����9  j"���9  j"����  i�����      D  , ,  k�����  k����9  lf���9  lf����  k�����      D  , ,  n(����  n(���9  n����9  n�����  n(����      D  , ,  pl����  pl���9  q���9  q����  pl����      D  , ,  r�����  r����9  sZ���9  sZ����  r�����      D  , ,  u����  u���9  u����9  u�����  u����      D  , ,  w`����  w`���9  w����9  w�����  w`����      D  , ,  y�����  y����9  z:���9  z:����  y�����      D  , ,  {�����  {����9  |����9  |�����  {�����      D  , ,  i����c  i�����  j"����  j"���c  i����c      D  , ,  k����c  k�����  lf����  lf���c  k����c      D  , ,  n(���c  n(����  n�����  n����c  n(���c      D  , ,  pl���c  pl����  q����  q���c  pl���c      D  , ,  d����c  d�����  e�����  e����c  d����c      D  , ,  g4���c  g4����  g�����  g����c  g4���c      D  , ,  i����c  i�����  j"����  j"���c  i����c      D  , ,  k����c  k�����  lf����  lf���c  k����c      D  , ,  n(���c  n(����  n�����  n����c  n(���c      D  , ,  pl���c  pl����  q����  q���c  pl���c      D  , ,  r����c  r�����  sZ����  sZ���c  r����c      D  , ,  u���c  u����  u�����  u����c  u���c      D  , ,  w`���c  w`����  w�����  w����c  w`���c      D  , ,  y����c  y�����  z:����  z:���c  y����c      D  , ,  {����c  {�����  |�����  |����c  {����c      D  , ,  r����c  r�����  sZ����  sZ���c  r����c      D  , ,  u���c  u����  u�����  u����c  u���c      D  , ,  w`���c  w`����  w�����  w����c  w`���c      D  , ,  � ��ՙ  � ���/  �����/  ����ՙ  � ��ՙ      D  , ,  �d��ՙ  �d���/  �����/  ����ՙ  �d��ՙ      D  , ,  ����ՙ  �����/  �R���/  �R��ՙ  ����ՙ      D  , ,  � ��ՙ  � ���/  �����/  ����ՙ  � ��ՙ      D  , ,  �X��ՙ  �X���/  �����/  ����ՙ  �X��ՙ      D  , ,  �����Y  ������  �&����  �&���Y  �����Y      D  , ,  �����Y  ������  �~����  �~���Y  �����Y      D  , ,  �,���Y  �,����  ������  �����Y  �,���Y      D  , ,  �����Y  ������  �����  ����Y  �����Y      D  , ,  �����Y  ������  �^����  �^���Y  �����Y      D  , ,  � ���Y  � ����  ������  �����Y  � ���Y      D  , ,  �d���Y  �d����  ������  �����Y  �d���Y      D  , ,  �����Y  ������  �&����  �&���Y  �����Y      D  , ,  �����Y  ������  �~����  �~���Y  �����Y      D  , ,  �,���Y  �,����  ������  �����Y  �,���Y      D  , ,  �����Y  ������  �����  ����Y  �����Y      D  , ,  �����Y  ������  �^����  �^���Y  �����Y      D  , ,  � ���Y  � ����  ������  �����Y  � ���Y      D  , ,  �d���Y  �d����  ������  �����Y  �d���Y      D  , ,  �����Y  ������  �R����  �R���Y  �����Y      D  , ,  � ���Y  � ����  ������  �����Y  � ���Y      D  , ,  �X���Y  �X����  ������  �����Y  �X���Y      D  , ,  �����Y  ������  �R����  �R���Y  �����Y      D  , ,  � ���Y  � ����  ������  �����Y  � ���Y      D  , ,  �X���Y  �X����  ������  �����Y  �X���Y      D  , ,  ������  �����o  �&���o  �&����  ������      D  , ,  ������  �����o  �~���o  �~����  ������      D  , ,  �,����  �,���o  �����o  ������  �,����      D  , ,  ������  �����]  �~���]  �~����  ������      D  , ,  ������  �����]  ����]  �����  ������      D  , ,  � ����  � ���]  �����]  ������  � ����      D  , ,  ������  �����]  �R���]  �R����  ������      D  , ,  �X����  �X���]  �����]  ������  �X����      D  , ,  ������  �����o  ����o  �����  ������      D  , ,  ����·  �����  �~���  �~��·  ����·      D  , ,  ����·  �����  ����  ���·  ����·      D  , ,  � ��·  � ���  �����  ����·  � ��·      D  , ,  ����·  �����  �R���  �R��·  ����·      D  , ,  �X��·  �X���  �����  ����·  �X��·      D  , ,  �����  ����د  �&��د  �&���  �����      D  , ,  �����  ����د  �~��د  �~���  �����      D  , ,  �,���  �,��د  ����د  �����  �,���      D  , ,  �����  ����د  ���د  ����  �����      D  , ,  �����  ����د  �^��د  �^���  �����      D  , ,  � ���  � ��د  ����د  �����  � ���      D  , ,  �d���  �d��د  ����د  �����  �d���      D  , ,  �����  ����د  �R��د  �R���  �����      D  , ,  � ���  � ��د  ����د  �����  � ���      D  , ,  �X���  �X��د  ����د  �����  �X���      D  , ,  ����ڙ  �����/  �&���/  �&��ڙ  ����ڙ      D  , ,  ����ڙ  �����/  �~���/  �~��ڙ  ����ڙ      D  , ,  �,��ڙ  �,���/  �����/  ����ڙ  �,��ڙ      D  , ,  ����ڙ  �����/  ����/  ���ڙ  ����ڙ      D  , ,  ����ڙ  �����/  �^���/  �^��ڙ  ����ڙ      D  , ,  � ��ڙ  � ���/  �����/  ����ڙ  � ��ڙ      D  , ,  �d��ڙ  �d���/  �����/  ����ڙ  �d��ڙ      D  , ,  ����ڙ  �����/  �R���/  �R��ڙ  ����ڙ      D  , ,  � ��ڙ  � ���/  �����/  ����ڙ  � ��ڙ      D  , ,  �X��ڙ  �X���/  �����/  ����ڙ  �X��ڙ      D  , ,  ������  �����o  �^���o  �^����  ������      D  , ,  � ����  � ���o  �����o  ������  � ����      D  , ,  �d����  �d���o  �����o  ������  �d����      D  , ,  ������  �����o  �&���o  �&����  ������      D  , ,  ������  �����o  �~���o  �~����  ������      D  , ,  �,����  �,���o  �����o  ������  �,����      D  , ,  ������  �����o  ����o  �����  ������      D  , ,  ������  �����o  �^���o  �^����  ������      D  , ,  � ����  � ���o  �����o  ������  � ����      D  , ,  �d����  �d���o  �����o  ������  �d����      D  , ,  ������  �����o  �R���o  �R����  ������      D  , ,  � ����  � ���o  �����o  ������  � ����      D  , ,  �X����  �X���o  �����o  ������  �X����      D  , ,  ������  �����o  �R���o  �R����  ������      D  , ,  � ����  � ���o  �����o  ������  � ����      D  , ,  �X����  �X���o  �����o  ������  �X����      D  , ,  ����ՙ  �����/  �&���/  �&��ՙ  ����ՙ      D  , ,  ����ՙ  �����/  �~���/  �~��ՙ  ����ՙ      D  , ,  �,��ՙ  �,���/  �����/  ����ՙ  �,��ՙ      D  , ,  ����ՙ  �����/  ����/  ���ՙ  ����ՙ      D  , ,  ����ՙ  �����/  �^���/  �^��ՙ  ����ՙ      D  , ,  ����ڙ  �����/  �F���/  �F��ڙ  ����ڙ      D  , ,  ~@���  ~@��د  ~���د  ~����  ~@���      D  , ,  �����  ����د  ���د  ����  �����      D  , ,  �����  ����د  �r��د  �r���  �����      D  , ,  � ���  � ��د  ����د  �����  � ���      D  , ,  �x���  �x��د  ���د  ����  �x���      D  , ,  �����  ����د  �R��د  �R���  �����      D  , ,  ����  ���د  ����د  �����  ����      D  , ,  �X���  �X��د  ����د  �����  �X���      D  , ,  �����  ����د  �F��د  �F���  �����      D  , ,  �����  ����د  ����د  �����  �����      D  , ,  �L���  �L��د  ����د  �����  �L���      D  , ,  ~@���Y  ~@����  ~�����  ~����Y  ~@���Y      D  , ,  �����Y  ������  �����  ����Y  �����Y      D  , ,  �����Y  ������  �r����  �r���Y  �����Y      D  , ,  � ���Y  � ����  ������  �����Y  � ���Y      D  , ,  �x���Y  �x����  �����  ����Y  �x���Y      D  , ,  ������  �����o  �����o  ������  ������      D  , ,  �L����  �L���o  �����o  ������  �L����      D  , ,  �����Y  ������  �R����  �R���Y  �����Y      D  , ,  ����Y  �����  ������  �����Y  ����Y      D  , ,  �X���Y  �X����  ������  �����Y  �X���Y      D  , ,  ����ڙ  �����/  �����/  ����ڙ  ����ڙ      D  , ,  �L��ڙ  �L���/  �����/  ����ڙ  �L��ڙ      D  , ,  ~@����  ~@���]  ~����]  ~�����  ~@����      D  , ,  ������  �����]  �r���]  �r����  ������      D  , ,  �x����  �x���]  ����]  �����  �x����      D  , ,  �����  ����]  �����]  ������  �����      D  , ,  ������  �����]  �F���]  �F����  ������      D  , ,  �L����  �L���]  �����]  ������  �L����      D  , ,  �����Y  ������  �F����  �F���Y  �����Y      D  , ,  �����Y  ������  ������  �����Y  �����Y      D  , ,  �L���Y  �L����  ������  �����Y  �L���Y      D  , ,  �L���Y  �L����  ������  �����Y  �L���Y      D  , ,  � ���Y  � ����  ������  �����Y  � ���Y      D  , ,  �x���Y  �x����  �����  ����Y  �x���Y      D  , ,  ~@��ڙ  ~@���/  ~����/  ~���ڙ  ~@��ڙ      D  , ,  ~@����  ~@���o  ~����o  ~�����  ~@����      D  , ,  ������  �����o  ����o  �����  ������      D  , ,  ������  �����o  �r���o  �r����  ������      D  , ,  � ����  � ���o  �����o  ������  � ����      D  , ,  �x����  �x���o  ����o  �����  �x����      D  , ,  ������  �����o  �R���o  �R����  ������      D  , ,  �����  ����o  �����o  ������  �����      D  , ,  �X����  �X���o  �����o  ������  �X����      D  , ,  ������  �����o  �F���o  �F����  ������      D  , ,  ������  �����o  �����o  ������  ������      D  , ,  �L����  �L���o  �����o  ������  �L����      D  , ,  ����ڙ  �����/  ����/  ���ڙ  ����ڙ      D  , ,  ����ڙ  �����/  �r���/  �r��ڙ  ����ڙ      D  , ,  � ��ڙ  � ���/  �����/  ����ڙ  � ��ڙ      D  , ,  �x��ڙ  �x���/  ����/  ���ڙ  �x��ڙ      D  , ,  ����ڙ  �����/  �R���/  �R��ڙ  ����ڙ      D  , ,  ~@��·  ~@���  ~����  ~���·  ~@��·      D  , ,  ����·  �����  �r���  �r��·  ����·      D  , ,  �x��·  �x���  ����  ���·  �x��·      D  , ,  ���·  ����  �����  ����·  ���·      D  , ,  ����·  �����  �F���  �F��·  ����·      D  , ,  �L��·  �L���  �����  ����·  �L��·      D  , ,  �����Y  ������  �R����  �R���Y  �����Y      D  , ,  ����Y  �����  ������  �����Y  ����Y      D  , ,  ~@����  ~@���o  ~����o  ~�����  ~@����      D  , ,  ������  �����o  ����o  �����  ������      D  , ,  ������  �����o  �r���o  �r����  ������      D  , ,  � ����  � ���o  �����o  ������  � ����      D  , ,  �x����  �x���o  ����o  �����  �x����      D  , ,  ������  �����o  �R���o  �R����  ������      D  , ,  �����  ����o  �����o  ������  �����      D  , ,  �X����  �X���o  �����o  ������  �X����      D  , ,  ������  �����o  �F���o  �F����  ������      D  , ,  ~@���Y  ~@����  ~�����  ~����Y  ~@���Y      D  , ,  �����Y  ������  �����  ����Y  �����Y      D  , ,  �����Y  ������  �r����  �r���Y  �����Y      D  , ,  ~@��ՙ  ~@���/  ~����/  ~���ՙ  ~@��ՙ      D  , ,  ����ՙ  �����/  ����/  ���ՙ  ����ՙ      D  , ,  ����ՙ  �����/  �r���/  �r��ՙ  ����ՙ      D  , ,  � ��ՙ  � ���/  �����/  ����ՙ  � ��ՙ      D  , ,  �x��ՙ  �x���/  ����/  ���ՙ  �x��ՙ      D  , ,  ����ՙ  �����/  �R���/  �R��ՙ  ����ՙ      D  , ,  ���ՙ  ����/  �����/  ����ՙ  ���ՙ      D  , ,  �X��ՙ  �X���/  �����/  ����ՙ  �X��ՙ      D  , ,  ����ՙ  �����/  �F���/  �F��ՙ  ����ՙ      D  , ,  ����ՙ  �����/  �����/  ����ՙ  ����ՙ      D  , ,  �L��ՙ  �L���/  �����/  ����ՙ  �L��ՙ      D  , ,  �X���Y  �X����  ������  �����Y  �X���Y      D  , ,  �����Y  ������  �F����  �F���Y  �����Y      D  , ,  �����Y  ������  ������  �����Y  �����Y      D  , ,  ���ڙ  ����/  �����/  ����ڙ  ���ڙ      D  , ,  �X��ڙ  �X���/  �����/  ����ڙ  �X��ڙ      D  , ,  �x���  �x��̝  ���̝  ����  �x���      D  , ,  ~@����  ~@���y  ~����y  ~�����  ~@����      D  , ,  ������  �����y  �.���y  �.����  ������      D  , ,  ������  �����y  �r���y  �r����  ������      D  , ,  �4����  �4���y  �����y  ������  �4����      D  , ,  �x����  �x���y  ����y  �����  �x����      D  , ,  ������  �����y  �f���y  �f����  ������      D  , ,  �����  ����y  �����y  ������  �����      D  , ,  �l����  �l���y  ����y  �����  �l����      D  , ,  ������  �����y  �F���y  �F����  ������      D  , ,  �����  ����y  �����y  ������  �����      D  , ,  �L����  �L���y  �����y  ������  �L����      D  , ,  ����  ���̝  ����̝  �����  ����      D  , ,  �����  ����̝  �F��̝  �F���  �����      D  , ,  �L���  �L��̝  ����̝  �����  �L���      D  , ,  �����G  ������  �r����  �r���G  �����G      D  , ,  �x���G  �x����  �����  ����G  �x���G      D  , ,  ~@���c  ~@����  ~�����  ~����c  ~@���c      D  , ,  �����c  ������  �.����  �.���c  �����c      D  , ,  �����c  ������  �r����  �r���c  �����c      D  , ,  ~@���#  ~@��Ĺ  ~���Ĺ  ~����#  ~@���#      D  , ,  �����#  ����Ĺ  �.��Ĺ  �.���#  �����#      D  , ,  �����#  ����Ĺ  �r��Ĺ  �r���#  �����#      D  , ,  �4���#  �4��Ĺ  ����Ĺ  �����#  �4���#      D  , ,  �x���#  �x��Ĺ  ���Ĺ  ����#  �x���#      D  , ,  �����#  ����Ĺ  �f��Ĺ  �f���#  �����#      D  , ,  ����#  ���Ĺ  ����Ĺ  �����#  ����#      D  , ,  ~@����  ~@���9  ~����9  ~�����  ~@����      D  , ,  ������  �����9  �.���9  �.����  ������      D  , ,  ������  �����9  �r���9  �r����  ������      D  , ,  �4����  �4���9  �����9  ������  �4����      D  , ,  �x����  �x���9  ����9  �����  �x����      D  , ,  ������  �����9  �f���9  �f����  ������      D  , ,  �����  ����9  �����9  ������  �����      D  , ,  �l����  �l���9  ����9  �����  �l����      D  , ,  ������  �����9  �F���9  �F����  ������      D  , ,  �����  ����9  �����9  ������  �����      D  , ,  �L����  �L���9  �����9  ������  �L����      D  , ,  �l���#  �l��Ĺ  ���Ĺ  ����#  �l���#      D  , ,  �����#  ����Ĺ  �F��Ĺ  �F���#  �����#      D  , ,  ����#  ���Ĺ  ����Ĺ  �����#  ����#      D  , ,  �L���#  �L��Ĺ  ����Ĺ  �����#  �L���#      D  , ,  �4���c  �4����  ������  �����c  �4���c      D  , ,  �x���c  �x����  �����  ����c  �x���c      D  , ,  �����c  ������  �f����  �f���c  �����c      D  , ,  ����c  �����  ������  �����c  ����c      D  , ,  �l���c  �l����  �����  ����c  �l���c      D  , ,  �����c  ������  �F����  �F���c  �����c      D  , ,  ����c  �����  ������  �����c  ����c      D  , ,  �L���c  �L����  ������  �����c  �L���c      D  , ,  ����G  �����  ������  �����G  ����G      D  , ,  �����G  ������  �F����  �F���G  �����G      D  , ,  �L���G  �L����  ������  �����G  �L���G      D  , ,  ~@���c  ~@����  ~�����  ~����c  ~@���c      D  , ,  �����c  ������  �.����  �.���c  �����c      D  , ,  �����c  ������  �r����  �r���c  �����c      D  , ,  �4���c  �4����  ������  �����c  �4���c      D  , ,  �x���c  �x����  �����  ����c  �x���c      D  , ,  �����c  ������  �f����  �f���c  �����c      D  , ,  ����c  �����  ������  �����c  ����c      D  , ,  �l���c  �l����  �����  ����c  �l���c      D  , ,  �����c  ������  �F����  �F���c  �����c      D  , ,  ����c  �����  ������  �����c  ����c      D  , ,  �L���c  �L����  ������  �����c  �L���c      D  , ,  ~@���G  ~@����  ~�����  ~����G  ~@���G      D  , ,  ~@���  ~@��̝  ~���̝  ~����  ~@���      D  , ,  �����  ����̝  �r��̝  �r���  �����      D  , ,  �����c  ������  �R����  �R���c  �����c      D  , ,  ����c  �����  ������  �����c  ����c      D  , ,  �X���c  �X����  ������  �����c  �X���c      D  , ,  �����  ����̝  �~��̝  �~���  �����      D  , ,  �����  ����̝  ���̝  ����  �����      D  , ,  � ���  � ��̝  ����̝  �����  � ���      D  , ,  �����  ����̝  �R��̝  �R���  �����      D  , ,  �X���  �X��̝  ����̝  �����  �X���      D  , ,  �����G  ������  �R����  �R���G  �����G      D  , ,  �����#  ����Ĺ  �:��Ĺ  �:���#  �����#      D  , ,  �����#  ����Ĺ  �~��Ĺ  �~���#  �����#      D  , ,  ������  �����9  �:���9  �:����  ������      D  , ,  ������  �����9  �~���9  �~����  ������      D  , ,  �@����  �@���9  �����9  ������  �@����      D  , ,  ������  �����9  ����9  �����  ������      D  , ,  ������  �����9  �r���9  �r����  ������      D  , ,  � ����  � ���9  �����9  ������  � ����      D  , ,  �x����  �x���9  ����9  �����  �x����      D  , ,  ������  �����9  �R���9  �R����  ������      D  , ,  �����  ����9  �����9  ������  �����      D  , ,  �X����  �X���9  �����9  ������  �X����      D  , ,  �@���#  �@��Ĺ  ����Ĺ  �����#  �@���#      D  , ,  �����#  ����Ĺ  ���Ĺ  ����#  �����#      D  , ,  �����#  ����Ĺ  �r��Ĺ  �r���#  �����#      D  , ,  � ���#  � ��Ĺ  ����Ĺ  �����#  � ���#      D  , ,  ������  �����y  �:���y  �:����  ������      D  , ,  ������  �����y  �~���y  �~����  ������      D  , ,  �@����  �@���y  �����y  ������  �@����      D  , ,  ������  �����y  ����y  �����  ������      D  , ,  ������  �����y  �r���y  �r����  ������      D  , ,  � ����  � ���y  �����y  ������  � ����      D  , ,  �x����  �x���y  ����y  �����  �x����      D  , ,  ������  �����y  �R���y  �R����  ������      D  , ,  �����  ����y  �����y  ������  �����      D  , ,  �X����  �X���y  �����y  ������  �X����      D  , ,  �x���#  �x��Ĺ  ���Ĺ  ����#  �x���#      D  , ,  �����#  ����Ĺ  �R��Ĺ  �R���#  �����#      D  , ,  ����#  ���Ĺ  ����Ĺ  �����#  ����#      D  , ,  �X���#  �X��Ĺ  ����Ĺ  �����#  �X���#      D  , ,  �X���G  �X����  ������  �����G  �X���G      D  , ,  �����G  ������  �~����  �~���G  �����G      D  , ,  �����G  ������  �����  ����G  �����G      D  , ,  � ���G  � ����  ������  �����G  � ���G      D  , ,  �����c  ������  �:����  �:���c  �����c      D  , ,  �����c  ������  �~����  �~���c  �����c      D  , ,  �@���c  �@����  ������  �����c  �@���c      D  , ,  �����c  ������  �����  ����c  �����c      D  , ,  �����c  ������  �:����  �:���c  �����c      D  , ,  �����c  ������  �~����  �~���c  �����c      D  , ,  �@���c  �@����  ������  �����c  �@���c      D  , ,  �����c  ������  �����  ����c  �����c      D  , ,  �����c  ������  �r����  �r���c  �����c      D  , ,  � ���c  � ����  ������  �����c  � ���c      D  , ,  �x���c  �x����  �����  ����c  �x���c      D  , ,  �����c  ������  �R����  �R���c  �����c      D  , ,  ����c  �����  ������  �����c  ����c      D  , ,  �X���c  �X����  ������  �����c  �X���c      D  , ,  �����c  ������  �r����  �r���c  �����c      D  , ,  � ���c  � ����  ������  �����c  � ���c      D  , ,  �x���c  �x����  �����  ����c  �x���c      D  , ,  � ���m  � ���  Ȗ���  Ȗ���m  � ���m      D  , ,  � ����  � ���  Ȗ���  Ȗ����  � ����      D  , ,  � ���  � ���C  Ȗ���C  Ȗ���  � ���      D  , ,  �D����  �D���  �����  ������  �D����      D  , ,  ̜����  ̜���  �2���  �2����  ̜����      D  , ,  ������  �����  �v���  �v����  ������      D  , ,  �8����  �8���  �����  ������  �8����      D  , ,  � ���  � ����  Ȗ����  Ȗ���  � ���      D  , ,  � ���Q  � ����  Ȗ����  Ȗ���Q  � ���Q      D  , ,  � ���-  � ����  Ȗ����  Ȗ���-  � ���-      D  , ,  � ���-  � ����  Ȗ����  Ȗ���-  � ���-      D  , ,  � ���m  � ���  Ȗ���  Ȗ���m  � ���m      D  , ,  � ���  � ���C  Ȗ���C  Ȗ���  � ���      D  , ,  � ����  � ���g  Ȗ���g  Ȗ����  � ����      D  , ,  � ����  � ���'  Ȗ���'  Ȗ����  � ����      D  , ,  � ����  � ���  Ȗ���  Ȗ����  � ����      D  , ,  � ���  � ��ݯ  Ȗ��ݯ  Ȗ���  � ���      D  , ,  ������  �����  �����  ������  ������      D  , ,  �8����  �8���  �����  ������  �8����      D  , ,  ������  �����  �&���  �&����  ������      D  , ,  ������  �����  �j���  �j����  ������      D  , ,  �,����  �,���  �����  ������  �,����      D  , ,  �p����  �p���  ����  �����  �p����      D  , ,  ������  �����  �^���  �^����  ������      D  , ,  �����  ����  �����  ������  �����      D  , ,  �d����  �d���  �����  ������  �d����      D  , ,  Ũ����  Ũ���  �>���  �>����  Ũ����      D  , ,  �8����  �8���g  �����g  ������  �8����      D  , ,  �����-  ������  �v����  �v���-  �����-      D  , ,  ̜����  ̜���'  �2���'  �2����  ̜����      D  , ,  �8���-  �8����  ������  �����-  �8���-      D  , ,  �8����  �8���'  �����'  ������  �8����      D  , ,  ̜���  ̜����  �2����  �2���  ̜���      D  , ,  �8���  �8����  ������  �����  �8���      D  , ,  �D���m  �D���  �����  �����m  �D���m      D  , ,  ̜���m  ̜���  �2���  �2���m  ̜���m      D  , ,  �����m  �����  �v���  �v���m  �����m      D  , ,  �D���-  �D����  ������  �����-  �D���-      D  , ,  �8���m  �8���  �����  �����m  �8���m      D  , ,  ̜���Q  ̜����  �2����  �2���Q  ̜���Q      D  , ,  �8���Q  �8����  ������  �����Q  �8���Q      D  , ,  ̜���-  ̜����  �2����  �2���-  ̜���-      D  , ,  ̜����  ̜���g  �2���g  �2����  ̜����      D  , ,  �����-  ������  �&����  �&���-  �����-      D  , ,  �����-  ������  �j����  �j���-  �����-      D  , ,  �,���-  �,����  ������  �����-  �,���-      D  , ,  �p���-  �p����  �����  ����-  �p���-      D  , ,  �����-  ������  �^����  �^���-  �����-      D  , ,  �d����  �d���g  �����g  ������  �d����      D  , ,  ����-  �����  ������  �����-  ����-      D  , ,  �d���-  �d����  ������  �����-  �d���-      D  , ,  Ũ���-  Ũ����  �>����  �>���-  Ũ���-      D  , ,  ������  �����g  �����g  ������  ������      D  , ,  ������  �����g  �&���g  �&����  ������      D  , ,  ������  �����'  �����'  ������  ������      D  , ,  ������  �����'  �&���'  �&����  ������      D  , ,  �,����  �,���'  �����'  ������  �,����      D  , ,  ������  �����'  �^���'  �^����  ������      D  , ,  �d����  �d���'  �����'  ������  �d����      D  , ,  �����Q  ������  �^����  �^���Q  �����Q      D  , ,  �d���Q  �d����  ������  �����Q  �d���Q      D  , ,  �,���Q  �,����  ������  �����Q  �,���Q      D  , ,  �����m  �����  �����  �����m  �����m      D  , ,  �,����  �,���g  �����g  ������  �,����      D  , ,  ������  �����g  �^���g  �^����  ������      D  , ,  �����Q  ������  ������  �����Q  �����Q      D  , ,  �����Q  ������  �&����  �&���Q  �����Q      D  , ,  �8���m  �8���  �����  �����m  �8���m      D  , ,  �����  ������  ������  �����  �����      D  , ,  �����  ������  �&����  �&���  �����      D  , ,  �,���  �,����  ������  �����  �,���      D  , ,  �����  ������  �^����  �^���  �����      D  , ,  �d���  �d����  ������  �����  �d���      D  , ,  �,���m  �,���  �����  �����m  �,���m      D  , ,  �p���m  �p���  ����  ����m  �p���m      D  , ,  �����m  �����  �^���  �^���m  �����m      D  , ,  ����m  ����  �����  �����m  ����m      D  , ,  �d���m  �d���  �����  �����m  �d���m      D  , ,  �����m  �����  �&���  �&���m  �����m      D  , ,  Ũ���m  Ũ���  �>���  �>���m  Ũ���m      D  , ,  �����m  �����  �j���  �j���m  �����m      D  , ,  �����-  ������  ������  �����-  �����-      D  , ,  �8���-  �8����  ������  �����-  �8���-      D  , ,  �p���  �p���C  ����C  ����  �p���      D  , ,  �����  �����C  �^���C  �^���  �����      D  , ,  ����  ����C  �����C  �����  ����      D  , ,  �d���  �d���C  �����C  �����  �d���      D  , ,  Ũ���  Ũ���C  �>���C  �>���  Ũ���      D  , ,  �����  �����C  �����C  �����  �����      D  , ,  �����C  ������  �c����  �c���C  �����C      D  , ,  ����C  �����  ������  �����C  ����C      D  , ,  �i���C  �i����  ������  �����C  �i���C      D  , ,  �����C  ������  �M����  �M���C  �����C      D  , ,  ����C  �����  ������  �����C  ����C      D  , ,  �S���C  �S����  ������  �����C  �S���C      D  , ,  �����C  ������  �7����  �7���C  �����C      D  , ,  �����C  ������  ������  �����C  �����C      D  , ,  �=���C  �=����  ������  �����C  �=���C      D  , ,  ċ���C  ċ����  �!����  �!���C  ċ���C      D  , ,  �����C  ������  �o����  �o���C  �����C      D  , ,  �8���  �8���C  �����C  �����  �8���      D  , ,  �����  �����C  �&���C  �&���  �����      D  , ,  �����  �����C  �j���C  �j���  �����      D  , ,  �,���  �,���C  �����C  �����  �,���      D  , ,  �p���  �p���C  ����C  ����  �p���      D  , ,  �����  �����C  �^���C  �^���  �����      D  , ,  �����  �����  �c���  �c���  �����      D  , ,  ����  ����  �����  �����  ����      D  , ,  �i���  �i���  �����  �����  �i���      D  , ,  �����  �����  �M���  �M���  �����      D  , ,  ����  ����  �����  �����  ����      D  , ,  �S���  �S���  �����  �����  �S���      D  , ,  �����  �����  �7���  �7���  �����      D  , ,  �����  �����  �����  �����  �����      D  , ,  �=���  �=���  �����  �����  �=���      D  , ,  ċ���  ċ���  �!���  �!���  ċ���      D  , ,  ������  �����  �����  ������  ������      D  , ,  �8����  �8���  �����  ������  �8����      D  , ,  ������  �����  �&���  �&����  ������      D  , ,  ������  �����  �j���  �j����  ������      D  , ,  �,����  �,���  �����  ������  �,����      D  , ,  �p����  �p���  ����  �����  �p����      D  , ,  ������  �����  �^���  �^����  ������      D  , ,  �����  ����  �����  ������  �����      D  , ,  �d����  �d���  �����  ������  �d����      D  , ,  Ũ����  Ũ���  �>���  �>����  Ũ����      D  , ,  �����  �����  �o���  �o���  �����      D  , ,  �����-  ������  ������  �����-  �����-      D  , ,  �8���-  �8����  ������  �����-  �8���-      D  , ,  �����-  ������  �&����  �&���-  �����-      D  , ,  �����-  ������  �j����  �j���-  �����-      D  , ,  �,���-  �,����  ������  �����-  �,���-      D  , ,  �����  ����ݯ  ����ݯ  �����  �����      D  , ,  �8���  �8��ݯ  ����ݯ  �����  �8���      D  , ,  �����  ����ݯ  �&��ݯ  �&���  �����      D  , ,  �����  ����ݯ  �j��ݯ  �j���  �����      D  , ,  �,���  �,��ݯ  ����ݯ  �����  �,���      D  , ,  �p���  �p��ݯ  ���ݯ  ����  �p���      D  , ,  �����  ����ݯ  �^��ݯ  �^���  �����      D  , ,  ����  ���ݯ  ����ݯ  �����  ����      D  , ,  �d���  �d��ݯ  ����ݯ  �����  �d���      D  , ,  Ũ���  Ũ��ݯ  �>��ݯ  �>���  Ũ���      D  , ,  �p���-  �p����  �����  ����-  �p���-      D  , ,  �����-  ������  �^����  �^���-  �����-      D  , ,  ����-  �����  ������  �����-  ����-      D  , ,  �d���-  �d����  ������  �����-  �d���-      D  , ,  Ũ���-  Ũ����  �>����  �>���-  Ũ���-      D  , ,  ����  ����C  �����C  �����  ����      D  , ,  �d���  �d���C  �����C  �����  �d���      D  , ,  Ũ���  Ũ���C  �>���C  �>���  Ũ���      D  , ,  Ũ���m  Ũ���  �>���  �>���m  Ũ���m      D  , ,  ����m  ����  �����  �����m  ����m      D  , ,  �d���m  �d���  �����  �����m  �d���m      D  , ,  �����  �����C  �����C  �����  �����      D  , ,  �8���  �8���C  �����C  �����  �8���      D  , ,  �����  �����C  �&���C  �&���  �����      D  , ,  �����  �����C  �j���C  �j���  �����      D  , ,  �,���  �,���C  �����C  �����  �,���      D  , ,  �����m  �����  �����  �����m  �����m      D  , ,  �8���m  �8���  �����  �����m  �8���m      D  , ,  �����m  �����  �&���  �&���m  �����m      D  , ,  �����m  �����  �j���  �j���m  �����m      D  , ,  �,���m  �,���  �����  �����m  �,���m      D  , ,  �p���m  �p���  ����  ����m  �p���m      D  , ,  �����m  �����  �^���  �^���m  �����m      D  , ,  ̜���m  ̜���  �2���  �2���m  ̜���m      D  , ,  �����m  �����  �v���  �v���m  �����m      D  , ,  �8���m  �8���  �����  �����m  �8���m      D  , ,  �D���  �D���C  �����C  �����  �D���      D  , ,  ̜���  ̜���C  �2���C  �2���  ̜���      D  , ,  �'���  �'���  ɽ���  ɽ���  �'���      D  , ,  �D���  �D��ݯ  ����ݯ  �����  �D���      D  , ,  ̜���  ̜��ݯ  �2��ݯ  �2���  ̜���      D  , ,  �����  ����ݯ  �v��ݯ  �v���  �����      D  , ,  �8���  �8��ݯ  ����ݯ  �����  �8���      D  , ,  �u���  �u���  ����  ����  �u���      D  , ,  �'���C  �'����  ɽ����  ɽ���C  �'���C      D  , ,  �u���C  �u����  �����  ����C  �u���C      D  , ,  �����C  ������  �Y����  �Y���C  �����C      D  , ,  ����C  �����  Ч����  Ч���C  ����C      D  , ,  �����  �����  �Y���  �Y���  �����      D  , ,  �D���-  �D����  ������  �����-  �D���-      D  , ,  ̜���-  ̜����  �2����  �2���-  ̜���-      D  , ,  �D����  �D���  �����  ������  �D����      D  , ,  ̜����  ̜���  �2���  �2����  ̜����      D  , ,  ������  �����  �v���  �v����  ������      D  , ,  �8����  �8���  �����  ������  �8����      D  , ,  �����-  ������  �v����  �v���-  �����-      D  , ,  �8���-  �8����  ������  �����-  �8���-      D  , ,  �D���  �D���C  �����C  �����  �D���      D  , ,  ̜���  ̜���C  �2���C  �2���  ̜���      D  , ,  �����  �����C  �v���C  �v���  �����      D  , ,  �8���  �8���C  �����C  �����  �8���      D  , ,  ����  ����  Ч���  Ч���  ����      D  , ,  �����  �����C  �v���C  �v���  �����      D  , ,  �8���  �8���C  �����C  �����  �8���      D  , ,  �D���m  �D���  �����  �����m  �D���m      D  , ,  � ���c  � ����  Ȗ����  Ȗ���c  � ���c      D  , ,  � ��·  � ���  Ȗ���  Ȗ��·  � ��·      D  , ,  � ��ڙ  � ���/  Ȗ���/  Ȗ��ڙ  � ��ڙ      D  , ,  � ����  � ���o  Ȗ���o  Ȗ����  � ����      D  , ,  � ���#  � ��Ĺ  Ȗ��Ĺ  Ȗ���#  � ���#      D  , ,  � ���  � ��د  Ȗ��د  Ȗ���  � ���      D  , ,  � ���G  � ����  Ȗ����  Ȗ���G  � ���G      D  , ,  � ����  � ���]  Ȗ���]  Ȗ����  � ����      D  , ,  � ���  � ��̝  Ȗ��̝  Ȗ���  � ���      D  , ,  � ����  � ���y  Ȗ���y  Ȗ����  � ����      D  , ,  � ����  � ���o  Ȗ���o  Ȗ����  � ����      D  , ,  � ���Y  � ����  Ȗ����  Ȗ���Y  � ���Y      D  , ,  � ���Y  � ����  Ȗ����  Ȗ���Y  � ���Y      D  , ,  � ����  � ���9  Ȗ���9  Ȗ����  � ����      D  , ,  � ��ՙ  � ���/  Ȗ���/  Ȗ��ՙ  � ��ՙ      D  , ,  � ���c  � ����  Ȗ����  Ȗ���c  � ���c      D  , ,  �����  ����د  �v��د  �v���  �����      D  , ,  �8���  �8��د  ����د  �����  �8���      D  , ,  ̜��ڙ  ̜���/  �2���/  �2��ڙ  ̜��ڙ      D  , ,  ������  �����o  �v���o  �v����  ������      D  , ,  �8����  �8���o  �����o  ������  �8����      D  , ,  ����ڙ  �����/  �v���/  �v��ڙ  ����ڙ      D  , ,  ̜����  ̜���]  �2���]  �2����  ̜����      D  , ,  �8����  �8���]  �����]  ������  �8����      D  , ,  �8��ڙ  �8���/  �����/  ����ڙ  �8��ڙ      D  , ,  �8��·  �8���  �����  ����·  �8��·      D  , ,  �D����  �D���o  �����o  ������  �D����      D  , ,  �D����  �D���o  �����o  ������  �D����      D  , ,  ̜����  ̜���o  �2���o  �2����  ̜����      D  , ,  ������  �����o  �v���o  �v����  ������      D  , ,  �8����  �8���o  �����o  ������  �8����      D  , ,  ̜����  ̜���o  �2���o  �2����  ̜����      D  , ,  �D���Y  �D����  ������  �����Y  �D���Y      D  , ,  ̜���Y  ̜����  �2����  �2���Y  ̜���Y      D  , ,  �����Y  ������  �v����  �v���Y  �����Y      D  , ,  �8���Y  �8����  ������  �����Y  �8���Y      D  , ,  ̜��·  ̜���  �2���  �2��·  ̜��·      D  , ,  �D��ڙ  �D���/  �����/  ����ڙ  �D��ڙ      D  , ,  �D���Y  �D����  ������  �����Y  �D���Y      D  , ,  ̜���Y  ̜����  �2����  �2���Y  ̜���Y      D  , ,  �����Y  ������  �v����  �v���Y  �����Y      D  , ,  �8���Y  �8����  ������  �����Y  �8���Y      D  , ,  �D���  �D��د  ����د  �����  �D���      D  , ,  �D��ՙ  �D���/  �����/  ����ՙ  �D��ՙ      D  , ,  ̜��ՙ  ̜���/  �2���/  �2��ՙ  ̜��ՙ      D  , ,  ����ՙ  �����/  �v���/  �v��ՙ  ����ՙ      D  , ,  �8��ՙ  �8���/  �����/  ����ՙ  �8��ՙ      D  , ,  ̜���  ̜��د  �2��د  �2���  ̜���      D  , ,  �����Y  ������  �&����  �&���Y  �����Y      D  , ,  ������  �����]  �����]  ������  ������      D  , ,  ������  �����]  �&���]  �&����  ������      D  , ,  �,����  �,���]  �����]  ������  �,����      D  , ,  ������  �����]  �^���]  �^����  ������      D  , ,  �d����  �d���]  �����]  ������  �d����      D  , ,  Ũ��ڙ  Ũ���/  �>���/  �>��ڙ  Ũ��ڙ      D  , ,  �d��·  �d���  �����  ����·  �d��·      D  , ,  �����  ����د  ����د  �����  �����      D  , ,  �����Y  ������  �j����  �j���Y  �����Y      D  , ,  �8���  �8��د  ����د  �����  �8���      D  , ,  �,���Y  �,����  ������  �����Y  �,���Y      D  , ,  �����  ����د  �&��د  �&���  �����      D  , ,  �p���Y  �p����  �����  ����Y  �p���Y      D  , ,  �����Y  ������  �^����  �^���Y  �����Y      D  , ,  ����Y  �����  ������  �����Y  ����Y      D  , ,  �d���Y  �d����  ������  �����Y  �d���Y      D  , ,  Ũ���Y  Ũ����  �>����  �>���Y  Ũ���Y      D  , ,  ������  �����o  �����o  ������  ������      D  , ,  �8����  �8���o  �����o  ������  �8����      D  , ,  ������  �����o  �&���o  �&����  ������      D  , ,  ������  �����o  �j���o  �j����  ������      D  , ,  �,����  �,���o  �����o  ������  �,����      D  , ,  �p����  �p���o  ����o  �����  �p����      D  , ,  ������  �����o  �^���o  �^����  ������      D  , ,  �����  ����o  �����o  ������  �����      D  , ,  �d����  �d���o  �����o  ������  �d����      D  , ,  Ũ����  Ũ���o  �>���o  �>����  Ũ����      D  , ,  �����  ����د  �j��د  �j���  �����      D  , ,  �,���  �,��د  ����د  �����  �,���      D  , ,  �p���  �p��د  ���د  ����  �p���      D  , ,  �����  ����د  �^��د  �^���  �����      D  , ,  ����  ���د  ����د  �����  ����      D  , ,  �d���  �d��د  ����د  �����  �d���      D  , ,  Ũ���  Ũ��د  �>��د  �>���  Ũ���      D  , ,  �,��ڙ  �,���/  �����/  ����ڙ  �,��ڙ      D  , ,  �p��ڙ  �p���/  ����/  ���ڙ  �p��ڙ      D  , ,  ����ڙ  �����/  �^���/  �^��ڙ  ����ڙ      D  , ,  �����Y  ������  ������  �����Y  �����Y      D  , ,  �8���Y  �8����  ������  �����Y  �8���Y      D  , ,  �����Y  ������  �&����  �&���Y  �����Y      D  , ,  �����Y  ������  �j����  �j���Y  �����Y      D  , ,  �,���Y  �,����  ������  �����Y  �,���Y      D  , ,  �p���Y  �p����  �����  ����Y  �p���Y      D  , ,  �����Y  ������  �^����  �^���Y  �����Y      D  , ,  ����Y  �����  ������  �����Y  ����Y      D  , ,  �d���Y  �d����  ������  �����Y  �d���Y      D  , ,  Ũ���Y  Ũ����  �>����  �>���Y  Ũ���Y      D  , ,  ���ڙ  ����/  �����/  ����ڙ  ���ڙ      D  , ,  ������  �����o  �^���o  �^����  ������      D  , ,  �����  ����o  �����o  ������  �����      D  , ,  �d����  �d���o  �����o  ������  �d����      D  , ,  Ũ����  Ũ���o  �>���o  �>����  Ũ����      D  , ,  �d��ڙ  �d���/  �����/  ����ڙ  �d��ڙ      D  , ,  �,����  �,���o  �����o  ������  �,����      D  , ,  �p����  �p���o  ����o  �����  �p����      D  , ,  ����ڙ  �����/  �����/  ����ڙ  ����ڙ      D  , ,  �8��ڙ  �8���/  �����/  ����ڙ  �8��ڙ      D  , ,  ����ڙ  �����/  �&���/  �&��ڙ  ����ڙ      D  , ,  ����ڙ  �����/  �j���/  �j��ڙ  ����ڙ      D  , ,  ����·  �����  �����  ����·  ����·      D  , ,  ����·  �����  �&���  �&��·  ����·      D  , ,  �,��·  �,���  �����  ����·  �,��·      D  , ,  ����·  �����  �^���  �^��·  ����·      D  , ,  ����ՙ  �����/  �����/  ����ՙ  ����ՙ      D  , ,  �8��ՙ  �8���/  �����/  ����ՙ  �8��ՙ      D  , ,  ����ՙ  �����/  �&���/  �&��ՙ  ����ՙ      D  , ,  ����ՙ  �����/  �j���/  �j��ՙ  ����ՙ      D  , ,  �,��ՙ  �,���/  �����/  ����ՙ  �,��ՙ      D  , ,  �p��ՙ  �p���/  ����/  ���ՙ  �p��ՙ      D  , ,  ����ՙ  �����/  �^���/  �^��ՙ  ����ՙ      D  , ,  ���ՙ  ����/  �����/  ����ՙ  ���ՙ      D  , ,  �d��ՙ  �d���/  �����/  ����ՙ  �d��ՙ      D  , ,  Ũ��ՙ  Ũ���/  �>���/  �>��ՙ  Ũ��ՙ      D  , ,  ������  �����o  �����o  ������  ������      D  , ,  �8����  �8���o  �����o  ������  �8����      D  , ,  ������  �����o  �&���o  �&����  ������      D  , ,  ������  �����o  �j���o  �j����  ������      D  , ,  �����Y  ������  ������  �����Y  �����Y      D  , ,  �8���Y  �8����  ������  �����Y  �8���Y      D  , ,  ������  �����9  �����9  ������  ������      D  , ,  �L����  �L���9  �����9  ������  �L����      D  , ,  ������  �����9  �&���9  �&����  ������      D  , ,  ������  �����9  �~���9  �~����  ������      D  , ,  �,����  �,���9  �����9  ������  �,����      D  , ,  ������  �����9  ����9  �����  ������      D  , ,  ������  �����9  �^���9  �^����  ������      D  , ,  � ����  � ���9  �����9  ������  � ����      D  , ,  �d����  �d���9  �����9  ������  �d����      D  , ,  ż����  ż���9  �R���9  �R����  ż����      D  , ,  �����G  ������  �&����  �&���G  �����G      D  , ,  �,���G  �,����  ������  �����G  �,���G      D  , ,  �����G  ������  �^����  �^���G  �����G      D  , ,  �����#  ����Ĺ  ����Ĺ  �����#  �����#      D  , ,  �d���G  �d����  ������  �����G  �d���G      D  , ,  �L���#  �L��Ĺ  ����Ĺ  �����#  �L���#      D  , ,  �����#  ����Ĺ  �&��Ĺ  �&���#  �����#      D  , ,  �����#  ����Ĺ  �~��Ĺ  �~���#  �����#      D  , ,  �����  ����̝  ����̝  �����  �����      D  , ,  �����  ����̝  �&��̝  �&���  �����      D  , ,  �,���  �,��̝  ����̝  �����  �,���      D  , ,  �����  ����̝  �^��̝  �^���  �����      D  , ,  �d���  �d��̝  ����̝  �����  �d���      D  , ,  �,���#  �,��Ĺ  ����Ĺ  �����#  �,���#      D  , ,  �����#  ����Ĺ  ���Ĺ  ����#  �����#      D  , ,  �����c  ������  ������  �����c  �����c      D  , ,  �L���c  �L����  ������  �����c  �L���c      D  , ,  �����c  ������  �&����  �&���c  �����c      D  , ,  �����c  ������  �~����  �~���c  �����c      D  , ,  �,���c  �,����  ������  �����c  �,���c      D  , ,  �����c  ������  �����  ����c  �����c      D  , ,  ������  �����y  �����y  ������  ������      D  , ,  �L����  �L���y  �����y  ������  �L����      D  , ,  ������  �����y  �&���y  �&����  ������      D  , ,  ������  �����y  �~���y  �~����  ������      D  , ,  �,����  �,���y  �����y  ������  �,����      D  , ,  ������  �����y  ����y  �����  ������      D  , ,  ������  �����y  �^���y  �^����  ������      D  , ,  � ����  � ���y  �����y  ������  � ����      D  , ,  �d����  �d���y  �����y  ������  �d����      D  , ,  ż����  ż���y  �R���y  �R����  ż����      D  , ,  �����#  ����Ĺ  �^��Ĺ  �^���#  �����#      D  , ,  � ���#  � ��Ĺ  ����Ĺ  �����#  � ���#      D  , ,  �d���#  �d��Ĺ  ����Ĺ  �����#  �d���#      D  , ,  ż���#  ż��Ĺ  �R��Ĺ  �R���#  ż���#      D  , ,  ż���c  ż����  �R����  �R���c  ż���c      D  , ,  �����c  ������  �^����  �^���c  �����c      D  , ,  �����c  ������  ������  �����c  �����c      D  , ,  �L���c  �L����  ������  �����c  �L���c      D  , ,  �����c  ������  �&����  �&���c  �����c      D  , ,  �����c  ������  �~����  �~���c  �����c      D  , ,  �,���c  �,����  ������  �����c  �,���c      D  , ,  �����c  ������  �����  ����c  �����c      D  , ,  �����c  ������  �^����  �^���c  �����c      D  , ,  � ���c  � ����  ������  �����c  � ���c      D  , ,  �d���c  �d����  ������  �����c  �d���c      D  , ,  ż���c  ż����  �R����  �R���c  ż���c      D  , ,  �����G  ������  ������  �����G  �����G      D  , ,  � ���c  � ����  ������  �����c  � ���c      D  , ,  �d���c  �d����  ������  �����c  �d���c      D  , ,  �X���c  �X����  ������  �����c  �X���c      D  , ,  ̜���c  ̜����  �2����  �2���c  ̜���c      D  , ,  ̜���  ̜��̝  �2��̝  �2���  ̜���      D  , ,  �8���  �8��̝  ����̝  �����  �8���      D  , ,  �X����  �X���y  �����y  ������  �X����      D  , ,  ̜����  ̜���y  �2���y  �2����  ̜����      D  , ,  ������  �����y  ϊ���y  ϊ����  ������      D  , ,  �X����  �X���9  �����9  ������  �X����      D  , ,  ̜����  ̜���9  �2���9  �2����  ̜����      D  , ,  ������  �����9  ϊ���9  ϊ����  ������      D  , ,  �8����  �8���9  �����9  ������  �8����      D  , ,  �8����  �8���y  �����y  ������  �8����      D  , ,  �����c  ������  ϊ����  ϊ���c  �����c      D  , ,  �X���#  �X��Ĺ  ����Ĺ  �����#  �X���#      D  , ,  ̜���#  ̜��Ĺ  �2��Ĺ  �2���#  ̜���#      D  , ,  �����#  ����Ĺ  ϊ��Ĺ  ϊ���#  �����#      D  , ,  ̜���G  ̜����  �2����  �2���G  ̜���G      D  , ,  �8���G  �8����  ������  �����G  �8���G      D  , ,  �X���c  �X����  ������  �����c  �X���c      D  , ,  ̜���c  ̜����  �2����  �2���c  ̜���c      D  , ,  �����c  ������  ϊ����  ϊ���c  �����c      D  , ,  �8���c  �8����  ������  �����c  �8���c      D  , ,  �8���#  �8��Ĺ  ����Ĺ  �����#  �8���#      D  , ,  �8���c  �8����  ������  �����c  �8���c      D  , ,  �����#  ������  �F����  �F���#  �����#      D  , ,  ������  �����y  �F���y  �F����  ������      D  , ,  ������  �����9  �F���9  �F����  ������      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ������  �����e  �F���e  �F����  ������      D  , ,  ������  �����%  �F���%  �F����  ������      D  , ,  �����O  ������  �F����  �F���O  �����O      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ������  �����e  �F���e  �F����  ������      D  , ,  ������  �����%  �F���%  �F����  ������      D  , ,  �����O  ������  �F����  �F���O  �����O      D  , ,  �����Y  ������  �F����  �F���Y  �����Y      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ������  �����o  �F���o  �F����  ������      D  , ,  ������  �����/  �F���/  �F����  ������      D  , ,  �����Y  ������  �F����  �F���Y  �����Y      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ������  �����o  �F���o  �F����  ������      D  , ,  ������  �����/  �F���/  �F����  ������      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ������  �����[  �F���[  �F����  ������      D  , ,  ������  �����  �F���  �F����  ������      D  , ,  �����E  ������  �F����  �F���E  �����E      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ������  �����[  �F���[  �F����  ������      D  , ,  ������  �����  �F���  �F����  ������      D  , ,  �����E  ������  �F����  �F���E  �����E      D  , ,  ����q�  ����r   �(��r   �(��q�  ����q�      D  , ,  ����pJ  ����p�  �(��p�  �(��pJ  ����pJ      D  , ,  ����o
  ����o�  �(��o�  �(��o
  ����o
      D  , ,  ����m�  ����n`  �(��n`  �(��m�  ����m�      D  , ,  ����l�  ����m   �(��m   �(��l�  ����l�      D  , ,  ����kJ  ����k�  �(��k�  �(��kJ  ����kJ      D  , ,  ����j
  ����j�  �(��j�  �(��j
  ����j
      D  , ,  ����h�  ����i`  �(��i`  �(��h�  ����h�      D  , ,  ����a�  ����b&  �(��b&  �(��a�  ����a�      D  , ,  ����`P  ����`�  �(��`�  �(��`P  ����`P      D  , ,  ����_  ����_�  �(��_�  �(��_  ����_      D  , ,  ����]�  ����^f  �(��^f  �(��]�  ����]�      D  , ,  ����\�  ����]&  �(��]&  �(��\�  ����\�      D  , ,  ����[P  ����[�  �(��[�  �(��[P  ����[P      D  , ,  ����Z  ����Z�  �(��Z�  �(��Z  ����Z      D  , ,  ����X�  ����Yf  �(��Yf  �(��X�  ����X�      D  , ,  � ����  � ���9  Ȗ���9  Ȗ����  � ����      D  , ,  � ���  � ����  Ȗ����  Ȗ���  � ���      D  , ,  � ����  � ���e  Ȗ���e  Ȗ����  � ����      D  , ,  � ����  � ���%  Ȗ���%  Ȗ����  � ����      D  , ,  �����O  ������  ������  �����O  �����O      D  , ,  �L���O  �L����  ������  �����O  �L���O      D  , ,  �����O  ������  �&����  �&���O  �����O      D  , ,  �����O  ������  �~����  �~���O  �����O      D  , ,  �,���O  �,����  ������  �����O  �,���O      D  , ,  �����O  ������  �����  ����O  �����O      D  , ,  �����O  ������  �^����  �^���O  �����O      D  , ,  � ���O  � ����  ������  �����O  � ���O      D  , ,  �d���O  �d����  ������  �����O  �d���O      D  , ,  ż���O  ż����  �R����  �R���O  ż���O      D  , ,  � ���O  � ����  Ȗ����  Ȗ���O  � ���O      D  , ,  �X���O  �X����  ������  �����O  �X���O      D  , ,  ̜���O  ̜����  �2����  �2���O  ̜���O      D  , ,  �����O  ������  ϊ����  ϊ���O  �����O      D  , ,  �8���O  �8����  ������  �����O  �8���O      D  , ,  � ���  � ����  Ȗ����  Ȗ���  � ���      D  , ,  � ����  � ���e  Ȗ���e  Ȗ����  � ����      D  , ,  � ����  � ���%  Ȗ���%  Ȗ����  � ����      D  , ,  � ���O  � ����  Ȗ����  Ȗ���O  � ���O      D  , ,  � ����  � ���S  Ȗ���S  Ȗ����  � ����      D  , ,  � ���}  � ���  Ȗ���  Ȗ���}  � ���}      D  , ,  � ���=  � ����  Ȗ����  Ȗ���=  � ���=      D  , ,  � ����  � ����  Ȗ����  Ȗ����  � ����      D  , ,  � ���#  � ����  Ȗ����  Ȗ���#  � ���#      D  , ,  � ����  � ���y  Ȗ���y  Ȗ����  � ����      D  , ,  �'���y  �'���  ɽ���  ɽ���y  �'���y      D  , ,  �u���y  �u���  ����  ����y  �u���y      D  , ,  �����y  �����  �Y���  �Y���y  �����y      D  , ,  ����y  ����  Ч���  Ч���y  ����y      D  , ,  �'���9  �'����  ɽ����  ɽ���9  �'���9      D  , ,  �u���9  �u����  �����  ����9  �u���9      D  , ,  �����9  ������  �Y����  �Y���9  �����9      D  , ,  ����9  �����  Ч����  Ч���9  ����9      D  , ,  �X����  �X���9  �����9  ������  �X����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  ̜���  ̜����  �2����  �2���  ̜���      D  , ,  �����  ������  ϊ����  ϊ���  �����      D  , ,  �8���  �8����  ������  �����  �8���      D  , ,  ̜����  ̜���9  �2���9  �2����  ̜����      D  , ,  �X����  �X���e  �����e  ������  �X����      D  , ,  ̜����  ̜���e  �2���e  �2����  ̜����      D  , ,  ������  �����e  ϊ���e  ϊ����  ������      D  , ,  �8����  �8���e  �����e  ������  �8����      D  , ,  ������  �����9  ϊ���9  ϊ����  ������      D  , ,  �X����  �X���%  �����%  ������  �X����      D  , ,  ̜����  ̜���%  �2���%  �2����  ̜����      D  , ,  ������  �����%  ϊ���%  ϊ����  ������      D  , ,  �8����  �8���%  �����%  ������  �8����      D  , ,  �X���#  �X����  ������  �����#  �X���#      D  , ,  ̜���#  ̜����  �2����  �2���#  ̜���#      D  , ,  �����#  ������  ϊ����  ϊ���#  �����#      D  , ,  �8���#  �8����  ������  �����#  �8���#      D  , ,  �8����  �8���9  �����9  ������  �8����      D  , ,  �X����  �X���y  �����y  ������  �X����      D  , ,  ̜����  ̜���y  �2���y  �2����  ̜����      D  , ,  ������  �����y  ϊ���y  ϊ����  ������      D  , ,  �8����  �8���y  �����y  ������  �8����      D  , ,  ż����  ż���e  �R���e  �R����  ż����      D  , ,  �i���y  �i���  �����  �����y  �i���y      D  , ,  �����y  �����  �M���  �M���y  �����y      D  , ,  �����9  ������  �c����  �c���9  �����9      D  , ,  ����9  �����  ������  �����9  ����9      D  , ,  �i���9  �i����  ������  �����9  �i���9      D  , ,  �,���#  �,����  ������  �����#  �,���#      D  , ,  ������  �����%  �����%  ������  ������      D  , ,  �L����  �L���%  �����%  ������  �L����      D  , ,  ������  �����%  �&���%  �&����  ������      D  , ,  ������  �����%  �~���%  �~����  ������      D  , ,  �,����  �,���%  �����%  ������  �,����      D  , ,  ������  �����%  ����%  �����  ������      D  , ,  ������  �����%  �^���%  �^����  ������      D  , ,  � ����  � ���%  �����%  ������  � ����      D  , ,  �d����  �d���%  �����%  ������  �d����      D  , ,  ż����  ż���%  �R���%  �R����  ż����      D  , ,  �����9  ������  �M����  �M���9  �����9      D  , ,  ����9  �����  ������  �����9  ����9      D  , ,  �S���9  �S����  ������  �����9  �S���9      D  , ,  �����9  ������  �7����  �7���9  �����9      D  , ,  �����9  ������  ������  �����9  �����9      D  , ,  �����#  ������  �����  ����#  �����#      D  , ,  �=���9  �=����  ������  �����9  �=���9      D  , ,  ċ���9  ċ����  �!����  �!���9  ċ���9      D  , ,  �����9  ������  �o����  �o���9  �����9      D  , ,  ����y  ����  �����  �����y  ����y      D  , ,  �S���y  �S���  �����  �����y  �S���y      D  , ,  �����y  �����  �7���  �7���y  �����y      D  , ,  �����y  �����  �����  �����y  �����y      D  , ,  �����#  ������  �&����  �&���#  �����#      D  , ,  �����  ������  ������  �����  �����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  �����  ������  �&����  �&���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �,���  �,����  ������  �����  �,���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����  ������  �^����  �^���  �����      D  , ,  �����#  ������  �^����  �^���#  �����#      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  � ���#  � ����  ������  �����#  � ���#      D  , ,  �d���  �d����  ������  �����  �d���      D  , ,  �d���#  �d����  ������  �����#  �d���#      D  , ,  ż���  ż����  �R����  �R���  ż���      D  , ,  ż���#  ż����  �R����  �R���#  ż���#      D  , ,  �=���y  �=���  �����  �����y  �=���y      D  , ,  ċ���y  ċ���  �!���  �!���y  ċ���y      D  , ,  �����y  �����  �o���  �o���y  �����y      D  , ,  �����y  �����  �c���  �c���y  �����y      D  , ,  ����y  ����  �����  �����y  ����y      D  , ,  �����#  ������  �~����  �~���#  �����#      D  , ,  ������  �����e  �����e  ������  ������      D  , ,  �L����  �L���e  �����e  ������  �L����      D  , ,  ������  �����e  �&���e  �&����  ������      D  , ,  ������  �����e  �~���e  �~����  ������      D  , ,  �����#  ������  ������  �����#  �����#      D  , ,  ������  �����y  �����y  ������  ������      D  , ,  �L����  �L���y  �����y  ������  �L����      D  , ,  ������  �����y  �&���y  �&����  ������      D  , ,  ������  �����y  �~���y  �~����  ������      D  , ,  �,����  �,���y  �����y  ������  �,����      D  , ,  ������  �����y  ����y  �����  ������      D  , ,  ������  �����y  �^���y  �^����  ������      D  , ,  � ����  � ���y  �����y  ������  � ����      D  , ,  �d����  �d���y  �����y  ������  �d����      D  , ,  ż����  ż���y  �R���y  �R����  ż����      D  , ,  �,����  �,���e  �����e  ������  �,����      D  , ,  ������  �����e  ����e  �����  ������      D  , ,  ������  �����e  �^���e  �^����  ������      D  , ,  � ����  � ���e  �����e  ������  � ����      D  , ,  �d����  �d���e  �����e  ������  �d����      D  , ,  �L���#  �L����  ������  �����#  �L���#      D  , ,  ������  �����9  �����9  ������  ������      D  , ,  �L����  �L���9  �����9  ������  �L����      D  , ,  ������  �����9  �&���9  �&����  ������      D  , ,  ������  �����9  �~���9  �~����  ������      D  , ,  �,����  �,���9  �����9  ������  �,����      D  , ,  ������  �����9  ����9  �����  ������      D  , ,  ������  �����9  �^���9  �^����  ������      D  , ,  � ����  � ���9  �����9  ������  � ����      D  , ,  �d����  �d���9  �����9  ������  �d����      D  , ,  ż����  ż���9  �R���9  �R����  ż����      D  , ,  � ���O  � ����  ������  �����O  � ���O      D  , ,  �d���O  �d����  ������  �����O  �d���O      D  , ,  ż���O  ż����  �R����  �R���O  ż���O      D  , ,  �����  ������  �^����  �^���  �����      D  , ,  ������  �����S  �����S  ������  ������      D  , ,  ������  �����S  �&���S  �&����  ������      D  , ,  �,����  �,���S  �����S  ������  �,����      D  , ,  ������  �����S  �^���S  �^����  ������      D  , ,  �d����  �d���S  �����S  ������  �d����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �����}  �����  �����  �����}  �����}      D  , ,  �����}  �����  �&���  �&���}  �����}      D  , ,  �,���}  �,���  �����  �����}  �,���}      D  , ,  �����}  �����  �^���  �^���}  �����}      D  , ,  �d���}  �d���  �����  �����}  �d���}      D  , ,  �d���  �d����  ������  �����  �d���      D  , ,  �����=  ������  ������  �����=  �����=      D  , ,  �����=  ������  �&����  �&���=  �����=      D  , ,  �,���=  �,����  ������  �����=  �,���=      D  , ,  �����=  ������  �^����  �^���=  �����=      D  , ,  �d���=  �d����  ������  �����=  �d���=      D  , ,  ż���  ż����  �R����  �R���  ż���      D  , ,  ������  ������  ������  ������  ������      D  , ,  ������  ������  �&����  �&����  ������      D  , ,  �,����  �,����  ������  ������  �,����      D  , ,  ������  ������  �^����  �^����  ������      D  , ,  �d����  �d����  ������  ������  �d����      D  , ,  �����  ������  ������  �����  �����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  ������  �����e  �����e  ������  ������      D  , ,  �L����  �L���e  �����e  ������  �L����      D  , ,  ������  �����e  �&���e  �&����  ������      D  , ,  ������  �����e  �~���e  �~����  ������      D  , ,  �,����  �,���e  �����e  ������  �,����      D  , ,  ������  �����e  ����e  �����  ������      D  , ,  ������  �����e  �^���e  �^����  ������      D  , ,  � ����  � ���e  �����e  ������  � ����      D  , ,  �d����  �d���e  �����e  ������  �d����      D  , ,  ż����  ż���e  �R���e  �R����  ż����      D  , ,  �����  ������  �&����  �&���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  ������  �����%  �����%  ������  ������      D  , ,  �L����  �L���%  �����%  ������  �L����      D  , ,  ������  �����%  �&���%  �&����  ������      D  , ,  ������  �����%  �~���%  �~����  ������      D  , ,  �,����  �,���%  �����%  ������  �,����      D  , ,  ������  �����%  ����%  �����  ������      D  , ,  ������  �����%  �^���%  �^����  ������      D  , ,  � ����  � ���%  �����%  ������  � ����      D  , ,  �d����  �d���%  �����%  ������  �d����      D  , ,  ż����  ż���%  �R���%  �R����  ż����      D  , ,  �,���  �,����  ������  �����  �,���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����O  ������  ������  �����O  �����O      D  , ,  �L���O  �L����  ������  �����O  �L���O      D  , ,  �����O  ������  �&����  �&���O  �����O      D  , ,  �����O  ������  �~����  �~���O  �����O      D  , ,  �,���O  �,����  ������  �����O  �,���O      D  , ,  �����O  ������  �����  ����O  �����O      D  , ,  �����O  ������  �^����  �^���O  �����O      D  , ,  �X���O  �X����  ������  �����O  �X���O      D  , ,  ̜���O  ̜����  �2����  �2���O  ̜���O      D  , ,  �����O  ������  ϊ����  ϊ���O  �����O      D  , ,  �8���O  �8����  ������  �����O  �8���O      D  , ,  �X����  �X���e  �����e  ������  �X����      D  , ,  ̜����  ̜���e  �2���e  �2����  ̜����      D  , ,  ̜���=  ̜����  �2����  �2���=  ̜���=      D  , ,  �8���=  �8����  ������  �����=  �8���=      D  , ,  ������  �����e  ϊ���e  ϊ����  ������      D  , ,  �8����  �8���e  �����e  ������  �8����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  ̜���  ̜����  �2����  �2���  ̜���      D  , ,  ̜����  ̜���S  �2���S  �2����  ̜����      D  , ,  �8����  �8���S  �����S  ������  �8����      D  , ,  ̜����  ̜����  �2����  �2����  ̜����      D  , ,  �8����  �8����  ������  ������  �8����      D  , ,  �����  ������  ϊ����  ϊ���  �����      D  , ,  �8���  �8����  ������  �����  �8���      D  , ,  �X����  �X���%  �����%  ������  �X����      D  , ,  ̜����  ̜���%  �2���%  �2����  ̜����      D  , ,  ������  �����%  ϊ���%  ϊ����  ������      D  , ,  �8����  �8���%  �����%  ������  �8����      D  , ,  ̜���}  ̜���  �2���  �2���}  ̜���}      D  , ,  �8���}  �8���  �����  �����}  �8���}      D  , ,  � ����  � ���o  Ȗ���o  Ȗ����  � ����      D  , ,  � ����  � ���/  Ȗ���/  Ȗ����  � ����      D  , ,  � ���Y  � ����  Ȗ����  Ȗ���Y  � ���Y      D  , ,  � ���  � ����  Ȗ����  Ȗ���  � ���      D  , ,  � ����  � ���o  Ȗ���o  Ȗ����  � ����      D  , ,  ������  �����/  �����/  ������  ������      D  , ,  �L����  �L���/  �����/  ������  �L����      D  , ,  ������  �����/  �&���/  �&����  ������      D  , ,  ������  �����/  �~���/  �~����  ������      D  , ,  �,����  �,���/  �����/  ������  �,����      D  , ,  ������  �����/  ����/  �����  ������      D  , ,  ������  �����/  �^���/  �^����  ������      D  , ,  � ����  � ���/  �����/  ������  � ����      D  , ,  �d����  �d���/  �����/  ������  �d����      D  , ,  ż����  ż���/  �R���/  �R����  ż����      D  , ,  � ����  � ���/  Ȗ���/  Ȗ����  � ����      D  , ,  �X����  �X���/  �����/  ������  �X����      D  , ,  ̜����  ̜���/  �2���/  �2����  ̜����      D  , ,  ������  �����/  ϊ���/  ϊ����  ������      D  , ,  �8����  �8���/  �����/  ������  �8����      D  , ,  � ���  � ����  Ȗ����  Ȗ���  � ���      D  , ,  � ����  � ���[  Ȗ���[  Ȗ����  � ����      D  , ,  � ����  � ���  Ȗ���  Ȗ����  � ����      D  , ,  � ���Y  � ����  Ȗ����  Ȗ���Y  � ���Y      D  , ,  � ���E  � ����  Ȗ����  Ȗ���E  � ���E      D  , ,  � ���  � ����  Ȗ����  Ȗ���  � ���      D  , ,  � ����  � ���[  Ȗ���[  Ȗ����  � ����      D  , ,  � ���  � ����  Ȗ����  Ȗ���  � ���      D  , ,  ������  �����/  ϊ���/  ϊ����  ������      D  , ,  �8����  �8���/  �����/  ������  �8����      D  , ,  ̜����  ̜���o  �2���o  �2����  ̜����      D  , ,  �X���Y  �X����  ������  �����Y  �X���Y      D  , ,  ̜���Y  ̜����  �2����  �2���Y  ̜���Y      D  , ,  �����Y  ������  ϊ����  ϊ���Y  �����Y      D  , ,  �8���Y  �8����  ������  �����Y  �8���Y      D  , ,  ������  �����o  ϊ���o  ϊ����  ������      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  ̜���  ̜����  �2����  �2���  ̜���      D  , ,  �����  ������  ϊ����  ϊ���  �����      D  , ,  �8���  �8����  ������  �����  �8���      D  , ,  �8����  �8���o  �����o  ������  �8����      D  , ,  �X����  �X���o  �����o  ������  �X����      D  , ,  ̜����  ̜���o  �2���o  �2����  ̜����      D  , ,  ������  �����o  ϊ���o  ϊ����  ������      D  , ,  �8����  �8���o  �����o  ������  �8����      D  , ,  �X���Y  �X����  ������  �����Y  �X���Y      D  , ,  �X����  �X���o  �����o  ������  �X����      D  , ,  ̜���Y  ̜����  �2����  �2���Y  ̜���Y      D  , ,  �X����  �X���/  �����/  ������  �X����      D  , ,  �����Y  ������  ϊ����  ϊ���Y  �����Y      D  , ,  �8���Y  �8����  ������  �����Y  �8���Y      D  , ,  ̜����  ̜���/  �2���/  �2����  ̜����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  ̜���  ̜����  �2����  �2���  ̜���      D  , ,  �����  ������  ϊ����  ϊ���  �����      D  , ,  �8���  �8����  ������  �����  �8���      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �d���  �d����  ������  �����  �d���      D  , ,  ż���  ż����  �R����  �R���  ż���      D  , ,  ������  �����o  �~���o  �~����  ������      D  , ,  �����Y  ������  �&����  �&���Y  �����Y      D  , ,  ������  �����/  �����/  ������  ������      D  , ,  �L����  �L���/  �����/  ������  �L����      D  , ,  ������  �����/  �&���/  �&����  ������      D  , ,  �����Y  ������  �����  ����Y  �����Y      D  , ,  ������  �����o  �����o  ������  ������      D  , ,  �L����  �L���o  �����o  ������  �L����      D  , ,  ������  �����o  �&���o  �&����  ������      D  , ,  ������  �����o  �~���o  �~����  ������      D  , ,  �,����  �,���o  �����o  ������  �,����      D  , ,  ������  �����o  ����o  �����  ������      D  , ,  ������  �����o  �^���o  �^����  ������      D  , ,  � ����  � ���o  �����o  ������  � ����      D  , ,  �d����  �d���o  �����o  ������  �d����      D  , ,  ż����  ż���o  �R���o  �R����  ż����      D  , ,  ������  �����/  �~���/  �~����  ������      D  , ,  �,����  �,���/  �����/  ������  �,����      D  , ,  ������  �����/  ����/  �����  ������      D  , ,  ������  �����/  �^���/  �^����  ������      D  , ,  � ����  � ���/  �����/  ������  � ����      D  , ,  �����Y  ������  �^����  �^���Y  �����Y      D  , ,  �d����  �d���/  �����/  ������  �d����      D  , ,  ż����  ż���/  �R���/  �R����  ż����      D  , ,  �,����  �,���o  �����o  ������  �,����      D  , ,  ������  �����o  ����o  �����  ������      D  , ,  ������  �����o  �^���o  �^����  ������      D  , ,  � ����  � ���o  �����o  ������  � ����      D  , ,  �d����  �d���o  �����o  ������  �d����      D  , ,  �����Y  ������  �~����  �~���Y  �����Y      D  , ,  �����Y  ������  ������  �����Y  �����Y      D  , ,  �L���Y  �L����  ������  �����Y  �L���Y      D  , ,  �����Y  ������  �&����  �&���Y  �����Y      D  , ,  �����Y  ������  �~����  �~���Y  �����Y      D  , ,  �,���Y  �,����  ������  �����Y  �,���Y      D  , ,  �����Y  ������  �����  ����Y  �����Y      D  , ,  �����Y  ������  �^����  �^���Y  �����Y      D  , ,  � ���Y  � ����  ������  �����Y  � ���Y      D  , ,  � ���Y  � ����  ������  �����Y  � ���Y      D  , ,  �d���Y  �d����  ������  �����Y  �d���Y      D  , ,  �d���Y  �d����  ������  �����Y  �d���Y      D  , ,  ż���Y  ż����  �R����  �R���Y  ż���Y      D  , ,  ż���Y  ż����  �R����  �R���Y  ż���Y      D  , ,  ż����  ż���o  �R���o  �R����  ż����      D  , ,  �L���Y  �L����  ������  �����Y  �L���Y      D  , ,  ������  �����o  �����o  ������  ������      D  , ,  �L����  �L���o  �����o  ������  �L����      D  , ,  ������  �����o  �&���o  �&����  ������      D  , ,  �,���Y  �,����  ������  �����Y  �,���Y      D  , ,  �����  ������  ������  �����  �����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  �����Y  ������  ������  �����Y  �����Y      D  , ,  �����  ������  ������  �����  �����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  �����  ������  �&����  �&���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �,���  �,����  ������  �����  �,���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����  ������  �^����  �^���  �����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �d���  �d����  ������  �����  �d���      D  , ,  ż���  ż����  �R����  �R���  ż���      D  , ,  �����  ������  �&����  �&���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �,���  �,����  ������  �����  �,���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����  ������  �^����  �^���  �����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �d���  �d����  ������  �����  �d���      D  , ,  ż���  ż����  �R����  �R���  ż���      D  , ,  ����o  ����  �����  �����o  ����o      D  , ,  �i���o  �i���  �����  �����o  �i���o      D  , ,  ������  �����[  �����[  ������  ������      D  , ,  �L����  �L���[  �����[  ������  �L����      D  , ,  ������  �����[  �&���[  �&����  ������      D  , ,  ������  �����[  �~���[  �~����  ������      D  , ,  �,����  �,���[  �����[  ������  �,����      D  , ,  ������  �����[  ����[  �����  ������      D  , ,  ������  �����[  �^���[  �^����  ������      D  , ,  � ����  � ���[  �����[  ������  � ����      D  , ,  �d����  �d���[  �����[  ������  �d����      D  , ,  ż����  ż���[  �R���[  �R����  ż����      D  , ,  �����o  �����  �M���  �M���o  �����o      D  , ,  ����o  ����  �����  �����o  ����o      D  , ,  ������  �����  �����  ������  ������      D  , ,  �L����  �L���  �����  ������  �L����      D  , ,  ������  �����  �&���  �&����  ������      D  , ,  ������  �����  �~���  �~����  ������      D  , ,  �,����  �,���  �����  ������  �,����      D  , ,  ������  �����  ����  �����  ������      D  , ,  ������  �����  �^���  �^����  ������      D  , ,  � ����  � ���  �����  ������  � ����      D  , ,  �d����  �d���  �����  ������  �d����      D  , ,  ż����  ż���  �R���  �R����  ż����      D  , ,  �S���o  �S���  �����  �����o  �S���o      D  , ,  �����o  �����  �7���  �7���o  �����o      D  , ,  �����E  ������  ������  �����E  �����E      D  , ,  �L���E  �L����  ������  �����E  �L���E      D  , ,  �����E  ������  �&����  �&���E  �����E      D  , ,  �����E  ������  �~����  �~���E  �����E      D  , ,  �,���E  �,����  ������  �����E  �,���E      D  , ,  �����E  ������  �����  ����E  �����E      D  , ,  �����E  ������  �^����  �^���E  �����E      D  , ,  � ���E  � ����  ������  �����E  � ���E      D  , ,  �d���E  �d����  ������  �����E  �d���E      D  , ,  ż���E  ż����  �R����  �R���E  ż���E      D  , ,  �����o  �����  �����  �����o  �����o      D  , ,  �=���o  �=���  �����  �����o  �=���o      D  , ,  �����  ������  ������  �����  �����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  �����  ������  �&����  �&���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �,���  �,����  ������  �����  �,���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����  ������  �^����  �^���  �����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �d���  �d����  ������  �����  �d���      D  , ,  ż���  ż����  �R����  �R���  ż���      D  , ,  ċ���o  ċ���  �!���  �!���o  ċ���o      D  , ,  �����o  �����  �o���  �o���o  �����o      D  , ,  ������  �����[  �����[  ������  ������      D  , ,  �L����  �L���[  �����[  ������  �L����      D  , ,  ������  �����[  �&���[  �&����  ������      D  , ,  ������  �����[  �~���[  �~����  ������      D  , ,  �,����  �,���[  �����[  ������  �,����      D  , ,  ������  �����[  ����[  �����  ������      D  , ,  ������  �����[  �^���[  �^����  ������      D  , ,  � ����  � ���[  �����[  ������  � ����      D  , ,  �d����  �d���[  �����[  ������  �d����      D  , ,  ż����  ż���[  �R���[  �R����  ż����      D  , ,  �����/  ������  �c����  �c���/  �����/      D  , ,  ����/  �����  ������  �����/  ����/      D  , ,  �i���/  �i����  ������  �����/  �i���/      D  , ,  �����/  ������  �M����  �M���/  �����/      D  , ,  ����/  �����  ������  �����/  ����/      D  , ,  �S���/  �S����  ������  �����/  �S���/      D  , ,  �����/  ������  �7����  �7���/  �����/      D  , ,  �����/  ������  ������  �����/  �����/      D  , ,  �=���/  �=����  ������  �����/  �=���/      D  , ,  ċ���/  ċ����  �!����  �!���/  ċ���/      D  , ,  �����/  ������  �o����  �o���/  �����/      D  , ,  �����o  �����  �c���  �c���o  �����o      D  , ,  �����  ������  ������  �����  �����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  �����  ������  �&����  �&���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �,���  �,����  ������  �����  �,���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����  ������  �^����  �^���  �����      D  , ,  �����/  ������  �Y����  �Y���/  �����/      D  , ,  ����/  �����  Ч����  Ч���/  ����/      D  , ,  ����o  ����  Ч���  Ч���o  ����o      D  , ,  �'���o  �'���  ɽ���  ɽ���o  �'���o      D  , ,  �u���o  �u���  ����  ����o  �u���o      D  , ,  �����o  �����  �Y���  �Y���o  �����o      D  , ,  �X���E  �X����  ������  �����E  �X���E      D  , ,  ̜���E  ̜����  �2����  �2���E  ̜���E      D  , ,  �����E  ������  ϊ����  ϊ���E  �����E      D  , ,  �8���E  �8����  ������  �����E  �8���E      D  , ,  �X����  �X���[  �����[  ������  �X����      D  , ,  ̜����  ̜���[  �2���[  �2����  ̜����      D  , ,  ������  �����[  ϊ���[  ϊ����  ������      D  , ,  �8����  �8���[  �����[  ������  �8����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  ̜���  ̜����  �2����  �2���  ̜���      D  , ,  �����  ������  ϊ����  ϊ���  �����      D  , ,  �8���  �8����  ������  �����  �8���      D  , ,  �X����  �X���  �����  ������  �X����      D  , ,  ̜����  ̜���  �2���  �2����  ̜����      D  , ,  ������  �����  ϊ���  ϊ����  ������      D  , ,  �8����  �8���  �����  ������  �8����      D  , ,  �X����  �X���[  �����[  ������  �X����      D  , ,  ̜����  ̜���[  �2���[  �2����  ̜����      D  , ,  ������  �����[  ϊ���[  ϊ����  ������      D  , ,  �8����  �8���[  �����[  ������  �8����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  ̜���  ̜����  �2����  �2���  ̜���      D  , ,  �����  ������  ϊ����  ϊ���  �����      D  , ,  �8���  �8����  ������  �����  �8���      D  , ,  �'���/  �'����  ɽ����  ɽ���/  �'���/      D  , ,  �u���/  �u����  �����  ����/  �u���/      D  , ,  ~@���O  ~@����  ~�����  ~����O  ~@���O      D  , ,  �����O  ������  �.����  �.���O  �����O      D  , ,  �����O  ������  �r����  �r���O  �����O      D  , ,  �4���O  �4����  ������  �����O  �4���O      D  , ,  �x���O  �x����  �����  ����O  �x���O      D  , ,  �����O  ������  �f����  �f���O  �����O      D  , ,  ����O  �����  ������  �����O  ����O      D  , ,  �l���O  �l����  �����  ����O  �l���O      D  , ,  �����O  ������  �F����  �F���O  �����O      D  , ,  ����O  �����  ������  �����O  ����O      D  , ,  �L���O  �L����  ������  �����O  �L���O      D  , ,  �����O  ������  �:����  �:���O  �����O      D  , ,  �����O  ������  �~����  �~���O  �����O      D  , ,  �@���O  �@����  ������  �����O  �@���O      D  , ,  �����O  ������  �����  ����O  �����O      D  , ,  �����O  ������  �r����  �r���O  �����O      D  , ,  � ���O  � ����  ������  �����O  � ���O      D  , ,  �x���O  �x����  �����  ����O  �x���O      D  , ,  �����O  ������  �R����  �R���O  �����O      D  , ,  ����O  �����  ������  �����O  ����O      D  , ,  �X���O  �X����  ������  �����O  �X���O      D  , ,  ����9  �����  �����  ����9  ����9      D  , ,  ������  �����y  �:���y  �:����  ������      D  , ,  ������  �����y  �~���y  �~����  ������      D  , ,  �@����  �@���y  �����y  ������  �@����      D  , ,  ������  �����y  ����y  �����  ������      D  , ,  �����  ������  �:����  �:���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �@���  �@����  ������  �����  �@���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �R����  �R���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  ������  �����y  �r���y  �r����  ������      D  , ,  � ����  � ���y  �����y  ������  � ����      D  , ,  �x����  �x���y  ����y  �����  �x����      D  , ,  ������  �����y  �R���y  �R����  ������      D  , ,  �����  ����y  �����y  ������  �����      D  , ,  �X����  �X���y  �����y  ������  �X����      D  , ,  �����#  ������  �:����  �:���#  �����#      D  , ,  �����#  ������  �~����  �~���#  �����#      D  , ,  �@���#  �@����  ������  �����#  �@���#      D  , ,  ������  �����e  �:���e  �:����  ������      D  , ,  ������  �����e  �~���e  �~����  ������      D  , ,  �@����  �@���e  �����e  ������  �@����      D  , ,  ������  �����e  ����e  �����  ������      D  , ,  ������  �����e  �r���e  �r����  ������      D  , ,  � ����  � ���e  �����e  ������  � ����      D  , ,  �x����  �x���e  ����e  �����  �x����      D  , ,  ������  �����e  �R���e  �R����  ������      D  , ,  �����  ����e  �����e  ������  �����      D  , ,  �X����  �X���e  �����e  ������  �X����      D  , ,  �����#  ������  �����  ����#  �����#      D  , ,  �����#  ������  �r����  �r���#  �����#      D  , ,  � ���#  � ����  ������  �����#  � ���#      D  , ,  �x���#  �x����  �����  ����#  �x���#      D  , ,  �����#  ������  �R����  �R���#  �����#      D  , ,  ����#  �����  ������  �����#  ����#      D  , ,  ������  �����%  �:���%  �:����  ������      D  , ,  ������  �����%  �~���%  �~����  ������      D  , ,  �@����  �@���%  �����%  ������  �@����      D  , ,  ������  �����%  ����%  �����  ������      D  , ,  ������  �����%  �r���%  �r����  ������      D  , ,  � ����  � ���%  �����%  ������  � ����      D  , ,  �x����  �x���%  ����%  �����  �x����      D  , ,  ������  �����%  �R���%  �R����  ������      D  , ,  �����  ����%  �����%  ������  �����      D  , ,  �X����  �X���%  �����%  ������  �X����      D  , ,  ������  �����9  �:���9  �:����  ������      D  , ,  �s���y  �s���  �	���  �	���y  �s���y      D  , ,  �����y  �����  �W���  �W���y  �����y      D  , ,  ����y  ����  �����  �����y  ����y      D  , ,  �]���y  �]���  �����  �����y  �]���y      D  , ,  �����y  �����  �A���  �A���y  �����y      D  , ,  �����y  �����  �����  �����y  �����y      D  , ,  �G���y  �G���  �����  �����y  �G���y      D  , ,  �����y  �����  �+���  �+���y  �����y      D  , ,  �����y  �����  �y���  �y���y  �����y      D  , ,  �1���y  �1���  �����  �����y  �1���y      D  , ,  ����y  ����  ����  ����y  ����y      D  , ,  �s���9  �s����  �	����  �	���9  �s���9      D  , ,  �����9  ������  �W����  �W���9  �����9      D  , ,  ����9  �����  ������  �����9  ����9      D  , ,  �]���9  �]����  ������  �����9  �]���9      D  , ,  �����9  ������  �A����  �A���9  �����9      D  , ,  �����9  ������  ������  �����9  �����9      D  , ,  �G���9  �G����  ������  �����9  �G���9      D  , ,  �����9  ������  �+����  �+���9  �����9      D  , ,  �����9  ������  �y����  �y���9  �����9      D  , ,  �1���9  �1����  ������  �����9  �1���9      D  , ,  ������  �����9  �~���9  �~����  ������      D  , ,  �@����  �@���9  �����9  ������  �@����      D  , ,  ������  �����9  ����9  �����  ������      D  , ,  ������  �����9  �r���9  �r����  ������      D  , ,  � ����  � ���9  �����9  ������  � ����      D  , ,  �x����  �x���9  ����9  �����  �x����      D  , ,  ������  �����9  �R���9  �R����  ������      D  , ,  �����  ����9  �����9  ������  �����      D  , ,  �X����  �X���9  �����9  ������  �X����      D  , ,  �X���#  �X����  ������  �����#  �X���#      D  , ,  �����  ����e  �����e  ������  �����      D  , ,  �l����  �l���e  ����e  �����  �l����      D  , ,  ������  �����e  �F���e  �F����  ������      D  , ,  �����  ����e  �����e  ������  �����      D  , ,  �L����  �L���e  �����e  ������  �L����      D  , ,  ~@����  ~@���y  ~����y  ~�����  ~@����      D  , ,  ������  �����y  �.���y  �.����  ������      D  , ,  ������  �����y  �r���y  �r����  ������      D  , ,  �4����  �4���y  �����y  ������  �4����      D  , ,  �x����  �x���y  ����y  �����  �x����      D  , ,  ������  �����y  �f���y  �f����  ������      D  , ,  �����  ����y  �����y  ������  �����      D  , ,  �l����  �l���y  ����y  �����  �l����      D  , ,  ������  �����y  �F���y  �F����  ������      D  , ,  �����  ����y  �����y  ������  �����      D  , ,  �L����  �L���y  �����y  ������  �L����      D  , ,  �4���#  �4����  ������  �����#  �4���#      D  , ,  }���9  }����  }�����  }����9  }���9      D  , ,  g���9  g����  �����  ����9  g���9      D  , ,  �����9  ������  �K����  �K���9  �����9      D  , ,  ~@���  ~@����  ~�����  ~����  ~@���      D  , ,  ~@����  ~@���%  ~����%  ~�����  ~@����      D  , ,  ������  �����%  �.���%  �.����  ������      D  , ,  ������  �����%  �r���%  �r����  ������      D  , ,  �4����  �4���%  �����%  ������  �4����      D  , ,  �x����  �x���%  ����%  �����  �x����      D  , ,  ������  �����%  �f���%  �f����  ������      D  , ,  �����  ����%  �����%  ������  �����      D  , ,  �l����  �l���%  ����%  �����  �l����      D  , ,  ������  �����%  �F���%  �F����  ������      D  , ,  �����  ����%  �����%  ������  �����      D  , ,  �L����  �L���%  �����%  ������  �L����      D  , ,  �����  ������  �.����  �.���  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  �4���  �4����  ������  �����  �4���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �f����  �f���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �l���  �l����  �����  ����  �l���      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  ~@����  ~@���9  ~����9  ~�����  ~@����      D  , ,  ������  �����9  �.���9  �.����  ������      D  , ,  ������  �����9  �r���9  �r����  ������      D  , ,  �4����  �4���9  �����9  ������  �4����      D  , ,  �x����  �x���9  ����9  �����  �x����      D  , ,  ������  �����9  �f���9  �f����  ������      D  , ,  �����  ����9  �����9  ������  �����      D  , ,  �l����  �l���9  ����9  �����  �l����      D  , ,  ������  �����9  �F���9  �F����  ������      D  , ,  �����  ����9  �����9  ������  �����      D  , ,  �L����  �L���9  �����9  ������  �L����      D  , ,  ����9  �����  ������  �����9  ����9      D  , ,  �Q���9  �Q����  ������  �����9  �Q���9      D  , ,  �����9  ������  �5����  �5���9  �����9      D  , ,  �����9  ������  ������  �����9  �����9      D  , ,  �;���9  �;����  ������  �����9  �;���9      D  , ,  �����9  ������  �����  ����9  �����9      D  , ,  �����9  ������  �m����  �m���9  �����9      D  , ,  �%���9  �%����  ������  �����9  �%���9      D  , ,  }���y  }���  }����  }����y  }���y      D  , ,  g���y  g���  ����  ����y  g���y      D  , ,  �����y  �����  �K���  �K���y  �����y      D  , ,  ����y  ����  �����  �����y  ����y      D  , ,  �Q���y  �Q���  �����  �����y  �Q���y      D  , ,  �����y  �����  �5���  �5���y  �����y      D  , ,  �����y  �����  �����  �����y  �����y      D  , ,  �;���y  �;���  �����  �����y  �;���y      D  , ,  �x���#  �x����  �����  ����#  �x���#      D  , ,  �����#  ������  �f����  �f���#  �����#      D  , ,  ����#  �����  ������  �����#  ����#      D  , ,  �l���#  �l����  �����  ����#  �l���#      D  , ,  �����#  ������  �F����  �F���#  �����#      D  , ,  ����#  �����  ������  �����#  ����#      D  , ,  �L���#  �L����  ������  �����#  �L���#      D  , ,  �����y  �����  ����  ����y  �����y      D  , ,  �����y  �����  �m���  �m���y  �����y      D  , ,  �%���y  �%���  �����  �����y  �%���y      D  , ,  ~@����  ~@���e  ~����e  ~�����  ~@����      D  , ,  ������  �����e  �.���e  �.����  ������      D  , ,  ������  �����e  �r���e  �r����  ������      D  , ,  �4����  �4���e  �����e  ������  �4����      D  , ,  �x����  �x���e  ����e  �����  �x����      D  , ,  ������  �����e  �f���e  �f����  ������      D  , ,  ~@���#  ~@����  ~�����  ~����#  ~@���#      D  , ,  �����#  ������  �.����  �.���#  �����#      D  , ,  �����#  ������  �r����  �r���#  �����#      D  , ,  �����=  ������  �r����  �r���=  �����=      D  , ,  �x���=  �x����  �����  ����=  �x���=      D  , ,  ����=  �����  ������  �����=  ����=      D  , ,  �����=  ������  �F����  �F���=  �����=      D  , ,  �L���=  �L����  ������  �����=  �L���=      D  , ,  �L����  �L���%  �����%  ������  �L����      D  , ,  �L����  �L���e  �����e  ������  �L����      D  , ,  ~@����  ~@���e  ~����e  ~�����  ~@����      D  , ,  ������  �����e  �.���e  �.����  ������      D  , ,  ������  �����e  �r���e  �r����  ������      D  , ,  �4����  �4���e  �����e  ������  �4����      D  , ,  �x����  �x���e  ����e  �����  �x����      D  , ,  ������  �����e  �f���e  �f����  ������      D  , ,  ~@����  ~@����  ~�����  ~�����  ~@����      D  , ,  ������  ������  �r����  �r����  ������      D  , ,  �x����  �x����  �����  �����  �x����      D  , ,  �����  �����  ������  ������  �����      D  , ,  ������  ������  �F����  �F����  ������      D  , ,  �L����  �L����  ������  ������  �L����      D  , ,  �����  ����e  �����e  ������  �����      D  , ,  �l����  �l���e  ����e  �����  �l����      D  , ,  ������  �����e  �F���e  �F����  ������      D  , ,  �����  ����e  �����e  ������  �����      D  , ,  ~@����  ~@���%  ~����%  ~�����  ~@����      D  , ,  ������  �����%  �.���%  �.����  ������      D  , ,  ~@���O  ~@����  ~�����  ~����O  ~@���O      D  , ,  �����O  ������  �.����  �.���O  �����O      D  , ,  �����O  ������  �r����  �r���O  �����O      D  , ,  �4���O  �4����  ������  �����O  �4���O      D  , ,  �x���O  �x����  �����  ����O  �x���O      D  , ,  �����O  ������  �f����  �f���O  �����O      D  , ,  ����O  �����  ������  �����O  ����O      D  , ,  �l���O  �l����  �����  ����O  �l���O      D  , ,  �����O  ������  �F����  �F���O  �����O      D  , ,  ����O  �����  ������  �����O  ����O      D  , ,  �L���O  �L����  ������  �����O  �L���O      D  , ,  ~@����  ~@���S  ~����S  ~�����  ~@����      D  , ,  ������  �����S  �r���S  �r����  ������      D  , ,  �x����  �x���S  ����S  �����  �x����      D  , ,  �����  ����S  �����S  ������  �����      D  , ,  ������  �����S  �F���S  �F����  ������      D  , ,  �L����  �L���S  �����S  ������  �L����      D  , ,  ~@���}  ~@���  ~����  ~����}  ~@���}      D  , ,  �����}  �����  �r���  �r���}  �����}      D  , ,  �x���}  �x���  ����  ����}  �x���}      D  , ,  ����}  ����  �����  �����}  ����}      D  , ,  �����}  �����  �F���  �F���}  �����}      D  , ,  �L���}  �L���  �����  �����}  �L���}      D  , ,  ������  �����%  �r���%  �r����  ������      D  , ,  �4����  �4���%  �����%  ������  �4����      D  , ,  �x����  �x���%  ����%  �����  �x����      D  , ,  ������  �����%  �f���%  �f����  ������      D  , ,  �����  ����%  �����%  ������  �����      D  , ,  �l����  �l���%  ����%  �����  �l����      D  , ,  ~@���  ~@����  ~�����  ~����  ~@���      D  , ,  �����  ������  �.����  �.���  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  �4���  �4����  ������  �����  �4���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �f����  �f���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �l���  �l����  �����  ����  �l���      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  ������  �����%  �F���%  �F����  ������      D  , ,  �����  ����%  �����%  ������  �����      D  , ,  ~@���=  ~@����  ~�����  ~����=  ~@���=      D  , ,  ������  �����%  �R���%  �R����  ������      D  , ,  �����  ����%  �����%  ������  �����      D  , ,  �X����  �X���%  �����%  ������  �X����      D  , ,  ������  �����e  �~���e  �~����  ������      D  , ,  �@����  �@���e  �����e  ������  �@����      D  , ,  ������  �����e  ����e  �����  ������      D  , ,  ������  �����e  �r���e  �r����  ������      D  , ,  �����O  ������  �:����  �:���O  �����O      D  , ,  �����O  ������  �~����  �~���O  �����O      D  , ,  �@���O  �@����  ������  �����O  �@���O      D  , ,  �����O  ������  �����  ����O  �����O      D  , ,  �����O  ������  �r����  �r���O  �����O      D  , ,  � ���O  � ����  ������  �����O  � ���O      D  , ,  �����=  ������  �~����  �~���=  �����=      D  , ,  �����=  ������  �����  ����=  �����=      D  , ,  � ���=  � ����  ������  �����=  � ���=      D  , ,  �����=  ������  �R����  �R���=  �����=      D  , ,  �X���=  �X����  ������  �����=  �X���=      D  , ,  �x���O  �x����  �����  ����O  �x���O      D  , ,  �����O  ������  �R����  �R���O  �����O      D  , ,  ����O  �����  ������  �����O  ����O      D  , ,  �X���O  �X����  ������  �����O  �X���O      D  , ,  � ����  � ���e  �����e  ������  � ����      D  , ,  �x����  �x���e  ����e  �����  �x����      D  , ,  ������  �����e  �R���e  �R����  ������      D  , ,  �����  ����e  �����e  ������  �����      D  , ,  �X����  �X���e  �����e  ������  �X����      D  , ,  ������  �����e  �:���e  �:����  ������      D  , ,  ������  �����S  �~���S  �~����  ������      D  , ,  ������  �����S  ����S  �����  ������      D  , ,  � ����  � ���S  �����S  ������  � ����      D  , ,  ������  �����S  �R���S  �R����  ������      D  , ,  ������  ������  �~����  �~����  ������      D  , ,  ������  ������  �����  �����  ������      D  , ,  � ����  � ����  ������  ������  � ����      D  , ,  ������  ������  �R����  �R����  ������      D  , ,  �X����  �X����  ������  ������  �X����      D  , ,  �X����  �X���S  �����S  ������  �X����      D  , ,  ������  �����%  �:���%  �:����  ������      D  , ,  ������  �����%  �~���%  �~����  ������      D  , ,  �@����  �@���%  �����%  ������  �@����      D  , ,  ������  �����%  ����%  �����  ������      D  , ,  ������  �����%  �r���%  �r����  ������      D  , ,  � ����  � ���%  �����%  ������  � ����      D  , ,  �����}  �����  �~���  �~���}  �����}      D  , ,  �����}  �����  ����  ����}  �����}      D  , ,  � ���}  � ���  �����  �����}  � ���}      D  , ,  �����  ������  �:����  �:���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �@���  �@����  ������  �����  �@���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �R����  �R���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  �����}  �����  �R���  �R���}  �����}      D  , ,  �X���}  �X���  �����  �����}  �X���}      D  , ,  �x����  �x���%  ����%  �����  �x����      D  , ,  c����9  c�����  dU����  dU���9  c����9      D  , ,  ]����O  ]�����  ^�����  ^����O  ]����O      D  , ,  `T���O  `T����  `�����  `����O  `T���O      D  , ,  b����O  b�����  c.����  c.���O  b����O      D  , ,  d����O  d�����  e�����  e����O  d����O      D  , ,  g4���O  g4����  g�����  g����O  g4���O      D  , ,  i����O  i�����  j"����  j"���O  i����O      D  , ,  k����O  k�����  lf����  lf���O  k����O      D  , ,  n(���O  n(����  n�����  n����O  n(���O      D  , ,  pl���O  pl����  q����  q���O  pl���O      D  , ,  r����O  r�����  sZ����  sZ���O  r����O      D  , ,  u���O  u����  u�����  u����O  u���O      D  , ,  w`���O  w`����  w�����  w����O  w`���O      D  , ,  y����O  y�����  z:����  z:���O  y����O      D  , ,  {����O  {�����  |�����  |����O  {����O      D  , ,  c����y  c����  dU���  dU���y  c����y      D  , ,  k�����  k����9  lf���9  lf����  k�����      D  , ,  n(����  n(���9  n����9  n�����  n(����      D  , ,  pl����  pl���9  q���9  q����  pl����      D  , ,  r�����  r����9  sZ���9  sZ����  r�����      D  , ,  d�����  d����%  e����%  e�����  d�����      D  , ,  g4����  g4���%  g����%  g�����  g4����      D  , ,  i�����  i����%  j"���%  j"����  i�����      D  , ,  k�����  k����%  lf���%  lf����  k�����      D  , ,  n(����  n(���%  n����%  n�����  n(����      D  , ,  pl����  pl���%  q���%  q����  pl����      D  , ,  r�����  r����%  sZ���%  sZ����  r�����      D  , ,  u����  u���%  u����%  u�����  u����      D  , ,  w`����  w`���%  w����%  w�����  w`����      D  , ,  y�����  y����%  z:���%  z:����  y�����      D  , ,  {�����  {����%  |����%  |�����  {�����      D  , ,  i�����  i����y  j"���y  j"����  i�����      D  , ,  k�����  k����y  lf���y  lf����  k�����      D  , ,  n(����  n(���y  n����y  n�����  n(����      D  , ,  pl����  pl���y  q���y  q����  pl����      D  , ,  r�����  r����y  sZ���y  sZ����  r�����      D  , ,  u����  u���y  u����y  u�����  u����      D  , ,  w`����  w`���y  w����y  w�����  w`����      D  , ,  y�����  y����y  z:���y  z:����  y�����      D  , ,  {�����  {����y  |����y  |�����  {�����      D  , ,  d�����  d����e  e����e  e�����  d�����      D  , ,  f���9  f����  f�����  f����9  f���9      D  , ,  h[���9  h[����  h�����  h����9  h[���9      D  , ,  u����  u���9  u����9  u�����  u����      D  , ,  w`����  w`���9  w����9  w�����  w`����      D  , ,  y�����  y����9  z:���9  z:����  y�����      D  , ,  {�����  {����9  |����9  |�����  {�����      D  , ,  oE���y  oE���  o����  o����y  oE���y      D  , ,  q����y  q����  r)���  r)���y  q����y      D  , ,  s����y  s����  tw���  tw���y  s����y      D  , ,  v/���y  v/���  v����  v����y  v/���y      D  , ,  g4����  g4���e  g����e  g�����  g4����      D  , ,  i�����  i����e  j"���e  j"����  i�����      D  , ,  k�����  k����e  lf���e  lf����  k�����      D  , ,  n(����  n(���e  n����e  n�����  n(����      D  , ,  pl����  pl���e  q���e  q����  pl����      D  , ,  r�����  r����e  sZ���e  sZ����  r�����      D  , ,  u����  u���e  u����e  u�����  u����      D  , ,  w`����  w`���e  w����e  w�����  w`����      D  , ,  y�����  y����e  z:���e  z:����  y�����      D  , ,  {�����  {����e  |����e  |�����  {�����      D  , ,  d�����  d����y  e����y  e�����  d�����      D  , ,  g4����  g4���y  g����y  g�����  g4����      D  , ,  d�����  d����9  e����9  e�����  d�����      D  , ,  g4����  g4���9  g����9  g�����  g4����      D  , ,  d����  d�����  e�����  e����  d����      D  , ,  g4���  g4����  g�����  g����  g4���      D  , ,  i����  i�����  j"����  j"���  i����      D  , ,  k����  k�����  lf����  lf���  k����      D  , ,  n(���  n(����  n�����  n����  n(���      D  , ,  pl���  pl����  q����  q���  pl���      D  , ,  r����  r�����  sZ����  sZ���  r����      D  , ,  u���  u����  u�����  u����  u���      D  , ,  w`���  w`����  w�����  w����  w`���      D  , ,  y����  y�����  z:����  z:���  y����      D  , ,  {����  {�����  |�����  |����  {����      D  , ,  j����9  j�����  k?����  k?���9  j����9      D  , ,  l����9  l�����  m�����  m����9  l����9      D  , ,  oE���9  oE����  o�����  o����9  oE���9      D  , ,  q����9  q�����  r)����  r)���9  q����9      D  , ,  s����9  s�����  tw����  tw���9  s����9      D  , ,  v/���9  v/����  v�����  v����9  v/���9      D  , ,  x}���9  x}����  y����  y���9  x}���9      D  , ,  z����9  z�����  {a����  {a���9  z����9      D  , ,  d����#  d�����  e�����  e����#  d����#      D  , ,  g4���#  g4����  g�����  g����#  g4���#      D  , ,  i����#  i�����  j"����  j"���#  i����#      D  , ,  k����#  k�����  lf����  lf���#  k����#      D  , ,  n(���#  n(����  n�����  n����#  n(���#      D  , ,  x}���y  x}���  y���  y���y  x}���y      D  , ,  z����y  z����  {a���  {a���y  z����y      D  , ,  pl���#  pl����  q����  q���#  pl���#      D  , ,  r����#  r�����  sZ����  sZ���#  r����#      D  , ,  u���#  u����  u�����  u����#  u���#      D  , ,  w`���#  w`����  w�����  w����#  w`���#      D  , ,  y����#  y�����  z:����  z:���#  y����#      D  , ,  {����#  {�����  |�����  |����#  {����#      D  , ,  i�����  i����9  j"���9  j"����  i�����      D  , ,  f���y  f���  f����  f����y  f���y      D  , ,  h[���y  h[���  h����  h����y  h[���y      D  , ,  j����y  j����  k?���  k?���y  j����y      D  , ,  l����y  l����  m����  m����y  l����y      D  , ,  `T����  `T���%  `����%  `�����  `T����      D  , ,  ]�����  ]����y  ^����y  ^�����  ]�����      D  , ,  b�����  b����y  c.���y  c.����  b�����      D  , ,  `T����  `T���y  `����y  `�����  `T����      D  , ,  ]����  ]�����  ^�����  ^����  ]����      D  , ,  `T���  `T����  `�����  `����  `T���      D  , ,  b����  b�����  c.����  c.���  b����      D  , ,  _#���9  _#����  _�����  _����9  _#���9      D  , ,  aq���9  aq����  b����  b���9  aq���9      D  , ,  b�����  b����%  c.���%  c.����  b�����      D  , ,  b�����  b����9  c.���9  c.����  b�����      D  , ,  ]�����  ]����e  ^����e  ^�����  ]�����      D  , ,  `T����  `T���e  `����e  `�����  `T����      D  , ,  _#���y  _#���  _����  _����y  _#���y      D  , ,  aq���y  aq���  b���  b���y  aq���y      D  , ,  b�����  b����e  c.���e  c.����  b�����      D  , ,  b����#  b�����  c.����  c.���#  b����#      D  , ,  ]�����  ]����9  ^����9  ^�����  ]�����      D  , ,  ]����#  ]�����  ^�����  ^����#  ]����#      D  , ,  `T����  `T���9  `����9  `�����  `T����      D  , ,  `T���#  `T����  `�����  `����#  `T���#      D  , ,  ]�����  ]����%  ^����%  ^�����  ]�����      D  , ,  `T����  `T���%  `����%  `�����  `T����      D  , ,  ]�����  ]����S  ^����S  ^�����  ]�����      D  , ,  b�����  b����S  c.���S  c.����  b�����      D  , ,  ]�����  ]�����  ^�����  ^�����  ]�����      D  , ,  b�����  b�����  c.����  c.����  b�����      D  , ,  b�����  b����%  c.���%  c.����  b�����      D  , ,  ]����  ]�����  ^�����  ^����  ]����      D  , ,  `T���  `T����  `�����  `����  `T���      D  , ,  b����  b�����  c.����  c.���  b����      D  , ,  ]�����  ]����%  ^����%  ^�����  ]�����      D  , ,  ]����O  ]�����  ^�����  ^����O  ]����O      D  , ,  `T���O  `T����  `�����  `����O  `T���O      D  , ,  b����O  b�����  c.����  c.���O  b����O      D  , ,  ]����}  ]����  ^����  ^����}  ]����}      D  , ,  b����}  b����  c.���  c.���}  b����}      D  , ,  ]����=  ]�����  ^�����  ^����=  ]����=      D  , ,  b����=  b�����  c.����  c.���=  b����=      D  , ,  ]�����  ]����e  ^����e  ^�����  ]�����      D  , ,  `T����  `T���e  `����e  `�����  `T����      D  , ,  b�����  b����e  c.���e  c.����  b�����      D  , ,  y����}  y����  z:���  z:���}  y����}      D  , ,  n(����  n(���%  n����%  n�����  n(����      D  , ,  pl����  pl���%  q���%  q����  pl����      D  , ,  y����=  y�����  z:����  z:���=  y����=      D  , ,  n(����  n(���e  n����e  n�����  n(����      D  , ,  pl����  pl���e  q���e  q����  pl����      D  , ,  r�����  r����e  sZ���e  sZ����  r�����      D  , ,  g4����  g4����  g�����  g�����  g4����      D  , ,  k�����  k�����  lf����  lf����  k�����      D  , ,  g4����  g4���S  g����S  g�����  g4����      D  , ,  d����  d�����  e�����  e����  d����      D  , ,  g4���  g4����  g�����  g����  g4���      D  , ,  i����  i�����  j"����  j"���  i����      D  , ,  k����  k�����  lf����  lf���  k����      D  , ,  n(���  n(����  n�����  n����  n(���      D  , ,  pl���  pl����  q����  q���  pl���      D  , ,  r����  r�����  sZ����  sZ���  r����      D  , ,  u���  u����  u�����  u����  u���      D  , ,  w`���  w`����  w�����  w����  w`���      D  , ,  y����  y�����  z:����  z:���  y����      D  , ,  {����  {�����  |�����  |����  {����      D  , ,  k�����  k����S  lf���S  lf����  k�����      D  , ,  u����  u���e  u����e  u�����  u����      D  , ,  w`����  w`���e  w����e  w�����  w`����      D  , ,  y�����  y����e  z:���e  z:����  y�����      D  , ,  d����O  d�����  e�����  e����O  d����O      D  , ,  g4���O  g4����  g�����  g����O  g4���O      D  , ,  i����O  i�����  j"����  j"���O  i����O      D  , ,  k����O  k�����  lf����  lf���O  k����O      D  , ,  n(���O  n(����  n�����  n����O  n(���O      D  , ,  pl���O  pl����  q����  q���O  pl���O      D  , ,  r����O  r�����  sZ����  sZ���O  r����O      D  , ,  u���O  u����  u�����  u����O  u���O      D  , ,  w`���O  w`����  w�����  w����O  w`���O      D  , ,  y����O  y�����  z:����  z:���O  y����O      D  , ,  {����O  {�����  |�����  |����O  {����O      D  , ,  {�����  {����e  |����e  |�����  {�����      D  , ,  pl����  pl���S  q���S  q����  pl����      D  , ,  i�����  i����e  j"���e  j"����  i�����      D  , ,  k�����  k����e  lf���e  lf����  k�����      D  , ,  u����  u���S  u����S  u�����  u����      D  , ,  y�����  y����S  z:���S  z:����  y�����      D  , ,  r�����  r����%  sZ���%  sZ����  r�����      D  , ,  u����  u���%  u����%  u�����  u����      D  , ,  w`����  w`���%  w����%  w�����  w`����      D  , ,  y�����  y����%  z:���%  z:����  y�����      D  , ,  {�����  {����%  |����%  |�����  {�����      D  , ,  pl����  pl����  q����  q����  pl����      D  , ,  g4���=  g4����  g�����  g����=  g4���=      D  , ,  u����  u����  u�����  u�����  u����      D  , ,  y�����  y�����  z:����  z:����  y�����      D  , ,  g4����  g4���e  g����e  g�����  g4����      D  , ,  k����=  k�����  lf����  lf���=  k����=      D  , ,  pl���=  pl����  q����  q���=  pl���=      D  , ,  u���=  u����  u�����  u����=  u���=      D  , ,  d�����  d����%  e����%  e�����  d�����      D  , ,  g4����  g4���%  g����%  g�����  g4����      D  , ,  i�����  i����%  j"���%  j"����  i�����      D  , ,  k�����  k����%  lf���%  lf����  k�����      D  , ,  g4���}  g4���  g����  g����}  g4���}      D  , ,  k����}  k����  lf���  lf���}  k����}      D  , ,  pl���}  pl���  q���  q���}  pl���}      D  , ,  u���}  u���  u����  u����}  u���}      D  , ,  d�����  d����e  e����e  e�����  d�����      D  , ,  ]�����  ]����/  ^����/  ^�����  ]�����      D  , ,  `T����  `T���/  `����/  `�����  `T����      D  , ,  b�����  b����/  c.���/  c.����  b�����      D  , ,  d�����  d����/  e����/  e�����  d�����      D  , ,  g4����  g4���/  g����/  g�����  g4����      D  , ,  i�����  i����/  j"���/  j"����  i�����      D  , ,  k�����  k����/  lf���/  lf����  k�����      D  , ,  n(����  n(���/  n����/  n�����  n(����      D  , ,  pl����  pl���/  q���/  q����  pl����      D  , ,  r�����  r����/  sZ���/  sZ����  r�����      D  , ,  u����  u���/  u����/  u�����  u����      D  , ,  w`����  w`���/  w����/  w�����  w`����      D  , ,  y�����  y����/  z:���/  z:����  y�����      D  , ,  {�����  {����/  |����/  |�����  {�����      D  , ,  c����o  c����  dU���  dU���o  c����o      D  , ,  c����/  c�����  dU����  dU���/  c����/      D  , ,  {����  {�����  |�����  |����  {����      D  , ,  pl���  pl����  q����  q���  pl���      D  , ,  r����  r�����  sZ����  sZ���  r����      D  , ,  u���  u����  u�����  u����  u���      D  , ,  w`���  w`����  w�����  w����  w`���      D  , ,  y����  y�����  z:����  z:���  y����      D  , ,  {����  {�����  |�����  |����  {����      D  , ,  d����Y  d�����  e�����  e����Y  d����Y      D  , ,  g4���Y  g4����  g�����  g����Y  g4���Y      D  , ,  i����Y  i�����  j"����  j"���Y  i����Y      D  , ,  d�����  d����/  e����/  e�����  d�����      D  , ,  g4����  g4���/  g����/  g�����  g4����      D  , ,  i�����  i����/  j"���/  j"����  i�����      D  , ,  d�����  d����o  e����o  e�����  d�����      D  , ,  g4����  g4���o  g����o  g�����  g4����      D  , ,  i�����  i����o  j"���o  j"����  i�����      D  , ,  k�����  k����o  lf���o  lf����  k�����      D  , ,  n(����  n(���o  n����o  n�����  n(����      D  , ,  pl����  pl���o  q���o  q����  pl����      D  , ,  r�����  r����o  sZ���o  sZ����  r�����      D  , ,  u����  u���o  u����o  u�����  u����      D  , ,  w`����  w`���o  w����o  w�����  w`����      D  , ,  y�����  y����o  z:���o  z:����  y�����      D  , ,  {�����  {����o  |����o  |�����  {�����      D  , ,  k�����  k����/  lf���/  lf����  k�����      D  , ,  n(����  n(���/  n����/  n�����  n(����      D  , ,  pl����  pl���/  q���/  q����  pl����      D  , ,  r�����  r����/  sZ���/  sZ����  r�����      D  , ,  u����  u���/  u����/  u�����  u����      D  , ,  w`����  w`���/  w����/  w�����  w`����      D  , ,  y�����  y����/  z:���/  z:����  y�����      D  , ,  {�����  {����/  |����/  |�����  {�����      D  , ,  k����Y  k�����  lf����  lf���Y  k����Y      D  , ,  n(���Y  n(����  n�����  n����Y  n(���Y      D  , ,  pl���Y  pl����  q����  q���Y  pl���Y      D  , ,  r����Y  r�����  sZ����  sZ���Y  r����Y      D  , ,  u���Y  u����  u�����  u����Y  u���Y      D  , ,  w`���Y  w`����  w�����  w����Y  w`���Y      D  , ,  y����Y  y�����  z:����  z:���Y  y����Y      D  , ,  {����Y  {�����  |�����  |����Y  {����Y      D  , ,  {�����  {����o  |����o  |�����  {�����      D  , ,  d����  d�����  e�����  e����  d����      D  , ,  g4���  g4����  g�����  g����  g4���      D  , ,  i����  i�����  j"����  j"���  i����      D  , ,  k����  k�����  lf����  lf���  k����      D  , ,  n(���  n(����  n�����  n����  n(���      D  , ,  d����  d�����  e�����  e����  d����      D  , ,  g4���  g4����  g�����  g����  g4���      D  , ,  i����  i�����  j"����  j"���  i����      D  , ,  k����  k�����  lf����  lf���  k����      D  , ,  n(���  n(����  n�����  n����  n(���      D  , ,  pl���  pl����  q����  q���  pl���      D  , ,  r����  r�����  sZ����  sZ���  r����      D  , ,  u���  u����  u�����  u����  u���      D  , ,  d�����  d����o  e����o  e�����  d�����      D  , ,  d����Y  d�����  e�����  e����Y  d����Y      D  , ,  g4���Y  g4����  g�����  g����Y  g4���Y      D  , ,  i����Y  i�����  j"����  j"���Y  i����Y      D  , ,  k����Y  k�����  lf����  lf���Y  k����Y      D  , ,  n(���Y  n(����  n�����  n����Y  n(���Y      D  , ,  w`���  w`����  w�����  w����  w`���      D  , ,  pl���Y  pl����  q����  q���Y  pl���Y      D  , ,  r����Y  r�����  sZ����  sZ���Y  r����Y      D  , ,  u���Y  u����  u�����  u����Y  u���Y      D  , ,  w`���Y  w`����  w�����  w����Y  w`���Y      D  , ,  y����Y  y�����  z:����  z:���Y  y����Y      D  , ,  {����Y  {�����  |�����  |����Y  {����Y      D  , ,  g4����  g4���o  g����o  g�����  g4����      D  , ,  i�����  i����o  j"���o  j"����  i�����      D  , ,  k�����  k����o  lf���o  lf����  k�����      D  , ,  n(����  n(���o  n����o  n�����  n(����      D  , ,  pl����  pl���o  q���o  q����  pl����      D  , ,  r�����  r����o  sZ���o  sZ����  r�����      D  , ,  u����  u���o  u����o  u�����  u����      D  , ,  w`����  w`���o  w����o  w�����  w`����      D  , ,  y�����  y����o  z:���o  z:����  y�����      D  , ,  y����  y�����  z:����  z:���  y����      D  , ,  b�����  b����o  c.���o  c.����  b�����      D  , ,  `T���  `T����  `�����  `����  `T���      D  , ,  b����  b�����  c.����  c.���  b����      D  , ,  ]�����  ]����/  ^����/  ^�����  ]�����      D  , ,  `T����  `T���/  `����/  `�����  `T����      D  , ,  b�����  b����/  c.���/  c.����  b�����      D  , ,  b����  b�����  c.����  c.���  b����      D  , ,  b����Y  b�����  c.����  c.���Y  b����Y      D  , ,  ]����  ]�����  ^�����  ^����  ]����      D  , ,  ]����Y  ]�����  ^�����  ^����Y  ]����Y      D  , ,  `T���Y  `T����  `�����  `����Y  `T���Y      D  , ,  ]����  ]�����  ^�����  ^����  ]����      D  , ,  `T���  `T����  `�����  `����  `T���      D  , ,  ]�����  ]����o  ^����o  ^�����  ]�����      D  , ,  `T����  `T���o  `����o  `�����  `T����      D  , ,  b�����  b����o  c.���o  c.����  b�����      D  , ,  ]�����  ]����o  ^����o  ^�����  ]�����      D  , ,  ]����Y  ]�����  ^�����  ^����Y  ]����Y      D  , ,  `T���Y  `T����  `�����  `����Y  `T���Y      D  , ,  b����Y  b�����  c.����  c.���Y  b����Y      D  , ,  `T����  `T���o  `����o  `�����  `T����      D  , ,  ]����  ]�����  ^�����  ^����  ]����      D  , ,  _#���o  _#���  _����  _����o  _#���o      D  , ,  aq���o  aq���  b���  b���o  aq���o      D  , ,  ]�����  ]����[  ^����[  ^�����  ]�����      D  , ,  ]�����  ]����  ^����  ^�����  ]�����      D  , ,  ]����E  ]�����  ^�����  ^����E  ]����E      D  , ,  `T���E  `T����  `�����  `����E  `T���E      D  , ,  b����E  b�����  c.����  c.���E  b����E      D  , ,  `T����  `T���  `����  `�����  `T����      D  , ,  b�����  b����  c.���  c.����  b�����      D  , ,  `T����  `T���[  `����[  `�����  `T����      D  , ,  b�����  b����[  c.���[  c.����  b�����      D  , ,  ]����  ]�����  ^�����  ^����  ]����      D  , ,  `T���  `T����  `�����  `����  `T���      D  , ,  b����  b�����  c.����  c.���  b����      D  , ,  `T���  `T����  `�����  `����  `T���      D  , ,  ]�����  ]����[  ^����[  ^�����  ]�����      D  , ,  `T����  `T���[  `����[  `�����  `T����      D  , ,  b�����  b����[  c.���[  c.����  b�����      D  , ,  _#���/  _#����  _�����  _����/  _#���/      D  , ,  aq���/  aq����  b����  b���/  aq���/      D  , ,  b����  b�����  c.����  c.���  b����      D  , ,  d�����  d����  e����  e�����  d�����      D  , ,  g4����  g4���  g����  g�����  g4����      D  , ,  i�����  i����  j"���  j"����  i�����      D  , ,  k�����  k����  lf���  lf����  k�����      D  , ,  n(����  n(���  n����  n�����  n(����      D  , ,  pl����  pl���  q���  q����  pl����      D  , ,  r�����  r����  sZ���  sZ����  r�����      D  , ,  u����  u���  u����  u�����  u����      D  , ,  w`����  w`���  w����  w�����  w`����      D  , ,  d����  d�����  e�����  e����  d����      D  , ,  g4���  g4����  g�����  g����  g4���      D  , ,  i����  i�����  j"����  j"���  i����      D  , ,  k����  k�����  lf����  lf���  k����      D  , ,  n(���  n(����  n�����  n����  n(���      D  , ,  pl���  pl����  q����  q���  pl���      D  , ,  r����  r�����  sZ����  sZ���  r����      D  , ,  u���  u����  u�����  u����  u���      D  , ,  w`���  w`����  w�����  w����  w`���      D  , ,  y����  y�����  z:����  z:���  y����      D  , ,  {����  {�����  |�����  |����  {����      D  , ,  y�����  y����  z:���  z:����  y�����      D  , ,  {�����  {����  |����  |�����  {�����      D  , ,  g4����  g4���[  g����[  g�����  g4����      D  , ,  i�����  i����[  j"���[  j"����  i�����      D  , ,  k�����  k����[  lf���[  lf����  k�����      D  , ,  n(����  n(���[  n����[  n�����  n(����      D  , ,  pl����  pl���[  q���[  q����  pl����      D  , ,  r�����  r����[  sZ���[  sZ����  r�����      D  , ,  u����  u���[  u����[  u�����  u����      D  , ,  w`����  w`���[  w����[  w�����  w`����      D  , ,  y�����  y����[  z:���[  z:����  y�����      D  , ,  {�����  {����[  |����[  |�����  {�����      D  , ,  x}���/  x}����  y����  y���/  x}���/      D  , ,  z����/  z�����  {a����  {a���/  z����/      D  , ,  l����/  l�����  m�����  m����/  l����/      D  , ,  oE���/  oE����  o�����  o����/  oE���/      D  , ,  q����/  q�����  r)����  r)���/  q����/      D  , ,  s����/  s�����  tw����  tw���/  s����/      D  , ,  d����  d�����  e�����  e����  d����      D  , ,  d�����  d����[  e����[  e�����  d�����      D  , ,  g4����  g4���[  g����[  g�����  g4����      D  , ,  i�����  i����[  j"���[  j"����  i�����      D  , ,  k�����  k����[  lf���[  lf����  k�����      D  , ,  n(����  n(���[  n����[  n�����  n(����      D  , ,  pl����  pl���[  q���[  q����  pl����      D  , ,  r�����  r����[  sZ���[  sZ����  r�����      D  , ,  u����  u���[  u����[  u�����  u����      D  , ,  w`����  w`���[  w����[  w�����  w`����      D  , ,  y�����  y����[  z:���[  z:����  y�����      D  , ,  {�����  {����[  |����[  |�����  {�����      D  , ,  g4���  g4����  g�����  g����  g4���      D  , ,  i����  i�����  j"����  j"���  i����      D  , ,  d����E  d�����  e�����  e����E  d����E      D  , ,  g4���E  g4����  g�����  g����E  g4���E      D  , ,  i����E  i�����  j"����  j"���E  i����E      D  , ,  f���o  f���  f����  f����o  f���o      D  , ,  h[���o  h[���  h����  h����o  h[���o      D  , ,  j����o  j����  k?���  k?���o  j����o      D  , ,  l����o  l����  m����  m����o  l����o      D  , ,  oE���o  oE���  o����  o����o  oE���o      D  , ,  q����o  q����  r)���  r)���o  q����o      D  , ,  s����o  s����  tw���  tw���o  s����o      D  , ,  v/���o  v/���  v����  v����o  v/���o      D  , ,  x}���o  x}���  y���  y���o  x}���o      D  , ,  z����o  z����  {a���  {a���o  z����o      D  , ,  k����E  k�����  lf����  lf���E  k����E      D  , ,  n(���E  n(����  n�����  n����E  n(���E      D  , ,  pl���E  pl����  q����  q���E  pl���E      D  , ,  r����E  r�����  sZ����  sZ���E  r����E      D  , ,  u���E  u����  u�����  u����E  u���E      D  , ,  w`���E  w`����  w�����  w����E  w`���E      D  , ,  y����E  y�����  z:����  z:���E  y����E      D  , ,  {����E  {�����  |�����  |����E  {����E      D  , ,  k����  k�����  lf����  lf���  k����      D  , ,  n(���  n(����  n�����  n����  n(���      D  , ,  pl���  pl����  q����  q���  pl���      D  , ,  r����  r�����  sZ����  sZ���  r����      D  , ,  u���  u����  u�����  u����  u���      D  , ,  w`���  w`����  w�����  w����  w`���      D  , ,  y����  y�����  z:����  z:���  y����      D  , ,  {����  {�����  |�����  |����  {����      D  , ,  v/���/  v/����  v�����  v����/  v/���/      D  , ,  d�����  d����[  e����[  e�����  d�����      D  , ,  f���/  f����  f�����  f����/  f���/      D  , ,  h[���/  h[����  h�����  h����/  h[���/      D  , ,  j����/  j�����  k?����  k?���/  j����/      D  , ,  ~@����  ~@���/  ~����/  ~�����  ~@����      D  , ,  ������  �����/  �.���/  �.����  ������      D  , ,  ������  �����/  �r���/  �r����  ������      D  , ,  �4����  �4���/  �����/  ������  �4����      D  , ,  �x����  �x���/  ����/  �����  �x����      D  , ,  ������  �����/  �f���/  �f����  ������      D  , ,  �����  ����/  �����/  ������  �����      D  , ,  �l����  �l���/  ����/  �����  �l����      D  , ,  ������  �����/  �F���/  �F����  ������      D  , ,  �����  ����/  �����/  ������  �����      D  , ,  �L����  �L���/  �����/  ������  �L����      D  , ,  ������  �����/  �:���/  �:����  ������      D  , ,  ������  �����/  �~���/  �~����  ������      D  , ,  �@����  �@���/  �����/  ������  �@����      D  , ,  ������  �����/  ����/  �����  ������      D  , ,  ������  �����/  �r���/  �r����  ������      D  , ,  � ����  � ���/  �����/  ������  � ����      D  , ,  �x����  �x���/  ����/  �����  �x����      D  , ,  ������  �����/  �R���/  �R����  ������      D  , ,  �����  ����/  �����/  ������  �����      D  , ,  �X����  �X���/  �����/  ������  �X����      D  , ,  � ����  � ���o  �����o  ������  � ����      D  , ,  �x����  �x���o  ����o  �����  �x����      D  , ,  ������  �����o  �R���o  �R����  ������      D  , ,  �����  ����o  �����o  ������  �����      D  , ,  �X����  �X���o  �����o  ������  �X����      D  , ,  ������  �����o  �:���o  �:����  ������      D  , ,  ������  �����o  �~���o  �~����  ������      D  , ,  �@����  �@���o  �����o  ������  �@����      D  , ,  ������  �����o  ����o  �����  ������      D  , ,  ������  �����o  �r���o  �r����  ������      D  , ,  � ����  � ���o  �����o  ������  � ����      D  , ,  �x����  �x���o  ����o  �����  �x����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �R����  �R���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  ������  �����/  �:���/  �:����  ������      D  , ,  ������  �����/  �~���/  �~����  ������      D  , ,  �@����  �@���/  �����/  ������  �@����      D  , ,  ������  �����/  ����/  �����  ������      D  , ,  ������  �����/  �r���/  �r����  ������      D  , ,  � ����  � ���/  �����/  ������  � ����      D  , ,  �x����  �x���/  ����/  �����  �x����      D  , ,  ������  �����/  �R���/  �R����  ������      D  , ,  �����  ����/  �����/  ������  �����      D  , ,  �X����  �X���/  �����/  ������  �X����      D  , ,  ������  �����o  �:���o  �:����  ������      D  , ,  ������  �����o  �~���o  �~����  ������      D  , ,  �@����  �@���o  �����o  ������  �@����      D  , ,  ������  �����o  ����o  �����  ������      D  , ,  ������  �����o  �r���o  �r����  ������      D  , ,  �����Y  ������  �:����  �:���Y  �����Y      D  , ,  �����Y  ������  �~����  �~���Y  �����Y      D  , ,  �@���Y  �@����  ������  �����Y  �@���Y      D  , ,  �����Y  ������  �����  ����Y  �����Y      D  , ,  �����Y  ������  �r����  �r���Y  �����Y      D  , ,  � ���Y  � ����  ������  �����Y  � ���Y      D  , ,  �x���Y  �x����  �����  ����Y  �x���Y      D  , ,  �����Y  ������  �R����  �R���Y  �����Y      D  , ,  ����Y  �����  ������  �����Y  ����Y      D  , ,  �X���Y  �X����  ������  �����Y  �X���Y      D  , ,  ������  �����o  �R���o  �R����  ������      D  , ,  �����  ����o  �����o  ������  �����      D  , ,  �X����  �X���o  �����o  ������  �X����      D  , ,  �����  ������  �:����  �:���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �@���  �@����  ������  �����  �@���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �R����  �R���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  �����Y  ������  �:����  �:���Y  �����Y      D  , ,  �����Y  ������  �~����  �~���Y  �����Y      D  , ,  �@���Y  �@����  ������  �����Y  �@���Y      D  , ,  �����Y  ������  �����  ����Y  �����Y      D  , ,  �����Y  ������  �r����  �r���Y  �����Y      D  , ,  � ���Y  � ����  ������  �����Y  � ���Y      D  , ,  �x���Y  �x����  �����  ����Y  �x���Y      D  , ,  �����Y  ������  �R����  �R���Y  �����Y      D  , ,  ����Y  �����  ������  �����Y  ����Y      D  , ,  �X���Y  �X����  ������  �����Y  �X���Y      D  , ,  �����  ������  �:����  �:���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �@���  �@����  ������  �����  �@���      D  , ,  �����  ������  �����  ����  �����      D  , ,  ������  �����o  �.���o  �.����  ������      D  , ,  ������  �����o  �r���o  �r����  ������      D  , ,  �4����  �4���o  �����o  ������  �4����      D  , ,  �x����  �x���o  ����o  �����  �x����      D  , ,  ������  �����o  �f���o  �f����  ������      D  , ,  �����  ����o  �����o  ������  �����      D  , ,  �l����  �l���o  ����o  �����  �l����      D  , ,  ������  �����o  �F���o  �F����  ������      D  , ,  �����  ����o  �����o  ������  �����      D  , ,  �L����  �L���o  �����o  ������  �L����      D  , ,  �l����  �l���/  ����/  �����  �l����      D  , ,  ������  �����/  �F���/  �F����  ������      D  , ,  �����  ����/  �����/  ������  �����      D  , ,  �L����  �L���/  �����/  ������  �L����      D  , ,  �4���Y  �4����  ������  �����Y  �4���Y      D  , ,  �x���Y  �x����  �����  ����Y  �x���Y      D  , ,  �����Y  ������  �f����  �f���Y  �����Y      D  , ,  ����Y  �����  ������  �����Y  ����Y      D  , ,  �l���Y  �l����  �����  ����Y  �l���Y      D  , ,  �����Y  ������  �F����  �F���Y  �����Y      D  , ,  ����Y  �����  ������  �����Y  ����Y      D  , ,  �L���Y  �L����  ������  �����Y  �L���Y      D  , ,  ~@����  ~@���/  ~����/  ~�����  ~@����      D  , ,  ������  �����/  �.���/  �.����  ������      D  , ,  ������  �����/  �r���/  �r����  ������      D  , ,  �4���  �4����  ������  �����  �4���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �f����  �f���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �l���  �l����  �����  ����  �l���      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ~@����  ~@���o  ~����o  ~�����  ~@����      D  , ,  ������  �����o  �.���o  �.����  ������      D  , ,  ������  �����o  �r���o  �r����  ������      D  , ,  �4����  �4���o  �����o  ������  �4����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  �x����  �x���o  ����o  �����  �x����      D  , ,  ������  �����o  �f���o  �f����  ������      D  , ,  �����  ����o  �����o  ������  �����      D  , ,  �l����  �l���o  ����o  �����  �l����      D  , ,  ������  �����o  �F���o  �F����  ������      D  , ,  �����  ����o  �����o  ������  �����      D  , ,  �L����  �L���o  �����o  ������  �L����      D  , ,  �4����  �4���/  �����/  ������  �4����      D  , ,  �x����  �x���/  ����/  �����  �x����      D  , ,  ������  �����/  �f���/  �f����  ������      D  , ,  ����Y  �����  ������  �����Y  ����Y      D  , ,  �L���Y  �L����  ������  �����Y  �L���Y      D  , ,  �����  ����/  �����/  ������  �����      D  , ,  ����Y  �����  ������  �����Y  ����Y      D  , ,  �l���Y  �l����  �����  ����Y  �l���Y      D  , ,  �����Y  ������  �F����  �F���Y  �����Y      D  , ,  ~@���Y  ~@����  ~�����  ~����Y  ~@���Y      D  , ,  �����Y  ������  �.����  �.���Y  �����Y      D  , ,  �����Y  ������  �r����  �r���Y  �����Y      D  , ,  �4���Y  �4����  ������  �����Y  �4���Y      D  , ,  �x���Y  �x����  �����  ����Y  �x���Y      D  , ,  �����Y  ������  �f����  �f���Y  �����Y      D  , ,  ~@���Y  ~@����  ~�����  ~����Y  ~@���Y      D  , ,  �����Y  ������  �.����  �.���Y  �����Y      D  , ,  �����Y  ������  �r����  �r���Y  �����Y      D  , ,  ~@���  ~@����  ~�����  ~����  ~@���      D  , ,  �����  ������  �.����  �.���  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  �4���  �4����  ������  �����  �4���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �f����  �f���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �l���  �l����  �����  ����  �l���      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  ~@���  ~@����  ~�����  ~����  ~@���      D  , ,  �����  ������  �.����  �.���  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  ~@����  ~@���o  ~����o  ~�����  ~@����      D  , ,  ������  �����[  �r���[  �r����  ������      D  , ,  �4����  �4���[  �����[  ������  �4����      D  , ,  �x����  �x���[  ����[  �����  �x����      D  , ,  ������  �����[  �f���[  �f����  ������      D  , ,  �����  ����[  �����[  ������  �����      D  , ,  �l����  �l���[  ����[  �����  �l����      D  , ,  ������  �����[  �F���[  �F����  ������      D  , ,  �����  ����[  �����[  ������  �����      D  , ,  �L����  �L���[  �����[  ������  �L����      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  ~@���  ~@����  ~�����  ~����  ~@���      D  , ,  }���o  }���  }����  }����o  }���o      D  , ,  g���o  g���  ����  ����o  g���o      D  , ,  �����o  �����  �K���  �K���o  �����o      D  , ,  ����o  ����  �����  �����o  ����o      D  , ,  �Q���o  �Q���  �����  �����o  �Q���o      D  , ,  �����o  �����  �5���  �5���o  �����o      D  , ,  �����o  �����  �����  �����o  �����o      D  , ,  �;���o  �;���  �����  �����o  �;���o      D  , ,  �����o  �����  ����  ����o  �����o      D  , ,  ~@���  ~@����  ~�����  ~����  ~@���      D  , ,  �����  ������  �.����  �.���  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  �4���  �4����  ������  �����  �4���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �f����  �f���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �l���  �l����  �����  ����  �l���      D  , ,  �����  ������  �F����  �F���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �L���  �L����  ������  �����  �L���      D  , ,  �����o  �����  �m���  �m���o  �����o      D  , ,  �%���o  �%���  �����  �����o  �%���o      D  , ,  �����  ������  �.����  �.���  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  �4���  �4����  ������  �����  �4���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  ~@����  ~@���  ~����  ~�����  ~@����      D  , ,  ������  �����  �.���  �.����  ������      D  , ,  ������  �����  �r���  �r����  ������      D  , ,  �4����  �4���  �����  ������  �4����      D  , ,  �x����  �x���  ����  �����  �x����      D  , ,  ������  �����  �f���  �f����  ������      D  , ,  �����  ����  �����  ������  �����      D  , ,  �l����  �l���  ����  �����  �l����      D  , ,  ~@���E  ~@����  ~�����  ~����E  ~@���E      D  , ,  �����E  ������  �.����  �.���E  �����E      D  , ,  �����E  ������  �r����  �r���E  �����E      D  , ,  �4���E  �4����  ������  �����E  �4���E      D  , ,  �x���E  �x����  �����  ����E  �x���E      D  , ,  ~@����  ~@���[  ~����[  ~�����  ~@����      D  , ,  ������  �����[  �.���[  �.����  ������      D  , ,  ������  �����[  �r���[  �r����  ������      D  , ,  �4����  �4���[  �����[  ������  �4����      D  , ,  �x����  �x���[  ����[  �����  �x����      D  , ,  ������  �����[  �f���[  �f����  ������      D  , ,  �����  ����[  �����[  ������  �����      D  , ,  �l����  �l���[  ����[  �����  �l����      D  , ,  ������  �����[  �F���[  �F����  ������      D  , ,  �����  ����[  �����[  ������  �����      D  , ,  �L����  �L���[  �����[  ������  �L����      D  , ,  �����E  ������  �f����  �f���E  �����E      D  , ,  ����E  �����  ������  �����E  ����E      D  , ,  �l���E  �l����  �����  ����E  �l���E      D  , ,  �����E  ������  �F����  �F���E  �����E      D  , ,  ����E  �����  ������  �����E  ����E      D  , ,  �L���E  �L����  ������  �����E  �L���E      D  , ,  ������  �����  �F���  �F����  ������      D  , ,  �����  ����  �����  ������  �����      D  , ,  �L����  �L���  �����  ������  �L����      D  , ,  �����  ������  �f����  �f���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  }���/  }����  }�����  }����/  }���/      D  , ,  g���/  g����  �����  ����/  g���/      D  , ,  �����/  ������  �K����  �K���/  �����/      D  , ,  ����/  �����  ������  �����/  ����/      D  , ,  �Q���/  �Q����  ������  �����/  �Q���/      D  , ,  �����/  ������  �5����  �5���/  �����/      D  , ,  �����/  ������  ������  �����/  �����/      D  , ,  �;���/  �;����  ������  �����/  �;���/      D  , ,  �����/  ������  �����  ����/  �����/      D  , ,  �����/  ������  �m����  �m���/  �����/      D  , ,  �%���/  �%����  ������  �����/  �%���/      D  , ,  �l���  �l����  �����  ����  �l���      D  , ,  ~@����  ~@���[  ~����[  ~�����  ~@����      D  , ,  ������  �����[  �.���[  �.����  ������      D  , ,  �]���o  �]���  �����  �����o  �]���o      D  , ,  �����o  �����  �A���  �A���o  �����o      D  , ,  �����o  �����  �����  �����o  �����o      D  , ,  �G���o  �G���  �����  �����o  �G���o      D  , ,  �����o  �����  �+���  �+���o  �����o      D  , ,  �����o  �����  �y���  �y���o  �����o      D  , ,  �1���o  �1���  �����  �����o  �1���o      D  , ,  ����o  ����  ����  ����o  ����o      D  , ,  � ����  � ���[  �����[  ������  � ����      D  , ,  �x����  �x���[  ����[  �����  �x����      D  , ,  ������  �����[  �R���[  �R����  ������      D  , ,  �����  ����[  �����[  ������  �����      D  , ,  �X����  �X���[  �����[  ������  �X����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  ������  �����  �:���  �:����  ������      D  , ,  ������  �����  �~���  �~����  ������      D  , ,  �@����  �@���  �����  ������  �@����      D  , ,  ������  �����  ����  �����  ������      D  , ,  ������  �����  �r���  �r����  ������      D  , ,  � ����  � ���  �����  ������  � ����      D  , ,  �x����  �x���  ����  �����  �x����      D  , ,  ������  �����  �R���  �R����  ������      D  , ,  �����  ����  �����  ������  �����      D  , ,  �X����  �X���  �����  ������  �X����      D  , ,  �@���  �@����  ������  �����  �@���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �R����  �R���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  �����  ������  �:����  �:���  �����      D  , ,  ������  �����[  �:���[  �:����  ������      D  , ,  ������  �����[  �~���[  �~����  ������      D  , ,  �����E  ������  �:����  �:���E  �����E      D  , ,  ������  �����[  �:���[  �:����  ������      D  , ,  ������  �����[  �~���[  �~����  ������      D  , ,  �@����  �@���[  �����[  ������  �@����      D  , ,  ������  �����[  ����[  �����  ������      D  , ,  ������  �����[  �r���[  �r����  ������      D  , ,  � ����  � ���[  �����[  ������  � ����      D  , ,  �x����  �x���[  ����[  �����  �x����      D  , ,  ������  �����[  �R���[  �R����  ������      D  , ,  �����  ����[  �����[  ������  �����      D  , ,  �X����  �X���[  �����[  ������  �X����      D  , ,  �����E  ������  �~����  �~���E  �����E      D  , ,  �@���E  �@����  ������  �����E  �@���E      D  , ,  �����E  ������  �����  ����E  �����E      D  , ,  �����E  ������  �r����  �r���E  �����E      D  , ,  � ���E  � ����  ������  �����E  � ���E      D  , ,  �x���E  �x����  �����  ����E  �x���E      D  , ,  �����E  ������  �R����  �R���E  �����E      D  , ,  ����E  �����  ������  �����E  ����E      D  , ,  �X���E  �X����  ������  �����E  �X���E      D  , ,  �@����  �@���[  �����[  ������  �@����      D  , ,  �����  ������  �:����  �:���  �����      D  , ,  �����  ������  �~����  �~���  �����      D  , ,  �@���  �@����  ������  �����  �@���      D  , ,  �����  ������  �����  ����  �����      D  , ,  �����  ������  �r����  �r���  �����      D  , ,  � ���  � ����  ������  �����  � ���      D  , ,  �x���  �x����  �����  ����  �x���      D  , ,  �����  ������  �R����  �R���  �����      D  , ,  ����  �����  ������  �����  ����      D  , ,  �X���  �X����  ������  �����  �X���      D  , ,  ������  �����[  ����[  �����  ������      D  , ,  ������  �����[  �r���[  �r����  ������      D  , ,  �s���/  �s����  �	����  �	���/  �s���/      D  , ,  �����/  ������  �W����  �W���/  �����/      D  , ,  ����/  �����  ������  �����/  ����/      D  , ,  �]���/  �]����  ������  �����/  �]���/      D  , ,  �����/  ������  �A����  �A���/  �����/      D  , ,  �����/  ������  ������  �����/  �����/      D  , ,  �G���/  �G����  ������  �����/  �G���/      D  , ,  �����/  ������  �+����  �+���/  �����/      D  , ,  �����/  ������  �y����  �y���/  �����/      D  , ,  �1���/  �1����  ������  �����/  �1���/      D  , ,  ����/  �����  �����  ����/  ����/      D  , ,  �s���o  �s���  �	���  �	���o  �s���o      D  , ,  �����o  �����  �W���  �W���o  �����o      D  , ,  ����o  ����  �����  �����o  ����o      D  , ,  ������  �����  �:���  �:����  ������      D  , ,  ������  �����  �~���  �~����  ������      D  , ,  �@����  �@���  �����  ������  �@����      D  , ,  ������  �����  ����  �����  ������      D  , ,  ������  �����  �r���  �r����  ������      D  , ,  � ����  � ���  �����  ������  � ����      D  , ,  �x����  �x���  ����  �����  �x����      D  , ,  ������  �����  �R���  �R����  ������      D  , ,  �����  ����  �����  ������  �����      D  , ,  �X����  �X���  �����  ������  �X����      D  , ,  �����E  ������  �:����  �:���E  �����E      D  , ,  �����E  ������  �~����  �~���E  �����E      D  , ,  �@���E  �@����  ������  �����E  �@���E      D  , ,  �����E  ������  �����  ����E  �����E      D  , ,  �����E  ������  �r����  �r���E  �����E      D  , ,  � ���E  � ����  ������  �����E  � ���E      D  , ,  �x���E  �x����  �����  ����E  �x���E      D  , ,  �����E  ������  �R����  �R���E  �����E      D  , ,  ����E  �����  ������  �����E  ����E      D  , ,  �X���E  �X����  ������  �����E  �X���E      D  , ,  �����  �����I  �~���I  �~���  �����      D  , ,  �����  �����I  ����I  ����  �����      D  , ,  � ���  � ���I  �����I  �����  � ���      D  , ,  �����  �����I  �R���I  �R���  �����      D  , ,  �X���  �X���I  �����I  �����  �X���      D  , ,  ����~s  ����	  �~��	  �~��~s  ����~s      D  , ,  ����~s  ����	  ���	  ���~s  ����~s      D  , ,  � ��~s  � ��	  ����	  ����~s  � ��~s      D  , ,  ����~s  ����	  �R��	  �R��~s  ����~s      D  , ,  �X��~s  �X��	  ����	  ����~s  �X��~s      D  , ,  ����}3  ����}�  �~��}�  �~��}3  ����}3      D  , ,  ����}3  ����}�  ���}�  ���}3  ����}3      D  , ,  � ��}3  � ��}�  ����}�  ����}3  � ��}3      D  , ,  ����}3  ����}�  �R��}�  �R��}3  ����}3      D  , ,  �X��}3  �X��}�  ����}�  ����}3  �X��}3      D  , ,  ����{�  ����|�  �~��|�  �~��{�  ����{�      D  , ,  ����{�  ����|�  ���|�  ���{�  ����{�      D  , ,  � ��{�  � ��|�  ����|�  ����{�  � ��{�      D  , ,  ����{�  ����|�  �R��|�  �R��{�  ����{�      D  , ,  �X��{�  �X��|�  ����|�  ����{�  �X��{�      D  , ,  �����  �����I  �F���I  �F���  �����      D  , ,  �L���  �L���I  �����I  �����  �L���      D  , ,  �����E  ������  �f����  �f���E  �����E      D  , ,  ����E  �����  ������  �����E  ����E      D  , ,  �l���E  �l����  �����  ����E  �l���E      D  , ,  �����E  ������  �F����  �F���E  �����E      D  , ,  ����E  �����  ������  �����E  ����E      D  , ,  ~@��~s  ~@��	  ~���	  ~���~s  ~@��~s      D  , ,  ����~s  ����	  �r��	  �r��~s  ����~s      D  , ,  �x��~s  �x��	  ���	  ���~s  �x��~s      D  , ,  ���~s  ���	  ����	  ����~s  ���~s      D  , ,  ����~s  ����	  �F��	  �F��~s  ����~s      D  , ,  �L��~s  �L��	  ����	  ����~s  �L��~s      D  , ,  �L���E  �L����  ������  �����E  �L���E      D  , ,  �����  ����  �����  ������  �����      D  , ,  �l����  �l���  ����  �����  �l����      D  , ,  ������  �����  �F���  �F����  ������      D  , ,  �����  ����  �����  ������  �����      D  , ,  ~@��}3  ~@��}�  ~���}�  ~���}3  ~@��}3      D  , ,  ����}3  ����}�  �r��}�  �r��}3  ����}3      D  , ,  �x��}3  �x��}�  ���}�  ���}3  �x��}3      D  , ,  ���}3  ���}�  ����}�  ����}3  ���}3      D  , ,  ����}3  ����}�  �F��}�  �F��}3  ����}3      D  , ,  �L��}3  �L��}�  ����}�  ����}3  �L��}3      D  , ,  �L����  �L���  �����  ������  �L����      D  , ,  ~@���E  ~@����  ~�����  ~����E  ~@���E      D  , ,  �����E  ������  �.����  �.���E  �����E      D  , ,  �����E  ������  �r����  �r���E  �����E      D  , ,  �4���E  �4����  ������  �����E  �4���E      D  , ,  ~@��{�  ~@��|�  ~���|�  ~���{�  ~@��{�      D  , ,  ����{�  ����|�  �r��|�  �r��{�  ����{�      D  , ,  �x��{�  �x��|�  ���|�  ���{�  �x��{�      D  , ,  ���{�  ���|�  ����|�  ����{�  ���{�      D  , ,  ����{�  ����|�  �F��|�  �F��{�  ����{�      D  , ,  �L��{�  �L��|�  ����|�  ����{�  �L��{�      D  , ,  �x���E  �x����  �����  ����E  �x���E      D  , ,  ~@���  ~@���I  ~����I  ~����  ~@���      D  , ,  �����  �����I  �r���I  �r���  �����      D  , ,  �x���  �x���I  ����I  ����  �x���      D  , ,  ����  ����I  �����I  �����  ����      D  , ,  ~@����  ~@���  ~����  ~�����  ~@����      D  , ,  ������  �����  �.���  �.����  ������      D  , ,  ������  �����  �r���  �r����  ������      D  , ,  �4����  �4���  �����  ������  �4����      D  , ,  �x����  �x���  ����  �����  �x����      D  , ,  ������  �����  �f���  �f����  ������      D  , ,  �(��q�  �(��r   ����r   ����q�  �(��q�      D  , ,  �v��q�  �v��r   ���r   ���q�  �v��q�      D  , ,  ����q�  ����r   �Z��r   �Z��q�  ����q�      D  , ,  ���q�  ���r   ����r   ����q�  ���q�      D  , ,  �`��q�  �`��r   ����r   ����q�  �`��q�      D  , ,  ~T��pJ  ~T��p�  ~���p�  ~���pJ  ~T��pJ      D  , ,  ����pJ  ����p�  �8��p�  �8��pJ  ����pJ      D  , ,  ����pJ  ����p�  ����p�  ����pJ  ����pJ      D  , ,  �>��pJ  �>��p�  ����p�  ����pJ  �>��pJ      D  , ,  ����pJ  ����p�  �"��p�  �"��pJ  ����pJ      D  , ,  ����pJ  ����p�  �p��p�  �p��pJ  ����pJ      D  , ,  �(��pJ  �(��p�  ����p�  ����pJ  �(��pJ      D  , ,  �v��pJ  �v��p�  ���p�  ���pJ  �v��pJ      D  , ,  ����pJ  ����p�  �Z��p�  �Z��pJ  ����pJ      D  , ,  ���pJ  ���p�  ����p�  ����pJ  ���pJ      D  , ,  �`��pJ  �`��p�  ����p�  ����pJ  �`��pJ      D  , ,  ~T��o
  ~T��o�  ~���o�  ~���o
  ~T��o
      D  , ,  ����o
  ����o�  �8��o�  �8��o
  ����o
      D  , ,  ����o
  ����o�  ����o�  ����o
  ����o
      D  , ,  �>��o
  �>��o�  ����o�  ����o
  �>��o
      D  , ,  ����o
  ����o�  �"��o�  �"��o
  ����o
      D  , ,  ����o
  ����o�  �p��o�  �p��o
  ����o
      D  , ,  �(��o
  �(��o�  ����o�  ����o
  �(��o
      D  , ,  �v��o
  �v��o�  ���o�  ���o
  �v��o
      D  , ,  ����o
  ����o�  �Z��o�  �Z��o
  ����o
      D  , ,  ���o
  ���o�  ����o�  ����o
  ���o
      D  , ,  �`��o
  �`��o�  ����o�  ����o
  �`��o
      D  , ,  ~T��m�  ~T��n`  ~���n`  ~���m�  ~T��m�      D  , ,  ����m�  ����n`  �8��n`  �8��m�  ����m�      D  , ,  ����m�  ����n`  ����n`  ����m�  ����m�      D  , ,  �>��m�  �>��n`  ����n`  ����m�  �>��m�      D  , ,  ����m�  ����n`  �"��n`  �"��m�  ����m�      D  , ,  ����m�  ����n`  �p��n`  �p��m�  ����m�      D  , ,  �(��m�  �(��n`  ����n`  ����m�  �(��m�      D  , ,  �v��m�  �v��n`  ���n`  ���m�  �v��m�      D  , ,  ����m�  ����n`  �Z��n`  �Z��m�  ����m�      D  , ,  ���m�  ���n`  ����n`  ����m�  ���m�      D  , ,  �`��m�  �`��n`  ����n`  ����m�  �`��m�      D  , ,  ~T��l�  ~T��m   ~���m   ~���l�  ~T��l�      D  , ,  ����l�  ����m   �8��m   �8��l�  ����l�      D  , ,  ����l�  ����m   ����m   ����l�  ����l�      D  , ,  �>��l�  �>��m   ����m   ����l�  �>��l�      D  , ,  ����l�  ����m   �"��m   �"��l�  ����l�      D  , ,  ����l�  ����m   �p��m   �p��l�  ����l�      D  , ,  �(��l�  �(��m   ����m   ����l�  �(��l�      D  , ,  �v��l�  �v��m   ���m   ���l�  �v��l�      D  , ,  ����l�  ����m   �Z��m   �Z��l�  ����l�      D  , ,  ���l�  ���m   ����m   ����l�  ���l�      D  , ,  �`��l�  �`��m   ����m   ����l�  �`��l�      D  , ,  ~T��kJ  ~T��k�  ~���k�  ~���kJ  ~T��kJ      D  , ,  ����kJ  ����k�  �8��k�  �8��kJ  ����kJ      D  , ,  ����kJ  ����k�  ����k�  ����kJ  ����kJ      D  , ,  �>��kJ  �>��k�  ����k�  ����kJ  �>��kJ      D  , ,  ����kJ  ����k�  �"��k�  �"��kJ  ����kJ      D  , ,  ����kJ  ����k�  �p��k�  �p��kJ  ����kJ      D  , ,  �(��kJ  �(��k�  ����k�  ����kJ  �(��kJ      D  , ,  �v��kJ  �v��k�  ���k�  ���kJ  �v��kJ      D  , ,  ����kJ  ����k�  �Z��k�  �Z��kJ  ����kJ      D  , ,  ���kJ  ���k�  ����k�  ����kJ  ���kJ      D  , ,  �`��kJ  �`��k�  ����k�  ����kJ  �`��kJ      D  , ,  ~T��j
  ~T��j�  ~���j�  ~���j
  ~T��j
      D  , ,  ����j
  ����j�  �8��j�  �8��j
  ����j
      D  , ,  ����j
  ����j�  ����j�  ����j
  ����j
      D  , ,  �>��j
  �>��j�  ����j�  ����j
  �>��j
      D  , ,  ����j
  ����j�  �"��j�  �"��j
  ����j
      D  , ,  ����j
  ����j�  �p��j�  �p��j
  ����j
      D  , ,  �(��j
  �(��j�  ����j�  ����j
  �(��j
      D  , ,  �v��j
  �v��j�  ���j�  ���j
  �v��j
      D  , ,  ����j
  ����j�  �Z��j�  �Z��j
  ����j
      D  , ,  ���j
  ���j�  ����j�  ����j
  ���j
      D  , ,  �`��j
  �`��j�  ����j�  ����j
  �`��j
      D  , ,  ~T��q�  ~T��r   ~���r   ~���q�  ~T��q�      D  , ,  ����q�  ����r   �8��r   �8��q�  ����q�      D  , ,  ����q�  ����r   ����r   ����q�  ����q�      D  , ,  �>��q�  �>��r   ����r   ����q�  �>��q�      D  , ,  ����q�  ����r   �"��r   �"��q�  ����q�      D  , ,  ����q�  ����r   �p��r   �p��q�  ����q�      D  , ,  ����q�  ����r   �j��r   �j��q�  ����q�      D  , ,  �"��q�  �"��r   ����r   ����q�  �"��q�      D  , ,  ����pJ  ����p�  �j��p�  �j��pJ  ����pJ      D  , ,  �"��pJ  �"��p�  ����p�  ����pJ  �"��pJ      D  , ,  ����o
  ����o�  �j��o�  �j��o
  ����o
      D  , ,  �"��o
  �"��o�  ����o�  ����o
  �"��o
      D  , ,  �p��o
  �p��o�  ���o�  ���o
  �p��o
      D  , ,  ����o
  ����o�  �T��o�  �T��o
  ����o
      D  , ,  ����l�  ����m   �j��m   �j��l�  ����l�      D  , ,  �"��l�  �"��m   ����m   ����l�  �"��l�      D  , ,  �p��l�  �p��m   ���m   ���l�  �p��l�      D  , ,  ����l�  ����m   �T��m   �T��l�  ����l�      D  , ,  ���l�  ���m   ����m   ����l�  ���l�      D  , ,  �Z��l�  �Z��m   ����m   ����l�  �Z��l�      D  , ,  ����l�  ����m   �>��m   �>��l�  ����l�      D  , ,  ����l�  ����m   ����m   ����l�  ����l�      D  , ,  �D��l�  �D��m   ����m   ����l�  �D��l�      D  , ,  ���o
  ���o�  ����o�  ����o
  ���o
      D  , ,  �Z��o
  �Z��o�  ����o�  ����o
  �Z��o
      D  , ,  ����o
  ����o�  �>��o�  �>��o
  ����o
      D  , ,  ����o
  ����o�  ����o�  ����o
  ����o
      D  , ,  �D��o
  �D��o�  ����o�  ����o
  �D��o
      D  , ,  �p��pJ  �p��p�  ���p�  ���pJ  �p��pJ      D  , ,  ����pJ  ����p�  �T��p�  �T��pJ  ����pJ      D  , ,  ���pJ  ���p�  ����p�  ����pJ  ���pJ      D  , ,  �Z��pJ  �Z��p�  ����p�  ����pJ  �Z��pJ      D  , ,  ����pJ  ����p�  �>��p�  �>��pJ  ����pJ      D  , ,  ����pJ  ����p�  ����p�  ����pJ  ����pJ      D  , ,  ����kJ  ����k�  �j��k�  �j��kJ  ����kJ      D  , ,  �"��kJ  �"��k�  ����k�  ����kJ  �"��kJ      D  , ,  �p��kJ  �p��k�  ���k�  ���kJ  �p��kJ      D  , ,  ����kJ  ����k�  �T��k�  �T��kJ  ����kJ      D  , ,  ���kJ  ���k�  ����k�  ����kJ  ���kJ      D  , ,  �Z��kJ  �Z��k�  ����k�  ����kJ  �Z��kJ      D  , ,  ����kJ  ����k�  �>��k�  �>��kJ  ����kJ      D  , ,  ����kJ  ����k�  ����k�  ����kJ  ����kJ      D  , ,  �D��kJ  �D��k�  ����k�  ����kJ  �D��kJ      D  , ,  �D��pJ  �D��p�  ����p�  ����pJ  �D��pJ      D  , ,  �p��q�  �p��r   ���r   ���q�  �p��q�      D  , ,  ����q�  ����r   �T��r   �T��q�  ����q�      D  , ,  ���q�  ���r   ����r   ����q�  ���q�      D  , ,  �Z��q�  �Z��r   ����r   ����q�  �Z��q�      D  , ,  ����m�  ����n`  �j��n`  �j��m�  ����m�      D  , ,  �"��m�  �"��n`  ����n`  ����m�  �"��m�      D  , ,  �p��m�  �p��n`  ���n`  ���m�  �p��m�      D  , ,  ����m�  ����n`  �T��n`  �T��m�  ����m�      D  , ,  ���m�  ���n`  ����n`  ����m�  ���m�      D  , ,  �Z��m�  �Z��n`  ����n`  ����m�  �Z��m�      D  , ,  ����j
  ����j�  �j��j�  �j��j
  ����j
      D  , ,  �"��j
  �"��j�  ����j�  ����j
  �"��j
      D  , ,  �p��j
  �p��j�  ���j�  ���j
  �p��j
      D  , ,  ����j
  ����j�  �T��j�  �T��j
  ����j
      D  , ,  ���j
  ���j�  ����j�  ����j
  ���j
      D  , ,  �Z��j
  �Z��j�  ����j�  ����j
  �Z��j
      D  , ,  ����j
  ����j�  �>��j�  �>��j
  ����j
      D  , ,  ����j
  ����j�  ����j�  ����j
  ����j
      D  , ,  �D��j
  �D��j�  ����j�  ����j
  �D��j
      D  , ,  ����m�  ����n`  �>��n`  �>��m�  ����m�      D  , ,  ����m�  ����n`  ����n`  ����m�  ����m�      D  , ,  �D��m�  �D��n`  ����n`  ����m�  �D��m�      D  , ,  ����q�  ����r   �>��r   �>��q�  ����q�      D  , ,  ����q�  ����r   ����r   ����q�  ����q�      D  , ,  �D��q�  �D��r   ����r   ����q�  �D��q�      D  , ,  g4���E  g4����  g�����  g����E  g4���E      D  , ,  g4���  g4���I  g����I  g����  g4���      D  , ,  k����  k����I  lf���I  lf���  k����      D  , ,  pl���  pl���I  q���I  q���  pl���      D  , ,  u���  u���I  u����I  u����  u���      D  , ,  g4��}3  g4��}�  g���}�  g���}3  g4��}3      D  , ,  k���}3  k���}�  lf��}�  lf��}3  k���}3      D  , ,  pl��}3  pl��}�  q��}�  q��}3  pl��}3      D  , ,  u��}3  u��}�  u���}�  u���}3  u��}3      D  , ,  y���}3  y���}�  z:��}�  z:��}3  y���}3      D  , ,  i�����  i����  j"���  j"����  i�����      D  , ,  y����  y����I  z:���I  z:���  y����      D  , ,  i����E  i�����  j"����  j"���E  i����E      D  , ,  k����E  k�����  lf����  lf���E  k����E      D  , ,  n(���E  n(����  n�����  n����E  n(���E      D  , ,  pl���E  pl����  q����  q���E  pl���E      D  , ,  r����E  r�����  sZ����  sZ���E  r����E      D  , ,  u���E  u����  u�����  u����E  u���E      D  , ,  w`���E  w`����  w�����  w����E  w`���E      D  , ,  y����E  y�����  z:����  z:���E  y����E      D  , ,  {����E  {�����  |�����  |����E  {����E      D  , ,  g4��{�  g4��|�  g���|�  g���{�  g4��{�      D  , ,  k�����  k����  lf���  lf����  k�����      D  , ,  k���{�  k���|�  lf��|�  lf��{�  k���{�      D  , ,  pl��{�  pl��|�  q��|�  q��{�  pl��{�      D  , ,  u��{�  u��|�  u���|�  u���{�  u��{�      D  , ,  y���{�  y���|�  z:��|�  z:��{�  y���{�      D  , ,  g4��~s  g4��	  g���	  g���~s  g4��~s      D  , ,  k���~s  k���	  lf��	  lf��~s  k���~s      D  , ,  pl��~s  pl��	  q��	  q��~s  pl��~s      D  , ,  u��~s  u��	  u���	  u���~s  u��~s      D  , ,  d�����  d����  e����  e�����  d�����      D  , ,  y���~s  y���	  z:��	  z:��~s  y���~s      D  , ,  n(����  n(���  n����  n�����  n(����      D  , ,  d����E  d�����  e�����  e����E  d����E      D  , ,  g4����  g4���  g����  g�����  g4����      D  , ,  pl����  pl���  q���  q����  pl����      D  , ,  r�����  r����  sZ���  sZ����  r�����      D  , ,  u����  u���  u����  u�����  u����      D  , ,  w`����  w`���  w����  w�����  w`����      D  , ,  y�����  y����  z:���  z:����  y�����      D  , ,  {�����  {����  |����  |�����  {�����      D  , ,  b�����  b����  c.���  c.����  b�����      D  , ,  b����  b����I  c.���I  c.���  b����      D  , ,  `T����  `T���  `����  `�����  `T����      D  , ,  `T���E  `T����  `�����  `����E  `T���E      D  , ,  b����E  b�����  c.����  c.���E  b����E      D  , ,  ]���}3  ]���}�  ^���}�  ^���}3  ]���}3      D  , ,  b���}3  b���}�  c.��}�  c.��}3  b���}3      D  , ,  J���y�  J���zT  K���zT  K���y�  J���y�      D  , ,  N���y�  N���zT  O[��zT  O[��y�  N���y�      D  , ,  J���x~  J���y  K���y  K���x~  J���x~      D  , ,  N���x~  N���y  O[��y  O[��x~  N���x~      D  , ,  ]����  ]����I  ^����I  ^����  ]����      D  , ,  ]����E  ]�����  ^�����  ^����E  ]����E      D  , ,  ]���~s  ]���	  ^���	  ^���~s  ]���~s      D  , ,  b���~s  b���	  c.��	  c.��~s  b���~s      D  , ,  ]�����  ]����  ^����  ^�����  ]�����      D  , ,  ]���{�  ]���|�  ^���|�  ^���{�  ]���{�      D  , ,  b���{�  b���|�  c.��|�  c.��{�  b���{�      D  , ,  N���s~  N���t  O[��t  O[��s~  N���s~      D  , ,  J���r>  J���r�  K���r�  K���r>  J���r>      D  , ,  N���r>  N���r�  O[��r�  O[��r>  N���r>      D  , ,  J���p�  J���q�  K���q�  K���p�  J���p�      D  , ,  N���p�  N���q�  O[��q�  O[��p�  N���p�      D  , ,  J���w>  J���w�  K���w�  K���w>  J���w>      D  , ,  N���w>  N���w�  O[��w�  O[��w>  N���w>      D  , ,  J���u�  J���v�  K���v�  K���u�  J���u�      D  , ,  N���u�  N���v�  O[��v�  O[��u�  N���u�      D  , ,  J���t�  J���uT  K���uT  K���t�  J���t�      D  , ,  N���t�  N���uT  O[��uT  O[��t�  N���t�      D  , ,  J���s~  J���t  K���t  K���s~  J���s~      D  , ,  wj��j
  wj��j�  x ��j�  x ��j
  wj��j
      D  , ,  y���j
  y���j�  zN��j�  zN��j
  y���j
      D  , ,  |��j
  |��j�  |���j�  |���j
  |��j
      D  , ,  |��kJ  |��k�  |���k�  |���kJ  |��kJ      D  , ,  y���pJ  y���p�  zN��p�  zN��pJ  y���pJ      D  , ,  |��pJ  |��p�  |���p�  |���pJ  |��pJ      D  , ,  |��l�  |��m   |���m   |���l�  |��l�      D  , ,  y���q�  y���r   zN��r   zN��q�  y���q�      D  , ,  |��q�  |��r   |���r   |���q�  |��q�      D  , ,  r���l�  r���m   sd��m   sd��l�  r���l�      D  , ,  u��l�  u��m   u���m   u���l�  u��l�      D  , ,  wj��l�  wj��m   x ��m   x ��l�  wj��l�      D  , ,  y���l�  y���m   zN��m   zN��l�  y���l�      D  , ,  r���pJ  r���p�  sd��p�  sd��pJ  r���pJ      D  , ,  u��pJ  u��p�  u���p�  u���pJ  u��pJ      D  , ,  wj��pJ  wj��p�  x ��p�  x ��pJ  wj��pJ      D  , ,  r���o
  r���o�  sd��o�  sd��o
  r���o
      D  , ,  u��o
  u��o�  u���o�  u���o
  u��o
      D  , ,  wj��o
  wj��o�  x ��o�  x ��o
  wj��o
      D  , ,  y���o
  y���o�  zN��o�  zN��o
  y���o
      D  , ,  |��o
  |��o�  |���o�  |���o
  |��o
      D  , ,  r���m�  r���n`  sd��n`  sd��m�  r���m�      D  , ,  u��m�  u��n`  u���n`  u���m�  u��m�      D  , ,  r���kJ  r���k�  sd��k�  sd��kJ  r���kJ      D  , ,  u��kJ  u��k�  u���k�  u���kJ  u��kJ      D  , ,  wj��kJ  wj��k�  x ��k�  x ��kJ  wj��kJ      D  , ,  y���kJ  y���k�  zN��k�  zN��kJ  y���kJ      D  , ,  r���j
  r���j�  sd��j�  sd��j
  r���j
      D  , ,  u��j
  u��j�  u���j�  u���j
  u��j
      D  , ,  wj��m�  wj��n`  x ��n`  x ��m�  wj��m�      D  , ,  y���m�  y���n`  zN��n`  zN��m�  y���m�      D  , ,  |��m�  |��n`  |���n`  |���m�  |��m�      D  , ,  r���q�  r���r   sd��r   sd��q�  r���q�      D  , ,  u��q�  u��r   u���r   u���q�  u��q�      D  , ,  wj��q�  wj��r   x ��r   x ��q�  wj��q�      D  , ,  vC��d�  vC��e#  v���e#  v���d�  vC��d�      D  , ,  x���d�  x���e#  y'��e#  y'��d�  x���d�      D  , ,  z���d�  z���e#  {u��e#  {u��d�  z���d�      D  , ,  r���a�  r���b&  sd��b&  sd��a�  r���a�      D  , ,  u��a�  u��b&  u���b&  u���a�  u��a�      D  , ,  wj��a�  wj��b&  x ��b&  x ��a�  wj��a�      D  , ,  y���a�  y���b&  zN��b&  zN��a�  y���a�      D  , ,  |��a�  |��b&  |���b&  |���a�  |��a�      D  , ,  u��h�  u��i`  u���i`  u���h�  u��h�      D  , ,  r���`P  r���`�  sd��`�  sd��`P  r���`P      D  , ,  u��`P  u��`�  u���`�  u���`P  u��`P      D  , ,  wj��`P  wj��`�  x ��`�  x ��`P  wj��`P      D  , ,  y���`P  y���`�  zN��`�  zN��`P  y���`P      D  , ,  |��`P  |��`�  |���`�  |���`P  |��`P      D  , ,  wj��h�  wj��i`  x ��i`  x ��h�  wj��h�      D  , ,  y���h�  y���i`  zN��i`  zN��h�  y���h�      D  , ,  r���_  r���_�  sd��_�  sd��_  r���_      D  , ,  u��_  u��_�  u���_�  u���_  u��_      D  , ,  wj��_  wj��_�  x ��_�  x ��_  wj��_      D  , ,  y���_  y���_�  zN��_�  zN��_  y���_      D  , ,  |��_  |��_�  |���_�  |���_  |��_      D  , ,  |��h�  |��i`  |���i`  |���h�  |��h�      D  , ,  r���h�  r���i`  sd��i`  sd��h�  r���h�      D  , ,  r���]�  r���^f  sd��^f  sd��]�  r���]�      D  , ,  u��]�  u��^f  u���^f  u���]�  u��]�      D  , ,  wj��]�  wj��^f  x ��^f  x ��]�  wj��]�      D  , ,  y���]�  y���^f  zN��^f  zN��]�  y���]�      D  , ,  |��]�  |��^f  |���^f  |���]�  |��]�      D  , ,  s���e�  s���fc  t���fc  t���e�  s���e�      D  , ,  r���\�  r���]&  sd��]&  sd��\�  r���\�      D  , ,  u��\�  u��]&  u���]&  u���\�  u��\�      D  , ,  wj��\�  wj��]&  x ��]&  x ��\�  wj��\�      D  , ,  y���\�  y���]&  zN��]&  zN��\�  y���\�      D  , ,  |��\�  |��]&  |���]&  |���\�  |��\�      D  , ,  vC��e�  vC��fc  v���fc  v���e�  vC��e�      D  , ,  r���[P  r���[�  sd��[�  sd��[P  r���[P      D  , ,  u��[P  u��[�  u���[�  u���[P  u��[P      D  , ,  wj��[P  wj��[�  x ��[�  x ��[P  wj��[P      D  , ,  y���[P  y���[�  zN��[�  zN��[P  y���[P      D  , ,  |��[P  |��[�  |���[�  |���[P  |��[P      D  , ,  x���e�  x���fc  y'��fc  y'��e�  x���e�      D  , ,  r���Z  r���Z�  sd��Z�  sd��Z  r���Z      D  , ,  u��Z  u��Z�  u���Z�  u���Z  u��Z      D  , ,  wj��Z  wj��Z�  x ��Z�  x ��Z  wj��Z      D  , ,  y���Z  y���Z�  zN��Z�  zN��Z  y���Z      D  , ,  |��Z  |��Z�  |���Z�  |���Z  |��Z      D  , ,  z���e�  z���fc  {u��fc  {u��e�  z���e�      D  , ,  r���X�  r���Yf  sd��Yf  sd��X�  r���X�      D  , ,  u��X�  u��Yf  u���Yf  u���X�  u��X�      D  , ,  wj��X�  wj��Yf  x ��Yf  x ��X�  wj��X�      D  , ,  y���X�  y���Yf  zN��Yf  zN��X�  y���X�      D  , ,  |��X�  |��Yf  |���Yf  |���X�  |��X�      D  , ,  s���d�  s���e#  t���e#  t���d�  s���d�      D  , ,  ����d�  ����e#  ����e#  ����d�  ����d�      D  , ,  �I��d�  �I��e#  ����e#  ����d�  �I��d�      D  , ,  ����d�  ����e#  �-��e#  �-��d�  ����d�      D  , ,  ����d�  ����e#  �{��e#  �{��d�  ����d�      D  , ,  �3��d�  �3��e#  ����e#  ����d�  �3��d�      D  , ,  ����d�  ����e#  ���e#  ���d�  ����d�      D  , ,  ����d�  ����e#  �e��e#  �e��d�  ����d�      D  , ,  ���d�  ���e#  ����e#  ����d�  ���d�      D  , ,  �k��d�  �k��e#  ���e#  ���d�  �k��d�      D  , ,  ����h�  ����i`  �j��i`  �j��h�  ����h�      D  , ,  �"��h�  �"��i`  ����i`  ����h�  �"��h�      D  , ,  �p��h�  �p��i`  ���i`  ���h�  �p��h�      D  , ,  ����a�  ����b&  �j��b&  �j��a�  ����a�      D  , ,  �"��a�  �"��b&  ����b&  ����a�  �"��a�      D  , ,  �p��a�  �p��b&  ���b&  ���a�  �p��a�      D  , ,  ����a�  ����b&  �T��b&  �T��a�  ����a�      D  , ,  ���a�  ���b&  ����b&  ����a�  ���a�      D  , ,  �Z��a�  �Z��b&  ����b&  ����a�  �Z��a�      D  , ,  ����a�  ����b&  �>��b&  �>��a�  ����a�      D  , ,  ����a�  ����b&  ����b&  ����a�  ����a�      D  , ,  �D��a�  �D��b&  ����b&  ����a�  �D��a�      D  , ,  ����h�  ����i`  �T��i`  �T��h�  ����h�      D  , ,  ���h�  ���i`  ����i`  ����h�  ���h�      D  , ,  �Z��h�  �Z��i`  ����i`  ����h�  �Z��h�      D  , ,  ����h�  ����i`  �>��i`  �>��h�  ����h�      D  , ,  ����h�  ����i`  ����i`  ����h�  ����h�      D  , ,  �D��h�  �D��i`  ����i`  ����h�  �D��h�      D  , ,  ����`P  ����`�  �j��`�  �j��`P  ����`P      D  , ,  �"��`P  �"��`�  ����`�  ����`P  �"��`P      D  , ,  �p��`P  �p��`�  ���`�  ���`P  �p��`P      D  , ,  ����`P  ����`�  �T��`�  �T��`P  ����`P      D  , ,  ���`P  ���`�  ����`�  ����`P  ���`P      D  , ,  �Z��`P  �Z��`�  ����`�  ����`P  �Z��`P      D  , ,  ����`P  ����`�  �>��`�  �>��`P  ����`P      D  , ,  ����`P  ����`�  ����`�  ����`P  ����`P      D  , ,  �D��`P  �D��`�  ����`�  ����`P  �D��`P      D  , ,  ����_  ����_�  �j��_�  �j��_  ����_      D  , ,  �"��_  �"��_�  ����_�  ����_  �"��_      D  , ,  �p��_  �p��_�  ���_�  ���_  �p��_      D  , ,  ����_  ����_�  �T��_�  �T��_  ����_      D  , ,  ���_  ���_�  ����_�  ����_  ���_      D  , ,  �Z��_  �Z��_�  ����_�  ����_  �Z��_      D  , ,  ����_  ����_�  �>��_�  �>��_  ����_      D  , ,  ����_  ����_�  ����_�  ����_  ����_      D  , ,  �D��_  �D��_�  ����_�  ����_  �D��_      D  , ,  ����]�  ����^f  �j��^f  �j��]�  ����]�      D  , ,  �"��]�  �"��^f  ����^f  ����]�  �"��]�      D  , ,  �p��]�  �p��^f  ���^f  ���]�  �p��]�      D  , ,  ����]�  ����^f  �T��^f  �T��]�  ����]�      D  , ,  ���]�  ���^f  ����^f  ����]�  ���]�      D  , ,  �Z��]�  �Z��^f  ����^f  ����]�  �Z��]�      D  , ,  ����]�  ����^f  �>��^f  �>��]�  ����]�      D  , ,  ����]�  ����^f  ����^f  ����]�  ����]�      D  , ,  �D��]�  �D��^f  ����^f  ����]�  �D��]�      D  , ,  ����e�  ����fc  ����fc  ����e�  ����e�      D  , ,  �I��e�  �I��fc  ����fc  ����e�  �I��e�      D  , ,  ����e�  ����fc  �-��fc  �-��e�  ����e�      D  , ,  ����e�  ����fc  �{��fc  �{��e�  ����e�      D  , ,  ����\�  ����]&  �j��]&  �j��\�  ����\�      D  , ,  �"��\�  �"��]&  ����]&  ����\�  �"��\�      D  , ,  �p��\�  �p��]&  ���]&  ���\�  �p��\�      D  , ,  ����\�  ����]&  �T��]&  �T��\�  ����\�      D  , ,  ���\�  ���]&  ����]&  ����\�  ���\�      D  , ,  �Z��\�  �Z��]&  ����]&  ����\�  �Z��\�      D  , ,  ����\�  ����]&  �>��]&  �>��\�  ����\�      D  , ,  ����\�  ����]&  ����]&  ����\�  ����\�      D  , ,  �D��\�  �D��]&  ����]&  ����\�  �D��\�      D  , ,  �3��e�  �3��fc  ����fc  ����e�  �3��e�      D  , ,  ����e�  ����fc  ���fc  ���e�  ����e�      D  , ,  ����e�  ����fc  �e��fc  �e��e�  ����e�      D  , ,  ���e�  ���fc  ����fc  ����e�  ���e�      D  , ,  �k��e�  �k��fc  ���fc  ���e�  �k��e�      D  , ,  ����[P  ����[�  �j��[�  �j��[P  ����[P      D  , ,  �"��[P  �"��[�  ����[�  ����[P  �"��[P      D  , ,  �p��[P  �p��[�  ���[�  ���[P  �p��[P      D  , ,  ����[P  ����[�  �T��[�  �T��[P  ����[P      D  , ,  ���[P  ���[�  ����[�  ����[P  ���[P      D  , ,  �Z��[P  �Z��[�  ����[�  ����[P  �Z��[P      D  , ,  ����[P  ����[�  �>��[�  �>��[P  ����[P      D  , ,  ����[P  ����[�  ����[�  ����[P  ����[P      D  , ,  �D��[P  �D��[�  ����[�  ����[P  �D��[P      D  , ,  ���a�  ���b&  ����b&  ����a�  ���a�      D  , ,  �`��a�  �`��b&  ����b&  ����a�  �`��a�      D  , ,  �9��d�  �9��e#  ����e#  ����d�  �9��d�      D  , ,  ~T��`P  ~T��`�  ~���`�  ~���`P  ~T��`P      D  , ,  ����`P  ����`�  �8��`�  �8��`P  ����`P      D  , ,  ����`P  ����`�  ����`�  ����`P  ����`P      D  , ,  �>��`P  �>��`�  ����`�  ����`P  �>��`P      D  , ,  ����e�  ����fc  �_��fc  �_��e�  ����e�      D  , ,  ���e�  ���fc  ����fc  ����e�  ���e�      D  , ,  �e��e�  �e��fc  ����fc  ����e�  �e��e�      D  , ,  ����e�  ����fc  �I��fc  �I��e�  ����e�      D  , ,  ���e�  ���fc  ����fc  ����e�  ���e�      D  , ,  �O��e�  �O��fc  ����fc  ����e�  �O��e�      D  , ,  ����e�  ����fc  �3��fc  �3��e�  ����e�      D  , ,  ~T��]�  ~T��^f  ~���^f  ~���]�  ~T��]�      D  , ,  ����]�  ����^f  �8��^f  �8��]�  ����]�      D  , ,  ����]�  ����^f  ����^f  ����]�  ����]�      D  , ,  �>��]�  �>��^f  ����^f  ����]�  �>��]�      D  , ,  ����]�  ����^f  �"��^f  �"��]�  ����]�      D  , ,  ����]�  ����^f  �p��^f  �p��]�  ����]�      D  , ,  �(��]�  �(��^f  ����^f  ����]�  �(��]�      D  , ,  �v��]�  �v��^f  ���^f  ���]�  �v��]�      D  , ,  ����]�  ����^f  �Z��^f  �Z��]�  ����]�      D  , ,  ���]�  ���^f  ����^f  ����]�  ���]�      D  , ,  �`��]�  �`��^f  ����^f  ����]�  �`��]�      D  , ,  ����`P  ����`�  �"��`�  �"��`P  ����`P      D  , ,  ����`P  ����`�  �p��`�  �p��`P  ����`P      D  , ,  �(��`P  �(��`�  ����`�  ����`P  �(��`P      D  , ,  �v��`P  �v��`�  ���`�  ���`P  �v��`P      D  , ,  ����`P  ����`�  �Z��`�  �Z��`P  ����`P      D  , ,  ���`P  ���`�  ����`�  ����`P  ���`P      D  , ,  �`��`P  �`��`�  ����`�  ����`P  �`��`P      D  , ,  ���h�  ���i`  ����i`  ����h�  ���h�      D  , ,  �`��h�  �`��i`  ����i`  ����h�  �`��h�      D  , ,  ����e�  ����fc  ����fc  ����e�  ����e�      D  , ,  �9��e�  �9��fc  ����fc  ����e�  �9��e�      D  , ,  ~T��a�  ~T��b&  ~���b&  ~���a�  ~T��a�      D  , ,  ����a�  ����b&  �8��b&  �8��a�  ����a�      D  , ,  ����a�  ����b&  ����b&  ����a�  ����a�      D  , ,  �>��a�  �>��b&  ����b&  ����a�  �>��a�      D  , ,  ~T��\�  ~T��]&  ~���]&  ~���\�  ~T��\�      D  , ,  ����\�  ����]&  �8��]&  �8��\�  ����\�      D  , ,  ����\�  ����]&  ����]&  ����\�  ����\�      D  , ,  �>��\�  �>��]&  ����]&  ����\�  �>��\�      D  , ,  ����\�  ����]&  �"��]&  �"��\�  ����\�      D  , ,  ����\�  ����]&  �p��]&  �p��\�  ����\�      D  , ,  �(��\�  �(��]&  ����]&  ����\�  �(��\�      D  , ,  �v��\�  �v��]&  ���]&  ���\�  �v��\�      D  , ,  ����\�  ����]&  �Z��]&  �Z��\�  ����\�      D  , ,  ���\�  ���]&  ����]&  ����\�  ���\�      D  , ,  �`��\�  �`��]&  ����]&  ����\�  �`��\�      D  , ,  ����a�  ����b&  �"��b&  �"��a�  ����a�      D  , ,  ����a�  ����b&  �p��b&  �p��a�  ����a�      D  , ,  �(��a�  �(��b&  ����b&  ����a�  �(��a�      D  , ,  ~T��h�  ~T��i`  ~���i`  ~���h�  ~T��h�      D  , ,  ����h�  ����i`  �8��i`  �8��h�  ����h�      D  , ,  ����h�  ����i`  ����i`  ����h�  ����h�      D  , ,  �>��h�  �>��i`  ����i`  ����h�  �>��h�      D  , ,  ����h�  ����i`  �"��i`  �"��h�  ����h�      D  , ,  }-��e�  }-��fc  }���fc  }���e�  }-��e�      D  , ,  {��e�  {��fc  ���fc  ���e�  {��e�      D  , ,  ~T��_  ~T��_�  ~���_�  ~���_  ~T��_      D  , ,  ����_  ����_�  �8��_�  �8��_  ����_      D  , ,  ����_  ����_�  ����_�  ����_  ����_      D  , ,  �>��_  �>��_�  ����_�  ����_  �>��_      D  , ,  ����h�  ����i`  �p��i`  �p��h�  ����h�      D  , ,  ~T��[P  ~T��[�  ~���[�  ~���[P  ~T��[P      D  , ,  ����[P  ����[�  �8��[�  �8��[P  ����[P      D  , ,  ����[P  ����[�  ����[�  ����[P  ����[P      D  , ,  �>��[P  �>��[�  ����[�  ����[P  �>��[P      D  , ,  ����[P  ����[�  �"��[�  �"��[P  ����[P      D  , ,  ����[P  ����[�  �p��[�  �p��[P  ����[P      D  , ,  �(��[P  �(��[�  ����[�  ����[P  �(��[P      D  , ,  �v��[P  �v��[�  ���[�  ���[P  �v��[P      D  , ,  ����[P  ����[�  �Z��[�  �Z��[P  ����[P      D  , ,  ���[P  ���[�  ����[�  ����[P  ���[P      D  , ,  �`��[P  �`��[�  ����[�  ����[P  �`��[P      D  , ,  ����_  ����_�  �"��_�  �"��_  ����_      D  , ,  ����_  ����_�  �p��_�  �p��_  ����_      D  , ,  �(��_  �(��_�  ����_�  ����_  �(��_      D  , ,  �v��_  �v��_�  ���_�  ���_  �v��_      D  , ,  ����_  ����_�  �Z��_�  �Z��_  ����_      D  , ,  ���_  ���_�  ����_�  ����_  ���_      D  , ,  �`��_  �`��_�  ����_�  ����_  �`��_      D  , ,  �v��a�  �v��b&  ���b&  ���a�  �v��a�      D  , ,  ����a�  ����b&  �Z��b&  �Z��a�  ����a�      D  , ,  �(��h�  �(��i`  ����i`  ����h�  �(��h�      D  , ,  �v��h�  �v��i`  ���i`  ���h�  �v��h�      D  , ,  ����h�  ����i`  �Z��i`  �Z��h�  ����h�      D  , ,  }-��d�  }-��e#  }���e#  }���d�  }-��d�      D  , ,  {��d�  {��e#  ���e#  ���d�  {��d�      D  , ,  ����d�  ����e#  �_��e#  �_��d�  ����d�      D  , ,  ���d�  ���e#  ����e#  ����d�  ���d�      D  , ,  �e��d�  �e��e#  ����e#  ����d�  �e��d�      D  , ,  ����d�  ����e#  �I��e#  �I��d�  ����d�      D  , ,  ���d�  ���e#  ����e#  ����d�  ���d�      D  , ,  �O��d�  �O��e#  ����e#  ����d�  �O��d�      D  , ,  ����d�  ����e#  �3��e#  �3��d�  ����d�      D  , ,  ����d�  ����e#  ����e#  ����d�  ����d�      D  , ,  �v��Z  �v��Z�  ���Z�  ���Z  �v��Z      D  , ,  ����Z  ����Z�  �Z��Z�  �Z��Z  ����Z      D  , ,  ���Z  ���Z�  ����Z�  ����Z  ���Z      D  , ,  �`��Z  �`��Z�  ����Z�  ����Z  �`��Z      D  , ,  ~T��Z  ~T��Z�  ~���Z�  ~���Z  ~T��Z      D  , ,  ����Z  ����Z�  �8��Z�  �8��Z  ����Z      D  , ,  ����Z  ����Z�  ����Z�  ����Z  ����Z      D  , ,  �>��Z  �>��Z�  ����Z�  ����Z  �>��Z      D  , ,  ����Z  ����Z�  �"��Z�  �"��Z  ����Z      D  , ,  ����Z  ����Z�  �p��Z�  �p��Z  ����Z      D  , ,  ~T��X�  ~T��Yf  ~���Yf  ~���X�  ~T��X�      D  , ,  ����X�  ����Yf  �8��Yf  �8��X�  ����X�      D  , ,  ����X�  ����Yf  ����Yf  ����X�  ����X�      D  , ,  �>��X�  �>��Yf  ����Yf  ����X�  �>��X�      D  , ,  ����X�  ����Yf  �"��Yf  �"��X�  ����X�      D  , ,  ����X�  ����Yf  �p��Yf  �p��X�  ����X�      D  , ,  �(��X�  �(��Yf  ����Yf  ����X�  �(��X�      D  , ,  �v��X�  �v��Yf  ���Yf  ���X�  �v��X�      D  , ,  ����X�  ����Yf  �Z��Yf  �Z��X�  ����X�      D  , ,  ���X�  ���Yf  ����Yf  ����X�  ���X�      D  , ,  �`��X�  �`��Yf  ����Yf  ����X�  �`��X�      D  , ,  �(��Z  �(��Z�  ����Z�  ����Z  �(��Z      D  , ,  ����Z  ����Z�  �j��Z�  �j��Z  ����Z      D  , ,  �"��Z  �"��Z�  ����Z�  ����Z  �"��Z      D  , ,  �p��Z  �p��Z�  ���Z�  ���Z  �p��Z      D  , ,  ����Z  ����Z�  �T��Z�  �T��Z  ����Z      D  , ,  ���Z  ���Z�  ����Z�  ����Z  ���Z      D  , ,  �Z��Z  �Z��Z�  ����Z�  ����Z  �Z��Z      D  , ,  ����Z  ����Z�  �>��Z�  �>��Z  ����Z      D  , ,  ����Z  ����Z�  ����Z�  ����Z  ����Z      D  , ,  ����X�  ����Yf  �j��Yf  �j��X�  ����X�      D  , ,  �"��X�  �"��Yf  ����Yf  ����X�  �"��X�      D  , ,  �p��X�  �p��Yf  ���Yf  ���X�  �p��X�      D  , ,  ����X�  ����Yf  �T��Yf  �T��X�  ����X�      D  , ,  ���X�  ���Yf  ����Yf  ����X�  ���X�      D  , ,  �Z��X�  �Z��Yf  ����Yf  ����X�  �Z��X�      D  , ,  ����X�  ����Yf  �>��Yf  �>��X�  ����X�      D  , ,  ����X�  ����Yf  ����Yf  ����X�  ����X�      D  , ,  �D��X�  �D��Yf  ����Yf  ����X�  �D��X�      D  , ,  �D��Z  �D��Z�  ����Z�  ����Z  �D��Z      D  , ,  ����iB  ����i�  �n��i�  �n��iB  ����iB      D  , ,  ����iB  ����i�  �R��i�  �R��iB  ����iB      D  , ,  ����iB  ����i�  �6��i�  �6��iB  ����iB      D  , ,  ����iB  ����i�  ���i�  ���iB  ����iB      D  , ,  h��iB  h��i�  ���i�  ���iB  h��iB      D  , , L��iB L��i� ���i� ���iB L��iB      D  , , 0��iB 0��i� ���i� ���iB 0��iB      D  , , 	��iB 	��i� 	���i� 	���iB 	��iB      D  , , ���iB ���i� ���i� ���iB ���iB      D  , , ���iB ���i� r��i� r��iB ���iB      D  , , ���iB ���i� V��i� V��iB ���iB      D  , , ���m ���m� ���m� ���m ���m      D  , , ���m ���m� r��m� r��m ���m      D  , , ���m ���m� V��m� V��m ���m      D  , ,  ����p�  ����qX  �n��qX  �n��p�  ����p�      D  , ,  ����p�  ����qX  �R��qX  �R��p�  ����p�      D  , ,  ����p�  ����qX  �6��qX  �6��p�  ����p�      D  , ,  ����p�  ����qX  ���qX  ���p�  ����p�      D  , ,  h��p�  h��qX  ���qX  ���p�  h��p�      D  , , L��p� L��qX ���qX ���p� L��p�      D  , , 0��p� 0��qX ���qX ���p� 0��p�      D  , , 	��p� 	��qX 	���qX 	���p� 	��p�      D  , , ���p� ���qX ���qX ���p� ���p�      D  , , ���p� ���qX r��qX r��p� ���p�      D  , , ���p� ���qX V��qX V��p� ���p�      D  , ,  ����k�  ����lX  �n��lX  �n��k�  ����k�      D  , ,  ����k�  ����lX  �R��lX  �R��k�  ����k�      D  , ,  ����k�  ����lX  �6��lX  �6��k�  ����k�      D  , ,  ����k�  ����lX  ���lX  ���k�  ����k�      D  , ,  h��k�  h��lX  ���lX  ���k�  h��k�      D  , , L��k� L��lX ���lX ���k� L��k�      D  , , 0��k� 0��lX ���lX ���k� 0��k�      D  , , 	��k� 	��lX 	���lX 	���k� 	��k�      D  , , ���k� ���lX ���lX ���k� ���k�      D  , , ���k� ���lX r��lX r��k� ���k�      D  , , ���k� ���lX V��lX V��k� ���k�      D  , ,  ����o�  ����p  �n��p  �n��o�  ����o�      D  , ,  ����o�  ����p  �R��p  �R��o�  ����o�      D  , ,  ����j�  ����k  �n��k  �n��j�  ����j�      D  , ,  ����j�  ����k  �R��k  �R��j�  ����j�      D  , ,  ����j�  ����k  �6��k  �6��j�  ����j�      D  , ,  ����j�  ����k  ���k  ���j�  ����j�      D  , ,  h��j�  h��k  ���k  ���j�  h��j�      D  , , L��j� L��k ���k ���j� L��j�      D  , , 0��j� 0��k ���k ���j� 0��j�      D  , , 	��j� 	��k 	���k 	���j� 	��j�      D  , , ���j� ���k ���k ���j� ���j�      D  , , ���j� ���k r��k r��j� ���j�      D  , , ���j� ���k V��k V��j� ���j�      D  , ,  ����o�  ����p  �6��p  �6��o�  ����o�      D  , ,  ����o�  ����p  ���p  ���o�  ����o�      D  , ,  h��o�  h��p  ���p  ���o�  h��o�      D  , , L��o� L��p ���p ���o� L��o�      D  , , 0��o� 0��p ���p ���o� 0��o�      D  , , 	��o� 	��p 	���p 	���o� 	��o�      D  , , ���o� ���p ���p ���o� ���o�      D  , , ���o� ���p r��p r��o� ���o�      D  , , ���o� ���p V��p V��o� ���o�      D  , ,  ����r  ����r�  �n��r�  �n��r  ����r      D  , , ���nB ���n� r��n� r��nB ���nB      D  , , ���nB ���n� V��n� V��nB ���nB      D  , , ���r ���r� V��r� V��r ���r      D  , ,  ����m  ����m�  �n��m�  �n��m  ����m      D  , ,  ����m  ����m�  �R��m�  �R��m  ����m      D  , ,  ����m  ����m�  �6��m�  �6��m  ����m      D  , ,  ����m  ����m�  ���m�  ���m  ����m      D  , ,  h��m  h��m�  ���m�  ���m  h��m      D  , , L��m L��m� ���m� ���m L��m      D  , , 0��m 0��m� ���m� ���m 0��m      D  , , 	��m 	��m� 	���m� 	���m 	��m      D  , ,  ����r  ����r�  �R��r�  �R��r  ����r      D  , ,  ����r  ����r�  �6��r�  �6��r  ����r      D  , ,  ����r  ����r�  ���r�  ���r  ����r      D  , ,  h��r  h��r�  ���r�  ���r  h��r      D  , , L��r L��r� ���r� ���r L��r      D  , , 0��r 0��r� ���r� ���r 0��r      D  , , 	��r 	��r� 	���r� 	���r 	��r      D  , , ���r ���r� ���r� ���r ���r      D  , , ���r ���r� r��r� r��r ���r      D  , ,  ����nB  ����n�  �n��n�  �n��nB  ����nB      D  , ,  ����nB  ����n�  �R��n�  �R��nB  ����nB      D  , ,  ����nB  ����n�  �6��n�  �6��nB  ����nB      D  , ,  ����nB  ����n�  ���n�  ���nB  ����nB      D  , ,  h��nB  h��n�  ���n�  ���nB  h��nB      D  , , L��nB L��n� ���n� ���nB L��nB      D  , , 0��nB 0��n� ���n� ���nB 0��nB      D  , , 	��nB 	��n� 	���n� 	���nB 	��nB      D  , , ���nB ���n� ���n� ���nB ���nB      D  , ,  � ���  � ���I  Ȗ���I  Ȗ���  � ���      D  , ,  � ���E  � ����  Ȗ����  Ȗ���E  � ���E      D  , ,  � ��}3  � ��}�  Ȗ��}�  Ȗ��}3  � ��}3      D  , ,  � ��{�  � ��|�  Ȗ��|�  Ȗ��{�  � ��{�      D  , ,  � ����  � ���  Ȗ���  Ȗ����  � ����      D  , ,  � ��~s  � ��	  Ȗ��	  Ȗ��~s  � ��~s      D  , ,  �X���E  �X����  ������  �����E  �X���E      D  , ,  ̜��}3  ̜��}�  �2��}�  �2��}3  ̜��}3      D  , ,  �8��}3  �8��}�  ����}�  ����}3  �8��}3      D  , ,  ̜���  ̜���I  �2���I  �2���  ̜���      D  , ,  �8���  �8���I  �����I  �����  �8���      D  , ,  ̜���E  ̜����  �2����  �2���E  ̜���E      D  , ,  ̜��{�  ̜��|�  �2��|�  �2��{�  ̜��{�      D  , ,  �8��{�  �8��|�  ����|�  ����{�  �8��{�      D  , ,  �����E  ������  ϊ����  ϊ���E  �����E      D  , ,  �X����  �X���  �����  ������  �X����      D  , ,  �8���E  �8����  ������  �����E  �8���E      D  , ,  ̜��~s  ̜��	  �2��	  �2��~s  ̜��~s      D  , ,  �8��~s  �8��	  ����	  ����~s  �8��~s      D  , ,  ̜����  ̜���  �2���  �2����  ̜����      D  , ,  ������  �����  ϊ���  ϊ����  ������      D  , ,  �8����  �8���  �����  ������  �8����      D  , ,  ������  �����  ����  �����  ������      D  , ,  �����E  ������  ������  �����E  �����E      D  , ,  ������  �����  �^���  �^����  ������      D  , ,  � ����  � ���  �����  ������  � ����      D  , ,  �d����  �d���  �����  ������  �d����      D  , ,  ����~s  ����	  �^��	  �^��~s  ����~s      D  , ,  ż����  ż���  �R���  �R����  ż����      D  , ,  ����{�  ����|�  ����|�  ����{�  ����{�      D  , ,  ����{�  ����|�  �&��|�  �&��{�  ����{�      D  , ,  �,��{�  �,��|�  ����|�  ����{�  �,��{�      D  , ,  ����{�  ����|�  �^��|�  �^��{�  ����{�      D  , ,  �d��{�  �d��|�  ����|�  ����{�  �d��{�      D  , ,  �d��}3  �d��}�  ����}�  ����}3  �d��}3      D  , ,  �L���E  �L����  ������  �����E  �L���E      D  , ,  �����E  ������  �&����  �&���E  �����E      D  , ,  �����  �����I  �����I  �����  �����      D  , ,  �����  �����I  �&���I  �&���  �����      D  , ,  �,���  �,���I  �����I  �����  �,���      D  , ,  �����E  ������  �~����  �~���E  �����E      D  , ,  �,���E  �,����  ������  �����E  �,���E      D  , ,  �����E  ������  �����  ����E  �����E      D  , ,  �����E  ������  �^����  �^���E  �����E      D  , ,  �����  �����I  �^���I  �^���  �����      D  , ,  �d���  �d���I  �����I  �����  �d���      D  , ,  �L����  �L���  �����  ������  �L����      D  , ,  ����}3  ����}�  ����}�  ����}3  ����}3      D  , ,  ����}3  ����}�  �&��}�  �&��}3  ����}3      D  , ,  �d��~s  �d��	  ����	  ����~s  �d��~s      D  , ,  �,��}3  �,��}�  ����}�  ����}3  �,��}3      D  , ,  ����}3  ����}�  �^��}�  �^��}3  ����}3      D  , ,  ż���E  ż����  �R����  �R���E  ż���E      D  , ,  ������  �����  �&���  �&����  ������      D  , ,  ������  �����  �~���  �~����  ������      D  , ,  �,����  �,���  �����  ������  �,����      D  , ,  ������  �����  �����  ������  ������      D  , ,  ����~s  ����	  ����	  ����~s  ����~s      D  , ,  ����~s  ����	  �&��	  �&��~s  ����~s      D  , ,  �,��~s  �,��	  ����	  ����~s  �,��~s      D  , ,  � ���E  � ����  ������  �����E  � ���E      D  , ,  �d���E  �d����  ������  �����E  �d���E      D  , ,  ����q�  ����r   �v��r   �v��q�  ����q�      D  , ,  �.��q�  �.��r   ����r   ����q�  �.��q�      D  , ,  �|��q�  �|��r   ���r   ���q�  �|��q�      D  , ,  ����q�  ����r   �`��r   �`��q�  ����q�      D  , ,  ���q�  ���r   ����r   ����q�  ���q�      D  , ,  �f��q�  �f��r   ����r   ����q�  �f��q�      D  , ,  ���pJ  ���p�  ����p�  ����pJ  ���pJ      D  , ,  �f��pJ  �f��p�  ����p�  ����pJ  �f��pJ      D  , ,  �|��j
  �|��j�  ���j�  ���j
  �|��j
      D  , ,  ����j
  ����j�  �`��j�  �`��j
  ����j
      D  , ,  ���j
  ���j�  ����j�  ����j
  ���j
      D  , ,  �f��j
  �f��j�  ����j�  ����j
  �f��j
      D  , ,  �|��o
  �|��o�  ���o�  ���o
  �|��o
      D  , ,  ����o
  ����o�  �`��o�  �`��o
  ����o
      D  , ,  ���o
  ���o�  ����o�  ����o
  ���o
      D  , ,  �f��o
  �f��o�  ����o�  ����o
  �f��o
      D  , ,  ����o
  ����o�  �v��o�  �v��o
  ����o
      D  , ,  �.��o
  �.��o�  ����o�  ����o
  �.��o
      D  , ,  ����j
  ����j�  �v��j�  �v��j
  ����j
      D  , ,  ����kJ  ����k�  �v��k�  �v��kJ  ����kJ      D  , ,  �.��kJ  �.��k�  ����k�  ����kJ  �.��kJ      D  , ,  �|��kJ  �|��k�  ���k�  ���kJ  �|��kJ      D  , ,  ����kJ  ����k�  �`��k�  �`��kJ  ����kJ      D  , ,  ���kJ  ���k�  ����k�  ����kJ  ���kJ      D  , ,  �f��kJ  �f��k�  ����k�  ����kJ  �f��kJ      D  , ,  �.��j
  �.��j�  ����j�  ����j
  �.��j
      D  , ,  ����pJ  ����p�  �v��p�  �v��pJ  ����pJ      D  , ,  ����m�  ����n`  �v��n`  �v��m�  ����m�      D  , ,  �.��m�  �.��n`  ����n`  ����m�  �.��m�      D  , ,  �|��m�  �|��n`  ���n`  ���m�  �|��m�      D  , ,  ����m�  ����n`  �`��n`  �`��m�  ����m�      D  , ,  ���m�  ���n`  ����n`  ����m�  ���m�      D  , ,  �f��m�  �f��n`  ����n`  ����m�  �f��m�      D  , ,  �.��pJ  �.��p�  ����p�  ����pJ  �.��pJ      D  , ,  ����l�  ����m   �v��m   �v��l�  ����l�      D  , ,  �.��l�  �.��m   ����m   ����l�  �.��l�      D  , ,  �|��l�  �|��m   ���m   ���l�  �|��l�      D  , ,  ����l�  ����m   �`��m   �`��l�  ����l�      D  , ,  ���l�  ���m   ����m   ����l�  ���l�      D  , ,  �f��l�  �f��m   ����m   ����l�  �f��l�      D  , ,  �|��pJ  �|��p�  ���p�  ���pJ  �|��pJ      D  , ,  ����pJ  ����p�  �`��p�  �`��pJ  ����pJ      D  , ,  �|��]�  �|��^f  ���^f  ���]�  �|��]�      D  , ,  ����h�  ����i`  �v��i`  �v��h�  ����h�      D  , ,  �.��h�  �.��i`  ����i`  ����h�  �.��h�      D  , ,  �|��h�  �|��i`  ���i`  ���h�  �|��h�      D  , ,  ����h�  ����i`  �`��i`  �`��h�  ����h�      D  , ,  ���h�  ���i`  ����i`  ����h�  ���h�      D  , ,  �f��h�  �f��i`  ����i`  ����h�  �f��h�      D  , ,  ����]�  ����^f  �`��^f  �`��]�  ����]�      D  , ,  ���]�  ���^f  ����^f  ����]�  ���]�      D  , ,  �f��]�  �f��^f  ����^f  ����]�  �f��]�      D  , ,  ����`P  ����`�  �v��`�  �v��`P  ����`P      D  , ,  �.��`P  �.��`�  ����`�  ����`P  �.��`P      D  , ,  �|��`P  �|��`�  ���`�  ���`P  �|��`P      D  , ,  ����`P  ����`�  �`��`�  �`��`P  ����`P      D  , ,  ���`P  ���`�  ����`�  ����`P  ���`P      D  , ,  �f��`P  �f��`�  ����`�  ����`P  �f��`P      D  , ,  ����d�  ����e#  ����e#  ����d�  ����d�      D  , ,  �?��d�  �?��e#  ����e#  ����d�  �?��d�      D  , ,  ����[P  ����[�  �v��[�  �v��[P  ����[P      D  , ,  �.��[P  �.��[�  ����[�  ����[P  �.��[P      D  , ,  �|��[P  �|��[�  ���[�  ���[P  �|��[P      D  , ,  ����[P  ����[�  �`��[�  �`��[P  ����[P      D  , ,  ���[P  ���[�  ����[�  ����[P  ���[P      D  , ,  �f��[P  �f��[�  ����[�  ����[P  �f��[P      D  , ,  ����d�  ����e#  �O��e#  �O��d�  ����d�      D  , ,  ���d�  ���e#  ����e#  ����d�  ���d�      D  , ,  ����a�  ����b&  �v��b&  �v��a�  ����a�      D  , ,  �.��a�  �.��b&  ����b&  ����a�  �.��a�      D  , ,  �|��a�  �|��b&  ���b&  ���a�  �|��a�      D  , ,  ����a�  ����b&  �`��b&  �`��a�  ����a�      D  , ,  ���a�  ���b&  ����b&  ����a�  ���a�      D  , ,  ����_  ����_�  �v��_�  �v��_  ����_      D  , ,  �.��_  �.��_�  ����_�  ����_  �.��_      D  , ,  �|��_  �|��_�  ���_�  ���_  �|��_      D  , ,  ����_  ����_�  �`��_�  �`��_  ����_      D  , ,  ���_  ���_�  ����_�  ����_  ���_      D  , ,  ����Z  ����Z�  �v��Z�  �v��Z  ����Z      D  , ,  �.��Z  �.��Z�  ����Z�  ����Z  �.��Z      D  , ,  �|��Z  �|��Z�  ���Z�  ���Z  �|��Z      D  , ,  ����Z  ����Z�  �`��Z�  �`��Z  ����Z      D  , ,  ���Z  ���Z�  ����Z�  ����Z  ���Z      D  , ,  �f��Z  �f��Z�  ����Z�  ����Z  �f��Z      D  , ,  �f��_  �f��_�  ����_�  ����_  �f��_      D  , ,  �f��a�  �f��b&  ����b&  ����a�  �f��a�      D  , ,  �U��d�  �U��e#  ����e#  ����d�  �U��d�      D  , ,  ����d�  ����e#  �9��e#  �9��d�  ����d�      D  , ,  ����]�  ����^f  �v��^f  �v��]�  ����]�      D  , ,  �.��]�  �.��^f  ����^f  ����]�  �.��]�      D  , ,  ����\�  ����]&  �v��]&  �v��\�  ����\�      D  , ,  �.��\�  �.��]&  ����]&  ����\�  �.��\�      D  , ,  �|��\�  �|��]&  ���]&  ���\�  �|��\�      D  , ,  ����\�  ����]&  �`��]&  �`��\�  ����\�      D  , ,  ���\�  ���]&  ����]&  ����\�  ���\�      D  , ,  �f��\�  �f��]&  ����]&  ����\�  �f��\�      D  , ,  ����e�  ����fc  �O��fc  �O��e�  ����e�      D  , ,  ���e�  ���fc  ����fc  ����e�  ���e�      D  , ,  �U��e�  �U��fc  ����fc  ����e�  �U��e�      D  , ,  ����e�  ����fc  �9��fc  �9��e�  ����e�      D  , ,  ����e�  ����fc  ����fc  ����e�  ����e�      D  , ,  �?��e�  �?��fc  ����fc  ����e�  �?��e�      D  , ,  ����X�  ����Yf  �v��Yf  �v��X�  ����X�      D  , ,  �.��X�  �.��Yf  ����Yf  ����X�  �.��X�      D  , ,  �|��X�  �|��Yf  ���Yf  ���X�  �|��X�      D  , ,  ����X�  ����Yf  �`��Yf  �`��X�  ����X�      D  , ,  ���X�  ���Yf  ����Yf  ����X�  ���X�      D  , ,  �f��X�  �f��Yf  ����Yf  ����X�  �f��X�      D  , ,  ����h  ����h�  ���h�  ���h  ����h      D  , ,  h��h  h��h�  ���h�  ���h  h��h      D  , , L��h L��h� ���h� ���h L��h      D  , , 0��h 0��h� ���h� ���h 0��h      D  , , 	��h 	��h� 	���h� 	���h 	��h      D  , ,  ����^�  ����_G  ����_G  ����^�  ����^�      D  , , ���^� ���_G p��_G p��^� ���^�      D  , , ���^� ���_G T��_G T��^� ���^�      D  , , ���^� ���_G 8��_G 8��^� ���^�      D  , , 
���^� 
���_G ��_G ��^� 
���^�      D  , , j��^� j��_G  ��_G  ��^� j��^�      D  , ,  ����[�  ����\6  �6��\6  �6��[�  ����[�      D  , ,  ����[�  ����\6  ���\6  ���[�  ����[�      D  , ,  h��[�  h��\6  ���\6  ���[�  h��[�      D  , , L��[� L��\6 ���\6 ���[� L��[�      D  , , 0��[� 0��\6 ���\6 ���[� 0��[�      D  , , 	��[� 	��\6 	���\6 	���[� 	��[�      D  , , ���[� ���\6 ���\6 ���[� ���[�      D  , , ���[� ���\6 r��\6 r��[� ���[�      D  , , ���[� ���\6 V��\6 V��[� ���[�      D  , , ���h ���h� ���h� ���h ���h      D  , , ���h ���h� r��h� r��h ���h      D  , , ���h ���h� V��h� V��h ���h      D  , ,  ����f�  ����gX  �6��gX  �6��f�  ����f�      D  , ,  ����f�  ����gX  ���gX  ���f�  ����f�      D  , ,  h��f�  h��gX  ���gX  ���f�  h��f�      D  , , L��f� L��gX ���gX ���f� L��f�      D  , , 0��f� 0��gX ���gX ���f� 0��f�      D  , , 	��f� 	��gX 	���gX 	���f� 	��f�      D  , , ���f� ���gX ���gX ���f� ���f�      D  , , ���f� ���gX r��gX r��f� ���f�      D  , , ���f� ���gX V��gX V��f� ���f�      D  , , N��^� N��_G ���_G ���^� N��^�      D  , , j��_� j��`�  ��`�  ��_� j��_�      D  , , N��_� N��`� ���`� ���_� N��_�      D  , ,  ����c  ����c�  �6��c�  �6��c  ����c      D  , ,  ����c  ����c�  ���c�  ���c  ����c      D  , ,  h��c  h��c�  ���c�  ���c  h��c      D  , , L��c L��c� ���c� ���c L��c      D  , , 0��c 0��c� ���c� ���c 0��c      D  , , 	��c 	��c� 	���c� 	���c 	��c      D  , , ���c ���c� ���c� ���c ���c      D  , , ���c ���c� r��c� r��c ���c      D  , , ���c ���c� V��c� V��c ���c      D  , , ���e� ���f ���f ���e� ���e�      D  , , ���e� ���f r��f r��e� ���e�      D  , , ���e� ���f V��f V��e� ���e�      D  , ,  ����dB  ����d�  �6��d�  �6��dB  ����dB      D  , ,  ����dB  ����d�  ���d�  ���dB  ����dB      D  , ,  h��dB  h��d�  ���d�  ���dB  h��dB      D  , , L��dB L��d� ���d� ���dB L��dB      D  , , 0��dB 0��d� ���d� ���dB 0��dB      D  , , 	��dB 	��d� 	���d� 	���dB 	��dB      D  , , ���dB ���d� ���d� ���dB ���dB      D  , , ���dB ���d� r��d� r��dB ���dB      D  , , ���dB ���d� V��d� V��dB ���dB      D  , ,  ���_�  ���`�  ����`�  ����_�  ���_�      D  , ,  ����_�  ����`�  ����`�  ����_�  ����_�      D  , , ���_� ���`� p��`� p��_� ���_�      D  , , ���_� ���`� T��`� T��_� ���_�      D  , , ���_� ���`� 8��`� 8��_� ���_�      D  , , 
���_� 
���`� ��`� ��_� 
���_�      D  , ,  ����e�  ����f  �6��f  �6��e�  ����e�      D  , ,  ����e�  ����f  ���f  ���e�  ����e�      D  , ,  h��e�  h��f  ���f  ���e�  h��e�      D  , , L��e� L��f ���f ���e� L��e�      D  , , 0��e� 0��f ���f ���e� 0��e�      D  , , 	��e� 	��f 	���f 	���e� 	��e�      D  , ,  ���^�  ���_G  ����_G  ����^�  ���^�      D  , ,  ����h  ����h�  �6��h�  �6��h  ����h      D  , ,  ����c  ����c�  �R��c�  �R��c  ����c      D  , ,  ����dB  ����d�  �n��d�  �n��dB  ����dB      D  , ,  ����e�  ����f  �n��f  �n��e�  ����e�      D  , ,  ����e�  ����f  �R��f  �R��e�  ����e�      D  , ,  ����dB  ����d�  �R��d�  �R��dB  ����dB      D  , ,  ����[�  ����\6  �n��\6  �n��[�  ����[�      D  , ,  �J��_�  �J��`�  ����`�  ����_�  �J��_�      D  , ,  �.��_�  �.��`�  ����`�  ����_�  �.��_�      D  , ,  ����[�  ����\6  �R��\6  �R��[�  ����[�      D  , ,  ����f�  ����gX  �n��gX  �n��f�  ����f�      D  , ,  �J��^�  �J��_G  ����_G  ����^�  �J��^�      D  , ,  �.��^�  �.��_G  ����_G  ����^�  �.��^�      D  , ,  ����f�  ����gX  �R��gX  �R��f�  ����f�      D  , ,  ����h  ����h�  �n��h�  �n��h  ����h      D  , ,  ����h  ����h�  �R��h�  �R��h  ����h      D  , ,  ����c  ����c�  �n��c�  �n��c  ����c      D  , ,  ����Z`  ����Z�  �n��Z�  �n��Z`  ����Z`      D  , ,  ����Z`  ����Z�  �R��Z�  �R��Z`  ����Z`      D  , ,  ����Y   ����Y�  �n��Y�  �n��Y   ����Y       D  , ,  ����Y   ����Y�  �R��Y�  �R��Y   ����Y       D  , ,  ����W�  ����Xv  �n��Xv  �n��W�  ����W�      D  , ,  ����W�  ����Xv  �R��Xv  �R��W�  ����W�      D  , ,  ����V�  ����W6  �n��W6  �n��V�  ����V�      D  , ,  ����V�  ����W6  �R��W6  �R��V�  ����V�      D  , ,  ����U`  ����U�  �n��U�  �n��U`  ����U`      D  , ,  ����U`  ����U�  �R��U�  �R��U`  ����U`      D  , ,  ����T   ����T�  �n��T�  �n��T   ����T       D  , ,  ����T   ����T�  �R��T�  �R��T   ����T       D  , ,  ����R�  ����Sv  �n��Sv  �n��R�  ����R�      D  , ,  ����R�  ����Sv  �R��Sv  �R��R�  ����R�      D  , ,  ����Q�  ����R6  �n��R6  �n��Q�  ����Q�      D  , ,  ����Q�  ����R6  �R��R6  �R��Q�  ����Q�      D  , ,  ����P`  ����P�  �n��P�  �n��P`  ����P`      D  , ,  ����P`  ����P�  �R��P�  �R��P`  ����P`      D  , ,  ����O   ����O�  �n��O�  �n��O   ����O       D  , ,  ����O   ����O�  �R��O�  �R��O   ����O       D  , ,  ����M�  ����Nv  �n��Nv  �n��M�  ����M�      D  , ,  ����M�  ����Nv  �R��Nv  �R��M�  ����M�      D  , ,  ����L�  ����M6  �n��M6  �n��L�  ����L�      D  , ,  ����L�  ����M6  �R��M6  �R��L�  ����L�      D  , , 0��W� 0��Xv ���Xv ���W� 0��W�      D  , , 0��V� 0��W6 ���W6 ���V� 0��V�      D  , , 0��U` 0��U� ���U� ���U` 0��U`      D  , , 0��Z` 0��Z� ���Z� ���Z` 0��Z`      D  , , 0��T  0��T� ���T� ���T  0��T       D  , , 0��R� 0��Sv ���Sv ���R� 0��R�      D  , , 0��Q� 0��R6 ���R6 ���Q� 0��Q�      D  , , 0��Y  0��Y� ���Y� ���Y  0��Y       D  , , 0��P` 0��P� ���P� ���P` 0��P`      D  , , 0��O  0��O� ���O� ���O  0��O       D  , , 0��M� 0��Nv ���Nv ���M� 0��M�      D  , , 0��L� 0��M6 ���M6 ���L� 0��L�      D  , , ���U` ���U� ���U� ���U` ���U`      D  , , ���U` ���U� r��U� r��U` ���U`      D  , , ���U` ���U� V��U� V��U` ���U`      D  , , ���W� ���Xv r��Xv r��W� ���W�      D  , , 	��Z` 	��Z� 	���Z� 	���Z` 	��Z`      D  , , ���W� ���Xv V��Xv V��W� ���W�      D  , , 	��T  	��T� 	���T� 	���T  	��T       D  , , ���T  ���T� ���T� ���T  ���T       D  , , ���T  ���T� r��T� r��T  ���T       D  , , ���T  ���T� V��T� V��T  ���T       D  , , ���Z` ���Z� ���Z� ���Z` ���Z`      D  , , 	��W� 	��Xv 	���Xv 	���W� 	��W�      D  , , 	��V� 	��W6 	���W6 	���V� 	��V�      D  , , ���V� ���W6 ���W6 ���V� ���V�      D  , , ���V� ���W6 r��W6 r��V� ���V�      D  , , 	��Y  	��Y� 	���Y� 	���Y  	��Y       D  , , ���Y  ���Y� ���Y� ���Y  ���Y       D  , , ���V� ���W6 V��W6 V��V� ���V�      D  , , ���Y  ���Y� r��Y� r��Y  ���Y       D  , , ���Y  ���Y� V��Y� V��Y  ���Y       D  , , ���W� ���Xv ���Xv ���W� ���W�      D  , , ���Z` ���Z� r��Z� r��Z` ���Z`      D  , , ���Z` ���Z� V��Z� V��Z` ���Z`      D  , , 	��U` 	��U� 	���U� 	���U` 	��U`      D  , , L��T  L��T� ���T� ���T  L��T       D  , , L��W� L��Xv ���Xv ���W� L��W�      D  , ,  ����W�  ����Xv  �6��Xv  �6��W�  ����W�      D  , ,  ����Z`  ����Z�  �6��Z�  �6��Z`  ����Z`      D  , ,  h��Z`  h��Z�  ���Z�  ���Z`  h��Z`      D  , , L��Z` L��Z� ���Z� ���Z` L��Z`      D  , ,  ����U`  ����U�  �6��U�  �6��U`  ����U`      D  , ,  ����Y   ����Y�  �6��Y�  �6��Y   ����Y       D  , ,  ����U`  ����U�  ���U�  ���U`  ����U`      D  , ,  ����Y   ����Y�  ���Y�  ���Y   ����Y       D  , ,  h��Y   h��Y�  ���Y�  ���Y   h��Y       D  , ,  h��U`  h��U�  ���U�  ���U`  h��U`      D  , , L��Y  L��Y� ���Y� ���Y  L��Y       D  , , L��U` L��U� ���U� ���U` L��U`      D  , ,  ����Z`  ����Z�  ���Z�  ���Z`  ����Z`      D  , ,  ����V�  ����W6  �6��W6  �6��V�  ����V�      D  , ,  ����V�  ����W6  ���W6  ���V�  ����V�      D  , ,  h��V�  h��W6  ���W6  ���V�  h��V�      D  , , L��V� L��W6 ���W6 ���V� L��V�      D  , ,  ����W�  ����Xv  ���Xv  ���W�  ����W�      D  , ,  h��W�  h��Xv  ���Xv  ���W�  h��W�      D  , ,  ����T   ����T�  �6��T�  �6��T   ����T       D  , ,  ����T   ����T�  ���T�  ���T   ����T       D  , ,  h��T   h��T�  ���T�  ���T   h��T       D  , ,  h��P`  h��P�  ���P�  ���P`  h��P`      D  , , L��P` L��P� ���P� ���P` L��P`      D  , ,  h��R�  h��Sv  ���Sv  ���R�  h��R�      D  , ,  ����Q�  ����R6  �6��R6  �6��Q�  ����Q�      D  , ,  ����Q�  ����R6  ���R6  ���Q�  ����Q�      D  , ,  ����O   ����O�  �6��O�  �6��O   ����O       D  , ,  ����O   ����O�  ���O�  ���O   ����O       D  , ,  h��O   h��O�  ���O�  ���O   h��O       D  , , L��O  L��O� ���O� ���O  L��O       D  , ,  h��Q�  h��R6  ���R6  ���Q�  h��Q�      D  , , L��Q� L��R6 ���R6 ���Q� L��Q�      D  , , L��R� L��Sv ���Sv ���R� L��R�      D  , ,  ����M�  ����Nv  �6��Nv  �6��M�  ����M�      D  , ,  ����M�  ����Nv  ���Nv  ���M�  ����M�      D  , ,  h��M�  h��Nv  ���Nv  ���M�  h��M�      D  , , L��M� L��Nv ���Nv ���M� L��M�      D  , ,  ����R�  ����Sv  �6��Sv  �6��R�  ����R�      D  , ,  ����R�  ����Sv  ���Sv  ���R�  ����R�      D  , ,  ����P`  ����P�  �6��P�  �6��P`  ����P`      D  , ,  ����L�  ����M6  �6��M6  �6��L�  ����L�      D  , ,  ����L�  ����M6  ���M6  ���L�  ����L�      D  , ,  h��L�  h��M6  ���M6  ���L�  h��L�      D  , , L��L� L��M6 ���M6 ���L� L��L�      D  , ,  ����P`  ����P�  ���P�  ���P`  ����P`      D  , , ���O  ���O� r��O� r��O  ���O       D  , , ���O  ���O� V��O� V��O  ���O       D  , , ���Q� ���R6 r��R6 r��Q� ���Q�      D  , , 	��P` 	��P� 	���P� 	���P` 	��P`      D  , , ���P` ���P� ���P� ���P` ���P`      D  , , ���P` ���P� r��P� r��P` ���P`      D  , , ���P` ���P� V��P� V��P` ���P`      D  , , ���Q� ���R6 V��R6 V��Q� ���Q�      D  , , ���R� ���Sv V��Sv V��R� ���R�      D  , , 	��M� 	��Nv 	���Nv 	���M� 	��M�      D  , , ���M� ���Nv ���Nv ���M� ���M�      D  , , ���M� ���Nv r��Nv r��M� ���M�      D  , , ���M� ���Nv V��Nv V��M� ���M�      D  , , 	��R� 	��Sv 	���Sv 	���R� 	��R�      D  , , ���R� ���Sv ���Sv ���R� ���R�      D  , , ���R� ���Sv r��Sv r��R� ���R�      D  , , 	��Q� 	��R6 	���R6 	���Q� 	��Q�      D  , , ���Q� ���R6 ���R6 ���Q� ���Q�      D  , , 	��O  	��O� 	���O� 	���O  	��O       D  , , ���O  ���O� ���O� ���O  ���O       D  , , 	��L� 	��M6 	���M6 	���L� 	��L�      D  , , ���L� ���M6 ���M6 ���L� ���L�      D  , , ���L� ���M6 r��M6 r��L� ���L�      D  , , ���L� ���M6 V��M6 V��L� ���L�      D  , , v���h v���h� w���h� w���h v���h      D  , , v���f� v���gX w���gX w���f� v���f�      D  , , v���nB v���n� w���n� w���nB v���nB      D  , , v���e� v���f w���f w���e� v���e�      D  , , v���p� v���qX w���qX w���p� v���p�      D  , , v���dB v���d� w���d� w���dB v���dB      D  , , v���c v���c� w���c� w���c v���c      D  , , v���m v���m� w���m� w���m v���m      D  , , v���k� v���lX w���lX w���k� v���k�      D  , , v���o� v���p w���p w���o� v���o�      D  , , v���[� v���\6 w���\6 w���[� v���[�      D  , , v���j� v���k w���k w���j� v���j�      D  , , v���Z` v���Z� w���Z� w���Z` v���Z`      D  , , v���Y  v���Y� w���Y� w���Y  v���Y       D  , , v���W� v���Xv w���Xv w���W� v���W�      D  , , v���V� v���W6 w���W6 w���V� v���V�      D  , , v���r v���r� w���r� w���r v���r      D  , , v���U` v���U� w���U� w���U` v���U`      D  , , v���T  v���T� w���T� w���T  v���T       D  , , v���R� v���Sv w���Sv w���R� v���R�      D  , , v���iB v���i� w���i� w���iB v���iB      D  , , v���Q� v���R6 w���R6 w���Q� v���Q�      D  , , v���P` v���P� w���P� w���P` v���P`      D  , , v���O  v���O� w���O� w���O  v���O       D  , , v���M� v���Nv w���Nv w���M� v���M�      D  , , v���L� v���M6 w���M6 w���L� v���L�      D  , , ���iB ���i� :��i� :��iB ���iB      D  , , ���iB ���i� ��i� ��iB ���iB      D  , , l��iB l��i� ��i� ��iB l��iB      D  , , P��iB P��i� ���i� ���iB P��iB      D  , ,  4��iB  4��i�  ���i�  ���iB  4��iB      D  , , #��iB #��i� #���i� #���iB #��iB      D  , , %���iB %���i� &���i� &���iB %���iB      D  , , (���iB (���i� )v��i� )v��iB (���iB      D  , , +���iB +���i� ,Z��i� ,Z��iB +���iB      D  , , .���iB .���i� />��i� />��iB .���iB      D  , , 1���iB 1���i� 2"��i� 2"��iB 1���iB      D  , , 4p��iB 4p��i� 5��i� 5��iB 4p��iB      D  , , 7T��iB 7T��i� 7���i� 7���iB 7T��iB      D  , , :8��iB :8��i� :���i� :���iB :8��iB      D  , , =��iB =��i� =���i� =���iB =��iB      D  , , @ ��iB @ ��i� @���i� @���iB @ ��iB      D  , , B���iB B���i� Cz��i� Cz��iB B���iB      D  , , E���iB E���i� F^��i� F^��iB E���iB      D  , , H���iB H���i� IB��i� IB��iB H���iB      D  , , K���iB K���i� L&��i� L&��iB K���iB      D  , , Nt��iB Nt��i� O
��i� O
��iB Nt��iB      D  , , QX��iB QX��i� Q���i� Q���iB QX��iB      D  , , T<��iB T<��i� T���i� T���iB T<��iB      D  , , W ��iB W ��i� W���i� W���iB W ��iB      D  , , Z��iB Z��i� Z���i� Z���iB Z��iB      D  , , \���iB \���i� ]~��i� ]~��iB \���iB      D  , , _���iB _���i� `b��i� `b��iB _���iB      D  , , b���iB b���i� cF��i� cF��iB b���iB      D  , , e���iB e���i� f*��i� f*��iB e���iB      D  , , hx��iB hx��i� i��i� i��iB hx��iB      D  , , k\��iB k\��i� k���i� k���iB k\��iB      D  , , n@��iB n@��i� n���i� n���iB n@��iB      D  , , q$��iB q$��i� q���i� q���iB q$��iB      D  , , t��iB t��i� t���i� t���iB t��iB      D  , , E���m E���m� F^��m� F^��m E���m      D  , , H���m H���m� IB��m� IB��m H���m      D  , , K���m K���m� L&��m� L&��m K���m      D  , , Nt��m Nt��m� O
��m� O
��m Nt��m      D  , , QX��m QX��m� Q���m� Q���m QX��m      D  , , T<��m T<��m� T���m� T���m T<��m      D  , , W ��m W ��m� W���m� W���m W ��m      D  , , Z��m Z��m� Z���m� Z���m Z��m      D  , , \���m \���m� ]~��m� ]~��m \���m      D  , , E���r E���r� F^��r� F^��r E���r      D  , , H���r H���r� IB��r� IB��r H���r      D  , , K���r K���r� L&��r� L&��r K���r      D  , , E���k� E���lX F^��lX F^��k� E���k�      D  , , H���k� H���lX IB��lX IB��k� H���k�      D  , , K���k� K���lX L&��lX L&��k� K���k�      D  , , Nt��k� Nt��lX O
��lX O
��k� Nt��k�      D  , , QX��k� QX��lX Q���lX Q���k� QX��k�      D  , , T<��k� T<��lX T���lX T���k� T<��k�      D  , , W ��k� W ��lX W���lX W���k� W ��k�      D  , , Z��k� Z��lX Z���lX Z���k� Z��k�      D  , , \���k� \���lX ]~��lX ]~��k� \���k�      D  , , Nt��r Nt��r� O
��r� O
��r Nt��r      D  , , E���o� E���p F^��p F^��o� E���o�      D  , , H���o� H���p IB��p IB��o� H���o�      D  , , K���o� K���p L&��p L&��o� K���o�      D  , , Nt��o� Nt��p O
��p O
��o� Nt��o�      D  , , QX��o� QX��p Q���p Q���o� QX��o�      D  , , T<��o� T<��p T���p T���o� T<��o�      D  , , W ��o� W ��p W���p W���o� W ��o�      D  , , Z��o� Z��p Z���p Z���o� Z��o�      D  , , \���o� \���p ]~��p ]~��o� \���o�      D  , , E���j� E���k F^��k F^��j� E���j�      D  , , H���j� H���k IB��k IB��j� H���j�      D  , , K���j� K���k L&��k L&��j� K���j�      D  , , Nt��j� Nt��k O
��k O
��j� Nt��j�      D  , , QX��j� QX��k Q���k Q���j� QX��j�      D  , , T<��j� T<��k T���k T���j� T<��j�      D  , , W ��j� W ��k W���k W���j� W ��j�      D  , , Z��j� Z��k Z���k Z���j� Z��j�      D  , , \���j� \���k ]~��k ]~��j� \���j�      D  , , QX��r QX��r� Q���r� Q���r QX��r      D  , , T<��r T<��r� T���r� T���r T<��r      D  , , W ��r W ��r� W���r� W���r W ��r      D  , , Z��r Z��r� Z���r� Z���r Z��r      D  , , \���r \���r� ]~��r� ]~��r \���r      D  , , E���p� E���qX F^��qX F^��p� E���p�      D  , , H���p� H���qX IB��qX IB��p� H���p�      D  , , K���p� K���qX L&��qX L&��p� K���p�      D  , , Nt��p� Nt��qX O
��qX O
��p� Nt��p�      D  , , E���nB E���n� F^��n� F^��nB E���nB      D  , , H���nB H���n� IB��n� IB��nB H���nB      D  , , K���nB K���n� L&��n� L&��nB K���nB      D  , , Nt��nB Nt��n� O
��n� O
��nB Nt��nB      D  , , QX��nB QX��n� Q���n� Q���nB QX��nB      D  , , T<��nB T<��n� T���n� T���nB T<��nB      D  , , W ��nB W ��n� W���n� W���nB W ��nB      D  , , Z��nB Z��n� Z���n� Z���nB Z��nB      D  , , \���nB \���n� ]~��n� ]~��nB \���nB      D  , , QX��p� QX��qX Q���qX Q���p� QX��p�      D  , , T<��p� T<��qX T���qX T���p� T<��p�      D  , , W ��p� W ��qX W���qX W���p� W ��p�      D  , , Z��p� Z��qX Z���qX Z���p� Z��p�      D  , , \���p� \���qX ]~��qX ]~��p� \���p�      D  , , q$��m q$��m� q���m� q���m q$��m      D  , , _���j� _���k `b��k `b��j� _���j�      D  , , b���j� b���k cF��k cF��j� b���j�      D  , , e���j� e���k f*��k f*��j� e���j�      D  , , hx��j� hx��k i��k i��j� hx��j�      D  , , k\��j� k\��k k���k k���j� k\��j�      D  , , n@��j� n@��k n���k n���j� n@��j�      D  , , q$��j� q$��k q���k q���j� q$��j�      D  , , t��j� t��k t���k t���j� t��j�      D  , , t��m t��m� t���m� t���m t��m      D  , , _���m _���m� `b��m� `b��m _���m      D  , , b���m b���m� cF��m� cF��m b���m      D  , , e���m e���m� f*��m� f*��m e���m      D  , , hx��m hx��m� i��m� i��m hx��m      D  , , _���r _���r� `b��r� `b��r _���r      D  , , b���r b���r� cF��r� cF��r b���r      D  , , e���r e���r� f*��r� f*��r e���r      D  , , hx��r hx��r� i��r� i��r hx��r      D  , , k\��r k\��r� k���r� k���r k\��r      D  , , n@��r n@��r� n���r� n���r n@��r      D  , , q$��r q$��r� q���r� q���r q$��r      D  , , t��r t��r� t���r� t���r t��r      D  , , _���k� _���lX `b��lX `b��k� _���k�      D  , , b���k� b���lX cF��lX cF��k� b���k�      D  , , _���o� _���p `b��p `b��o� _���o�      D  , , b���o� b���p cF��p cF��o� b���o�      D  , , e���o� e���p f*��p f*��o� e���o�      D  , , hx��o� hx��p i��p i��o� hx��o�      D  , , k\��o� k\��p k���p k���o� k\��o�      D  , , n@��o� n@��p n���p n���o� n@��o�      D  , , q$��o� q$��p q���p q���o� q$��o�      D  , , t��o� t��p t���p t���o� t��o�      D  , , e���k� e���lX f*��lX f*��k� e���k�      D  , , hx��k� hx��lX i��lX i��k� hx��k�      D  , , k\��k� k\��lX k���lX k���k� k\��k�      D  , , _���nB _���n� `b��n� `b��nB _���nB      D  , , b���nB b���n� cF��n� cF��nB b���nB      D  , , e���nB e���n� f*��n� f*��nB e���nB      D  , , hx��nB hx��n� i��n� i��nB hx��nB      D  , , k\��nB k\��n� k���n� k���nB k\��nB      D  , , n@��nB n@��n� n���n� n���nB n@��nB      D  , , q$��nB q$��n� q���n� q���nB q$��nB      D  , , t��nB t��n� t���n� t���nB t��nB      D  , , n@��k� n@��lX n���lX n���k� n@��k�      D  , , q$��k� q$��lX q���lX q���k� q$��k�      D  , , t��k� t��lX t���lX t���k� t��k�      D  , , k\��m k\��m� k���m� k���m k\��m      D  , , n@��m n@��m� n���m� n���m n@��m      D  , , _���p� _���qX `b��qX `b��p� _���p�      D  , , b���p� b���qX cF��qX cF��p� b���p�      D  , , e���p� e���qX f*��qX f*��p� e���p�      D  , , hx��p� hx��qX i��qX i��p� hx��p�      D  , , k\��p� k\��qX k���qX k���p� k\��p�      D  , , n@��p� n@��qX n���qX n���p� n@��p�      D  , , q$��p� q$��qX q���qX q���p� q$��p�      D  , , t��p� t��qX t���qX t���p� t��p�      D  , , +���o� +���p ,Z��p ,Z��o� +���o�      D  , , +���nB +���n� ,Z��n� ,Z��nB +���nB      D  , , +���j� +���k ,Z��k ,Z��j� +���j�      D  , , +���r +���r� ,Z��r� ,Z��r +���r      D  , , +���k� +���lX ,Z��lX ,Z��k� +���k�      D  , , +���m +���m� ,Z��m� ,Z��m +���m      D  , , +���p� +���qX ,Z��qX ,Z��p� +���p�      D  , , P��nB P��n� ���n� ���nB P��nB      D  , ,  4��nB  4��n�  ���n�  ���nB  4��nB      D  , , #��nB #��n� #���n� #���nB #��nB      D  , , %���nB %���n� &���n� &���nB %���nB      D  , , (���nB (���n� )v��n� )v��nB (���nB      D  , , %���o� %���p &���p &���o� %���o�      D  , , ���j� ���k :��k :��j� ���j�      D  , , ���j� ���k ��k ��j� ���j�      D  , , l��j� l��k ��k ��j� l��j�      D  , , P��j� P��k ���k ���j� P��j�      D  , ,  4��j�  4��k  ���k  ���j�  4��j�      D  , , #��j� #��k #���k #���j� #��j�      D  , , %���j� %���k &���k &���j� %���j�      D  , , (���j� (���k )v��k )v��j� (���j�      D  , , (���o� (���p )v��p )v��o� (���o�      D  , , ���r ���r� :��r� :��r ���r      D  , , ���r ���r� ��r� ��r ���r      D  , , l��r l��r� ��r� ��r l��r      D  , , P��r P��r� ���r� ���r P��r      D  , ,  4��r  4��r�  ���r�  ���r  4��r      D  , , #��r #��r� #���r� #���r #��r      D  , , %���r %���r� &���r� &���r %���r      D  , , (���r (���r� )v��r� )v��r (���r      D  , , #��o� #��p #���p #���o� #��o�      D  , , ���k� ���lX :��lX :��k� ���k�      D  , , ���k� ���lX ��lX ��k� ���k�      D  , , l��k� l��lX ��lX ��k� l��k�      D  , , P��k� P��lX ���lX ���k� P��k�      D  , ,  4��k�  4��lX  ���lX  ���k�  4��k�      D  , , #��k� #��lX #���lX #���k� #��k�      D  , , %���k� %���lX &���lX &���k� %���k�      D  , , (���k� (���lX )v��lX )v��k� (���k�      D  , , ���nB ���n� :��n� :��nB ���nB      D  , , ���m ���m� :��m� :��m ���m      D  , , ���m ���m� ��m� ��m ���m      D  , , l��m l��m� ��m� ��m l��m      D  , , P��m P��m� ���m� ���m P��m      D  , ,  4��m  4��m�  ���m�  ���m  4��m      D  , , #��m #��m� #���m� #���m #��m      D  , , %���m %���m� &���m� &���m %���m      D  , , (���m (���m� )v��m� )v��m (���m      D  , , ���nB ���n� ��n� ��nB ���nB      D  , , ���o� ���p :��p :��o� ���o�      D  , , ���o� ���p ��p ��o� ���o�      D  , , l��o� l��p ��p ��o� l��o�      D  , , P��o� P��p ���p ���o� P��o�      D  , ,  4��o�  4��p  ���p  ���o�  4��o�      D  , , ���p� ���qX :��qX :��p� ���p�      D  , , ���p� ���qX ��qX ��p� ���p�      D  , , l��p� l��qX ��qX ��p� l��p�      D  , , P��p� P��qX ���qX ���p� P��p�      D  , ,  4��p�  4��qX  ���qX  ���p�  4��p�      D  , , #��p� #��qX #���qX #���p� #��p�      D  , , %���p� %���qX &���qX &���p� %���p�      D  , , (���p� (���qX )v��qX )v��p� (���p�      D  , , l��nB l��n� ��n� ��nB l��nB      D  , , :8��r :8��r� :���r� :���r :8��r      D  , , =��r =��r� =���r� =���r =��r      D  , , @ ��r @ ��r� @���r� @���r @ ��r      D  , , B���r B���r� Cz��r� Cz��r B���r      D  , , =��nB =��n� =���n� =���nB =��nB      D  , , @ ��nB @ ��n� @���n� @���nB @ ��nB      D  , , B���nB B���n� Cz��n� Cz��nB B���nB      D  , , B���m B���m� Cz��m� Cz��m B���m      D  , , 1���p� 1���qX 2"��qX 2"��p� 1���p�      D  , , 4p��p� 4p��qX 5��qX 5��p� 4p��p�      D  , , 7T��p� 7T��qX 7���qX 7���p� 7T��p�      D  , , .���o� .���p />��p />��o� .���o�      D  , , 1���o� 1���p 2"��p 2"��o� 1���o�      D  , , 4p��o� 4p��p 5��p 5��o� 4p��o�      D  , , .���j� .���k />��k />��j� .���j�      D  , , 1���j� 1���k 2"��k 2"��j� 1���j�      D  , , .���k� .���lX />��lX />��k� .���k�      D  , , 1���k� 1���lX 2"��lX 2"��k� 1���k�      D  , , 4p��k� 4p��lX 5��lX 5��k� 4p��k�      D  , , 7T��k� 7T��lX 7���lX 7���k� 7T��k�      D  , , :8��k� :8��lX :���lX :���k� :8��k�      D  , , =��k� =��lX =���lX =���k� =��k�      D  , , @ ��k� @ ��lX @���lX @���k� @ ��k�      D  , , B���k� B���lX Cz��lX Cz��k� B���k�      D  , , :8��p� :8��qX :���qX :���p� :8��p�      D  , , =��p� =��qX =���qX =���p� =��p�      D  , , @ ��p� @ ��qX @���qX @���p� @ ��p�      D  , , B���p� B���qX Cz��qX Cz��p� B���p�      D  , , .���p� .���qX />��qX />��p� .���p�      D  , , 4p��j� 4p��k 5��k 5��j� 4p��j�      D  , , 7T��j� 7T��k 7���k 7���j� 7T��j�      D  , , :8��j� :8��k :���k :���j� :8��j�      D  , , =��j� =��k =���k =���j� =��j�      D  , , @ ��j� @ ��k @���k @���j� @ ��j�      D  , , B���j� B���k Cz��k Cz��j� B���j�      D  , , 1���nB 1���n� 2"��n� 2"��nB 1���nB      D  , , 4p��nB 4p��n� 5��n� 5��nB 4p��nB      D  , , 7T��nB 7T��n� 7���n� 7���nB 7T��nB      D  , , .���m .���m� />��m� />��m .���m      D  , , 1���m 1���m� 2"��m� 2"��m 1���m      D  , , 4p��m 4p��m� 5��m� 5��m 4p��m      D  , , 7T��m 7T��m� 7���m� 7���m 7T��m      D  , , :8��nB :8��n� :���n� :���nB :8��nB      D  , , 7T��o� 7T��p 7���p 7���o� 7T��o�      D  , , :8��o� :8��p :���p :���o� :8��o�      D  , , =��o� =��p =���p =���o� =��o�      D  , , @ ��o� @ ��p @���p @���o� @ ��o�      D  , , B���o� B���p Cz��p Cz��o� B���o�      D  , , :8��m :8��m� :���m� :���m :8��m      D  , , .���nB .���n� />��n� />��nB .���nB      D  , , =��m =��m� =���m� =���m =��m      D  , , @ ��m @ ��m� @���m� @���m @ ��m      D  , , .���r .���r� />��r� />��r .���r      D  , , 1���r 1���r� 2"��r� 2"��r 1���r      D  , , 4p��r 4p��r� 5��r� 5��r 4p��r      D  , , 7T��r 7T��r� 7���r� 7���r 7T��r      D  , , +���[� +���\6 ,Z��\6 ,Z��[� +���[�      D  , , +���f� +���gX ,Z��gX ,Z��f� +���f�      D  , , +���dB +���d� ,Z��d� ,Z��dB +���dB      D  , , +���Z` +���Z� ,Z��Z� ,Z��Z` +���Z`      D  , , +���Y  +���Y� ,Z��Y� ,Z��Y  +���Y       D  , , +���W� +���Xv ,Z��Xv ,Z��W� +���W�      D  , , +���V� +���W6 ,Z��W6 ,Z��V� +���V�      D  , , +���U` +���U� ,Z��U� ,Z��U` +���U`      D  , , +���c +���c� ,Z��c� ,Z��c +���c      D  , , +���h +���h� ,Z��h� ,Z��h +���h      D  , , +���T  +���T� ,Z��T� ,Z��T  +���T       D  , , +���R� +���Sv ,Z��Sv ,Z��R� +���R�      D  , , +���e� +���f ,Z��f ,Z��e� +���e�      D  , , +���Q� +���R6 ,Z��R6 ,Z��Q� +���Q�      D  , , +���P` +���P� ,Z��P� ,Z��P` +���P`      D  , , +���O  +���O� ,Z��O� ,Z��O  +���O       D  , , +���M� +���Nv ,Z��Nv ,Z��M� +���M�      D  , , +���L� +���M6 ,Z��M6 ,Z��L� +���L�      D  , , >���_� >���`� ?$��`� ?$��_� >���_�      D  , , Ar��_� Ar��`� B��`� B��_� Ar��_�      D  , , DV��_� DV��`� D���`� D���_� DV��_�      D  , , -6��_� -6��`� -���`� -���_� -6��_�      D  , , 0��_� 0��`� 0���`� 0���_� 0��_�      D  , , -6��^� -6��_G -���_G -���^� -6��^�      D  , , 0��^� 0��_G 0���_G 0���^� 0��^�      D  , , 2���^� 2���_G 3���_G 3���^� 2���^�      D  , , 5���^� 5���_G 6x��_G 6x��^� 5���^�      D  , , 8���^� 8���_G 9\��_G 9\��^� 8���^�      D  , , ;���^� ;���_G <@��_G <@��^� ;���^�      D  , , >���^� >���_G ?$��_G ?$��^� >���^�      D  , , Ar��^� Ar��_G B��_G B��^� Ar��^�      D  , , :8��h :8��h� :���h� :���h :8��h      D  , , 2���_� 2���`� 3���`� 3���_� 2���_�      D  , , =��h =��h� =���h� =���h =��h      D  , , 5���_� 5���`� 6x��`� 6x��_� 5���_�      D  , , @ ��h @ ��h� @���h� @���h @ ��h      D  , , DV��^� DV��_G D���_G D���^� DV��^�      D  , , .���dB .���d� />��d� />��dB .���dB      D  , , 8���_� 8���`� 9\��`� 9\��_� 8���_�      D  , , B���h B���h� Cz��h� Cz��h B���h      D  , , 1���dB 1���d� 2"��d� 2"��dB 1���dB      D  , , 4p��dB 4p��d� 5��d� 5��dB 4p��dB      D  , , 7T��dB 7T��d� 7���d� 7���dB 7T��dB      D  , , :8��dB :8��d� :���d� :���dB :8��dB      D  , , =��dB =��d� =���d� =���dB =��dB      D  , , @ ��dB @ ��d� @���d� @���dB @ ��dB      D  , , B���dB B���d� Cz��d� Cz��dB B���dB      D  , , 4p��h 4p��h� 5��h� 5��h 4p��h      D  , , .���h .���h� />��h� />��h .���h      D  , , .���[� .���\6 />��\6 />��[� .���[�      D  , , .���c .���c� />��c� />��c .���c      D  , , 1���c 1���c� 2"��c� 2"��c 1���c      D  , , 4p��c 4p��c� 5��c� 5��c 4p��c      D  , , 7T��c 7T��c� 7���c� 7���c 7T��c      D  , , :8��c :8��c� :���c� :���c :8��c      D  , , =��c =��c� =���c� =���c =��c      D  , , @ ��c @ ��c� @���c� @���c @ ��c      D  , , B���c B���c� Cz��c� Cz��c B���c      D  , , 1���[� 1���\6 2"��\6 2"��[� 1���[�      D  , , 4p��[� 4p��\6 5��\6 5��[� 4p��[�      D  , , .���f� .���gX />��gX />��f� .���f�      D  , , 1���f� 1���gX 2"��gX 2"��f� 1���f�      D  , , 4p��f� 4p��gX 5��gX 5��f� 4p��f�      D  , , 7T��f� 7T��gX 7���gX 7���f� 7T��f�      D  , , :8��f� :8��gX :���gX :���f� :8��f�      D  , , =��f� =��gX =���gX =���f� =��f�      D  , , 7T��[� 7T��\6 7���\6 7���[� 7T��[�      D  , , 1���h 1���h� 2"��h� 2"��h 1���h      D  , , :8��[� :8��\6 :���\6 :���[� :8��[�      D  , , .���e� .���f />��f />��e� .���e�      D  , , 1���e� 1���f 2"��f 2"��e� 1���e�      D  , , =��[� =��\6 =���\6 =���[� =��[�      D  , , @ ��[� @ ��\6 @���\6 @���[� @ ��[�      D  , , B���[� B���\6 Cz��\6 Cz��[� B���[�      D  , , 7T��h 7T��h� 7���h� 7���h 7T��h      D  , , 4p��e� 4p��f 5��f 5��e� 4p��e�      D  , , 7T��e� 7T��f 7���f 7���e� 7T��e�      D  , , :8��e� :8��f :���f :���e� :8��e�      D  , , =��e� =��f =���f =���e� =��e�      D  , , @ ��e� @ ��f @���f @���e� @ ��e�      D  , , B���e� B���f Cz��f Cz��e� B���e�      D  , , @ ��f� @ ��gX @���gX @���f� @ ��f�      D  , , B���f� B���gX Cz��gX Cz��f� B���f�      D  , , ;���_� ;���`� <@��`� <@��_� ;���_�      D  , , ���f� ���gX ��gX ��f� ���f�      D  , , l��f� l��gX ��gX ��f� l��f�      D  , , P��f� P��gX ���gX ���f� P��f�      D  , , #��f� #��gX #���gX #���f� #��f�      D  , , %���f� %���gX &���gX &���f� %���f�      D  , , (���f� (���gX )v��gX )v��f� (���f�      D  , , (���h (���h� )v��h� )v��h (���h      D  , , ���c ���c� :��c� :��c ���c      D  , , ���c ���c� ��c� ��c ���c      D  , , l��c l��c� ��c� ��c l��c      D  , ,  4��f�  4��gX  ���gX  ���f�  4��f�      D  , , P��c P��c� ���c� ���c P��c      D  , ,  4��c  4��c�  ���c�  ���c  4��c      D  , , #��c #��c� #���c� #���c #��c      D  , , %���c %���c� &���c� &���c %���c      D  , , %���h %���h� &���h� &���h %���h      D  , , (���c (���c� )v��c� )v��c (���c      D  , , ���dB ���d� :��d� :��dB ���dB      D  , , ���dB ���d� ��d� ��dB ���dB      D  , , l��dB l��d� ��d� ��dB l��dB      D  , , P��dB P��d� ���d� ���dB P��dB      D  , ,  4��dB  4��d�  ���d�  ���dB  4��dB      D  , , #��dB #��d� #���d� #���dB #��dB      D  , , %���dB %���d� &���d� &���dB %���dB      D  , , (���dB (���d� )v��d� )v��dB (���dB      D  , , ���[� ���\6 :��\6 :��[� ���[�      D  , , ��^� ��_G ���_G ���^� ��^�      D  , , ���^� ���_G ���_G ���^� ���^�      D  , , ���^� ���_G t��_G t��^� ���^�      D  , , ���^� ���_G X��_G X��^� ���^�      D  , , !���^� !���_G "<��_G "<��^� !���^�      D  , , $���^� $���_G % ��_G % ��^� $���^�      D  , , 'n��^� 'n��_G (��_G (��^� 'n��^�      D  , , *R��^� *R��_G *���_G *���^� *R��^�      D  , ,  4��h  4��h�  ���h�  ���h  4��h      D  , , ���e� ���f :��f :��e� ���e�      D  , , ���e� ���f ��f ��e� ���e�      D  , , l��e� l��f ��f ��e� l��e�      D  , , P��e� P��f ���f ���e� P��e�      D  , , ���[� ���\6 ��\6 ��[� ���[�      D  , ,  4��e�  4��f  ���f  ���e�  4��e�      D  , , #��e� #��f #���f #���e� #��e�      D  , , l��[� l��\6 ��\6 ��[� l��[�      D  , , %���e� %���f &���f &���e� %���e�      D  , , (���e� (���f )v��f )v��e� (���e�      D  , , P��[� P��\6 ���\6 ���[� P��[�      D  , ,  4��[�  4��\6  ���\6  ���[�  4��[�      D  , , #��[� #��\6 #���\6 #���[� #��[�      D  , , %���[� %���\6 &���\6 &���[� %���[�      D  , , (���[� (���\6 )v��\6 )v��[� (���[�      D  , , P��h P��h� ���h� ���h P��h      D  , , ��_� ��`� ���`� ���_� ��_�      D  , , ���_� ���`� ���`� ���_� ���_�      D  , , ���_� ���`� t��`� t��_� ���_�      D  , , ���_� ���`� X��`� X��_� ���_�      D  , , !���_� !���`� "<��`� "<��_� !���_�      D  , , $���_� $���`� % ��`� % ��_� $���_�      D  , , 'n��_� 'n��`� (��`� (��_� 'n��_�      D  , , #��h #��h� #���h� #���h #��h      D  , , *R��_� *R��`� *���`� *���_� *R��_�      D  , , l��h l��h� ��h� ��h l��h      D  , , ���h ���h� :��h� :��h ���h      D  , , ���h ���h� ��h� ��h ���h      D  , , ���f� ���gX :��gX :��f� ���f�      D  , , ���Z` ���Z� ��Z� ��Z` ���Z`      D  , , ���Y  ���Y� :��Y� :��Y  ���Y       D  , , ���Y  ���Y� ��Y� ��Y  ���Y       D  , , ���T  ���T� :��T� :��T  ���T       D  , , ���T  ���T� ��T� ��T  ���T       D  , , l��T  l��T� ��T� ��T  l��T       D  , , P��T  P��T� ���T� ���T  P��T       D  , ,  4��T   4��T�  ���T�  ���T   4��T       D  , , #��T  #��T� #���T� #���T  #��T       D  , , %���T  %���T� &���T� &���T  %���T       D  , , (���T  (���T� )v��T� )v��T  (���T       D  , , l��Y  l��Y� ��Y� ��Y  l��Y       D  , , P��Y  P��Y� ���Y� ���Y  P��Y       D  , ,  4��Y   4��Y�  ���Y�  ���Y   4��Y       D  , , #��Y  #��Y� #���Y� #���Y  #��Y       D  , , %���Y  %���Y� &���Y� &���Y  %���Y       D  , , (���Y  (���Y� )v��Y� )v��Y  (���Y       D  , , l��Z` l��Z� ��Z� ��Z` l��Z`      D  , , ���V� ���W6 :��W6 :��V� ���V�      D  , , ���V� ���W6 ��W6 ��V� ���V�      D  , , l��V� l��W6 ��W6 ��V� l��V�      D  , , P��V� P��W6 ���W6 ���V� P��V�      D  , ,  4��V�  4��W6  ���W6  ���V�  4��V�      D  , , ���R� ���Sv :��Sv :��R� ���R�      D  , , ���R� ���Sv ��Sv ��R� ���R�      D  , , l��R� l��Sv ��Sv ��R� l��R�      D  , , P��R� P��Sv ���Sv ���R� P��R�      D  , ,  4��R�  4��Sv  ���Sv  ���R�  4��R�      D  , , #��R� #��Sv #���Sv #���R� #��R�      D  , , %���R� %���Sv &���Sv &���R� %���R�      D  , , (���R� (���Sv )v��Sv )v��R� (���R�      D  , , #��V� #��W6 #���W6 #���V� #��V�      D  , , %���V� %���W6 &���W6 &���V� %���V�      D  , , (���V� (���W6 )v��W6 )v��V� (���V�      D  , , P��Z` P��Z� ���Z� ���Z` P��Z`      D  , ,  4��Z`  4��Z�  ���Z�  ���Z`  4��Z`      D  , , #��Z` #��Z� #���Z� #���Z` #��Z`      D  , , ���W� ���Xv :��Xv :��W� ���W�      D  , , ���W� ���Xv ��Xv ��W� ���W�      D  , , ���U` ���U� :��U� :��U` ���U`      D  , , ���Q� ���R6 :��R6 :��Q� ���Q�      D  , , ���Q� ���R6 ��R6 ��Q� ���Q�      D  , , l��Q� l��R6 ��R6 ��Q� l��Q�      D  , , P��Q� P��R6 ���R6 ���Q� P��Q�      D  , ,  4��Q�  4��R6  ���R6  ���Q�  4��Q�      D  , , #��Q� #��R6 #���R6 #���Q� #��Q�      D  , , %���Q� %���R6 &���R6 &���Q� %���Q�      D  , , (���Q� (���R6 )v��R6 )v��Q� (���Q�      D  , , ���U` ���U� ��U� ��U` ���U`      D  , , ���P` ���P� :��P� :��P` ���P`      D  , , ���P` ���P� ��P� ��P` ���P`      D  , , l��P` l��P� ��P� ��P` l��P`      D  , , P��P` P��P� ���P� ���P` P��P`      D  , ,  4��P`  4��P�  ���P�  ���P`  4��P`      D  , , #��P` #��P� #���P� #���P` #��P`      D  , , %���P` %���P� &���P� &���P` %���P`      D  , , (���P` (���P� )v��P� )v��P` (���P`      D  , , l��U` l��U� ��U� ��U` l��U`      D  , , ���O  ���O� :��O� :��O  ���O       D  , , ���O  ���O� ��O� ��O  ���O       D  , , l��O  l��O� ��O� ��O  l��O       D  , , P��O  P��O� ���O� ���O  P��O       D  , ,  4��O   4��O�  ���O�  ���O   4��O       D  , , #��O  #��O� #���O� #���O  #��O       D  , , %���O  %���O� &���O� &���O  %���O       D  , , (���O  (���O� )v��O� )v��O  (���O       D  , , P��U` P��U� ���U� ���U` P��U`      D  , , ���M� ���Nv :��Nv :��M� ���M�      D  , , ���M� ���Nv ��Nv ��M� ���M�      D  , , l��M� l��Nv ��Nv ��M� l��M�      D  , , P��M� P��Nv ���Nv ���M� P��M�      D  , ,  4��M�  4��Nv  ���Nv  ���M�  4��M�      D  , , #��M� #��Nv #���Nv #���M� #��M�      D  , , %���M� %���Nv &���Nv &���M� %���M�      D  , , (���M� (���Nv )v��Nv )v��M� (���M�      D  , ,  4��U`  4��U�  ���U�  ���U`  4��U`      D  , , #��U` #��U� #���U� #���U` #��U`      D  , , %���U` %���U� &���U� &���U` %���U`      D  , , (���U` (���U� )v��U� )v��U` (���U`      D  , , l��W� l��Xv ��Xv ��W� l��W�      D  , , P��W� P��Xv ���Xv ���W� P��W�      D  , ,  4��W�  4��Xv  ���Xv  ���W�  4��W�      D  , , #��W� #��Xv #���Xv #���W� #��W�      D  , , %���W� %���Xv &���Xv &���W� %���W�      D  , , (���W� (���Xv )v��Xv )v��W� (���W�      D  , , %���Z` %���Z� &���Z� &���Z` %���Z`      D  , , (���Z` (���Z� )v��Z� )v��Z` (���Z`      D  , , ���L� ���M6 :��M6 :��L� ���L�      D  , , ���L� ���M6 ��M6 ��L� ���L�      D  , , l��L� l��M6 ��M6 ��L� l��L�      D  , , P��L� P��M6 ���M6 ���L� P��L�      D  , ,  4��L�  4��M6  ���M6  ���L�  4��L�      D  , , #��L� #��M6 #���M6 #���L� #��L�      D  , , %���L� %���M6 &���M6 &���L� %���L�      D  , , (���L� (���M6 )v��M6 )v��L� (���L�      D  , , ���Z` ���Z� :��Z� :��Z` ���Z`      D  , , 4p��W� 4p��Xv 5��Xv 5��W� 4p��W�      D  , , 7T��W� 7T��Xv 7���Xv 7���W� 7T��W�      D  , , :8��W� :8��Xv :���Xv :���W� :8��W�      D  , , .���V� .���W6 />��W6 />��V� .���V�      D  , , 1���V� 1���W6 2"��W6 2"��V� 1���V�      D  , , 4p��V� 4p��W6 5��W6 5��V� 4p��V�      D  , , 7T��V� 7T��W6 7���W6 7���V� 7T��V�      D  , , :8��V� :8��W6 :���W6 :���V� :8��V�      D  , , =��V� =��W6 =���W6 =���V� =��V�      D  , , .���Q� .���R6 />��R6 />��Q� .���Q�      D  , , 1���Q� 1���R6 2"��R6 2"��Q� 1���Q�      D  , , 4p��Q� 4p��R6 5��R6 5��Q� 4p��Q�      D  , , 7T��Q� 7T��R6 7���R6 7���Q� 7T��Q�      D  , , :8��Q� :8��R6 :���R6 :���Q� :8��Q�      D  , , =��Q� =��R6 =���R6 =���Q� =��Q�      D  , , @ ��Q� @ ��R6 @���R6 @���Q� @ ��Q�      D  , , B���Q� B���R6 Cz��R6 Cz��Q� B���Q�      D  , , @ ��V� @ ��W6 @���W6 @���V� @ ��V�      D  , , B���V� B���W6 Cz��W6 Cz��V� B���V�      D  , , =��W� =��Xv =���Xv =���W� =��W�      D  , , .���T  .���T� />��T� />��T  .���T       D  , , 1���T  1���T� 2"��T� 2"��T  1���T       D  , , 4p��T  4p��T� 5��T� 5��T  4p��T       D  , , 7T��T  7T��T� 7���T� 7���T  7T��T       D  , , :8��T  :8��T� :���T� :���T  :8��T       D  , , =��T  =��T� =���T� =���T  =��T       D  , , .���P` .���P� />��P� />��P` .���P`      D  , , 1���P` 1���P� 2"��P� 2"��P` 1���P`      D  , , 4p��P` 4p��P� 5��P� 5��P` 4p��P`      D  , , 7T��P` 7T��P� 7���P� 7���P` 7T��P`      D  , , :8��P` :8��P� :���P� :���P` :8��P`      D  , , =��P` =��P� =���P� =���P` =��P`      D  , , @ ��P` @ ��P� @���P� @���P` @ ��P`      D  , , B���P` B���P� Cz��P� Cz��P` B���P`      D  , , @ ��T  @ ��T� @���T� @���T  @ ��T       D  , , B���T  B���T� Cz��T� Cz��T  B���T       D  , , @ ��W� @ ��Xv @���Xv @���W� @ ��W�      D  , , B���W� B���Xv Cz��Xv Cz��W� B���W�      D  , , :8��Y  :8��Y� :���Y� :���Y  :8��Y       D  , , =��Y  =��Y� =���Y� =���Y  =��Y       D  , , @ ��Y  @ ��Y� @���Y� @���Y  @ ��Y       D  , , B���Y  B���Y� Cz��Y� Cz��Y  B���Y       D  , , 4p��Z` 4p��Z� 5��Z� 5��Z` 4p��Z`      D  , , .���O  .���O� />��O� />��O  .���O       D  , , 1���O  1���O� 2"��O� 2"��O  1���O       D  , , 4p��O  4p��O� 5��O� 5��O  4p��O       D  , , 7T��O  7T��O� 7���O� 7���O  7T��O       D  , , :8��O  :8��O� :���O� :���O  :8��O       D  , , =��O  =��O� =���O� =���O  =��O       D  , , @ ��O  @ ��O� @���O� @���O  @ ��O       D  , , B���O  B���O� Cz��O� Cz��O  B���O       D  , , 7T��Z` 7T��Z� 7���Z� 7���Z` 7T��Z`      D  , , :8��Z` :8��Z� :���Z� :���Z` :8��Z`      D  , , =��Z` =��Z� =���Z� =���Z` =��Z`      D  , , @ ��Z` @ ��Z� @���Z� @���Z` @ ��Z`      D  , , B���Z` B���Z� Cz��Z� Cz��Z` B���Z`      D  , , .���U` .���U� />��U� />��U` .���U`      D  , , 1���U` 1���U� 2"��U� 2"��U` 1���U`      D  , , 4p��U` 4p��U� 5��U� 5��U` 4p��U`      D  , , 7T��U` 7T��U� 7���U� 7���U` 7T��U`      D  , , .���M� .���Nv />��Nv />��M� .���M�      D  , , 1���M� 1���Nv 2"��Nv 2"��M� 1���M�      D  , , 4p��M� 4p��Nv 5��Nv 5��M� 4p��M�      D  , , 7T��M� 7T��Nv 7���Nv 7���M� 7T��M�      D  , , :8��M� :8��Nv :���Nv :���M� :8��M�      D  , , =��M� =��Nv =���Nv =���M� =��M�      D  , , @ ��M� @ ��Nv @���Nv @���M� @ ��M�      D  , , B���M� B���Nv Cz��Nv Cz��M� B���M�      D  , , :8��U` :8��U� :���U� :���U` :8��U`      D  , , =��U` =��U� =���U� =���U` =��U`      D  , , @ ��U` @ ��U� @���U� @���U` @ ��U`      D  , , B���U` B���U� Cz��U� Cz��U` B���U`      D  , , .���R� .���Sv />��Sv />��R� .���R�      D  , , 1���R� 1���Sv 2"��Sv 2"��R� 1���R�      D  , , 4p��R� 4p��Sv 5��Sv 5��R� 4p��R�      D  , , 7T��R� 7T��Sv 7���Sv 7���R� 7T��R�      D  , , :8��R� :8��Sv :���Sv :���R� :8��R�      D  , , =��R� =��Sv =���Sv =���R� =��R�      D  , , @ ��R� @ ��Sv @���Sv @���R� @ ��R�      D  , , B���R� B���Sv Cz��Sv Cz��R� B���R�      D  , , .���Z` .���Z� />��Z� />��Z` .���Z`      D  , , 1���Z` 1���Z� 2"��Z� 2"��Z` 1���Z`      D  , , .���Y  .���Y� />��Y� />��Y  .���Y       D  , , 1���Y  1���Y� 2"��Y� 2"��Y  1���Y       D  , , 4p��Y  4p��Y� 5��Y� 5��Y  4p��Y       D  , , 7T��Y  7T��Y� 7���Y� 7���Y  7T��Y       D  , , .���W� .���Xv />��Xv />��W� .���W�      D  , , 1���W� 1���Xv 2"��Xv 2"��W� 1���W�      D  , , .���L� .���M6 />��M6 />��L� .���L�      D  , , 1���L� 1���M6 2"��M6 2"��L� 1���L�      D  , , 4p��L� 4p��M6 5��M6 5��L� 4p��L�      D  , , 7T��L� 7T��M6 7���M6 7���L� 7T��L�      D  , , :8��L� :8��M6 :���M6 :���L� :8��L�      D  , , =��L� =��M6 =���M6 =���L� =��L�      D  , , @ ��L� @ ��M6 @���M6 @���L� @ ��L�      D  , , B���L� B���M6 Cz��M6 Cz��L� B���L�      D  , , hx��[� hx��\6 i��\6 i��[� hx��[�      D  , , k\��[� k\��\6 k���\6 k���[� k\��[�      D  , , n@��[� n@��\6 n���\6 n���[� n@��[�      D  , , q$��[� q$��\6 q���\6 q���[� q$��[�      D  , , t��[� t��\6 t���\6 t���[� t��[�      D  , , ^Z��^� ^Z��_G ^���_G ^���^� ^Z��^�      D  , , a>��^� a>��_G a���_G a���^� a>��^�      D  , , d"��^� d"��_G d���_G d���^� d"��^�      D  , , g��^� g��_G g���_G g���^� g��^�      D  , , i���^� i���_G j���_G j���^� i���^�      D  , , l���^� l���_G md��_G md��^� l���^�      D  , , o���^� o���_G pH��_G pH��^� o���^�      D  , , r���^� r���_G s,��_G s,��^� r���^�      D  , , uz��^� uz��_G v��_G v��^� uz��^�      D  , , q$��h q$��h� q���h� q���h q$��h      D  , , _���dB _���d� `b��d� `b��dB _���dB      D  , , b���dB b���d� cF��d� cF��dB b���dB      D  , , e���dB e���d� f*��d� f*��dB e���dB      D  , , hx��dB hx��d� i��d� i��dB hx��dB      D  , , k\��dB k\��d� k���d� k���dB k\��dB      D  , , n@��dB n@��d� n���d� n���dB n@��dB      D  , , q$��dB q$��d� q���d� q���dB q$��dB      D  , , t��dB t��d� t���d� t���dB t��dB      D  , , _���e� _���f `b��f `b��e� _���e�      D  , , b���e� b���f cF��f cF��e� b���e�      D  , , e���e� e���f f*��f f*��e� e���e�      D  , , hx��e� hx��f i��f i��e� hx��e�      D  , , k\��e� k\��f k���f k���e� k\��e�      D  , , n@��e� n@��f n���f n���e� n@��e�      D  , , q$��e� q$��f q���f q���e� q$��e�      D  , , t��e� t��f t���f t���e� t��e�      D  , , ^Z��_� ^Z��`� ^���`� ^���_� ^Z��_�      D  , , a>��_� a>��`� a���`� a���_� a>��_�      D  , , d"��_� d"��`� d���`� d���_� d"��_�      D  , , g��_� g��`� g���`� g���_� g��_�      D  , , i���_� i���`� j���`� j���_� i���_�      D  , , l���_� l���`� md��`� md��_� l���_�      D  , , o���_� o���`� pH��`� pH��_� o���_�      D  , , r���_� r���`� s,��`� s,��_� r���_�      D  , , uz��_� uz��`� v��`� v��_� uz��_�      D  , , _���f� _���gX `b��gX `b��f� _���f�      D  , , b���f� b���gX cF��gX cF��f� b���f�      D  , , e���f� e���gX f*��gX f*��f� e���f�      D  , , _���c _���c� `b��c� `b��c _���c      D  , , b���c b���c� cF��c� cF��c b���c      D  , , e���c e���c� f*��c� f*��c e���c      D  , , hx��c hx��c� i��c� i��c hx��c      D  , , k\��c k\��c� k���c� k���c k\��c      D  , , n@��c n@��c� n���c� n���c n@��c      D  , , q$��c q$��c� q���c� q���c q$��c      D  , , t��c t��c� t���c� t���c t��c      D  , , hx��f� hx��gX i��gX i��f� hx��f�      D  , , k\��f� k\��gX k���gX k���f� k\��f�      D  , , _���h _���h� `b��h� `b��h _���h      D  , , n@��f� n@��gX n���gX n���f� n@��f�      D  , , q$��f� q$��gX q���gX q���f� q$��f�      D  , , t��f� t��gX t���gX t���f� t��f�      D  , , t��h t��h� t���h� t���h t��h      D  , , e���h e���h� f*��h� f*��h e���h      D  , , hx��h hx��h� i��h� i��h hx��h      D  , , k\��h k\��h� k���h� k���h k\��h      D  , , n@��h n@��h� n���h� n���h n@��h      D  , , _���[� _���\6 `b��\6 `b��[� _���[�      D  , , b���[� b���\6 cF��\6 cF��[� b���[�      D  , , e���[� e���\6 f*��\6 f*��[� e���[�      D  , , b���h b���h� cF��h� cF��h b���h      D  , , Z��f� Z��gX Z���gX Z���f� Z��f�      D  , , G:��_� G:��`� G���`� G���_� G:��_�      D  , , J��_� J��`� J���`� J���_� J��_�      D  , , M��_� M��`� M���`� M���_� M��_�      D  , , O���_� O���`� P|��`� P|��_� O���_�      D  , , R���_� R���`� S`��`� S`��_� R���_�      D  , , U���_� U���`� VD��`� VD��_� U���_�      D  , , T<��h T<��h� T���h� T���h T<��h      D  , , X���_� X���`� Y(��`� Y(��_� X���_�      D  , , [v��_� [v��`� \��`� \��_� [v��_�      D  , , W ��e� W ��f W���f W���e� W ��e�      D  , , Z��e� Z��f Z���f Z���e� Z��e�      D  , , \���e� \���f ]~��f ]~��e� \���e�      D  , , E���dB E���d� F^��d� F^��dB E���dB      D  , , H���dB H���d� IB��d� IB��dB H���dB      D  , , K���dB K���d� L&��d� L&��dB K���dB      D  , , W ��h W ��h� W���h� W���h W ��h      D  , , Nt��dB Nt��d� O
��d� O
��dB Nt��dB      D  , , QX��dB QX��d� Q���d� Q���dB QX��dB      D  , , T<��dB T<��d� T���d� T���dB T<��dB      D  , , \���f� \���gX ]~��gX ]~��f� \���f�      D  , , W ��dB W ��d� W���d� W���dB W ��dB      D  , , Z��dB Z��d� Z���d� Z���dB Z��dB      D  , , \���dB \���d� ]~��d� ]~��dB \���dB      D  , , E���c E���c� F^��c� F^��c E���c      D  , , H���c H���c� IB��c� IB��c H���c      D  , , Z��h Z��h� Z���h� Z���h Z��h      D  , , K���c K���c� L&��c� L&��c K���c      D  , , Nt��c Nt��c� O
��c� O
��c Nt��c      D  , , QX��c QX��c� Q���c� Q���c QX��c      D  , , T<��c T<��c� T���c� T���c T<��c      D  , , W ��c W ��c� W���c� W���c W ��c      D  , , Z��c Z��c� Z���c� Z���c Z��c      D  , , \���c \���c� ]~��c� ]~��c \���c      D  , , R���^� R���_G S`��_G S`��^� R���^�      D  , , U���^� U���_G VD��_G VD��^� U���^�      D  , , X���^� X���_G Y(��_G Y(��^� X���^�      D  , , [v��^� [v��_G \��_G \��^� [v��^�      D  , , \���h \���h� ]~��h� ]~��h \���h      D  , , H���h H���h� IB��h� IB��h H���h      D  , , E���h E���h� F^��h� F^��h E���h      D  , , O���^� O���_G P|��_G P|��^� O���^�      D  , , E���f� E���gX F^��gX F^��f� E���f�      D  , , K���h K���h� L&��h� L&��h K���h      D  , , Nt��h Nt��h� O
��h� O
��h Nt��h      D  , , H���f� H���gX IB��gX IB��f� H���f�      D  , , E���e� E���f F^��f F^��e� E���e�      D  , , H���e� H���f IB��f IB��e� H���e�      D  , , K���e� K���f L&��f L&��e� K���e�      D  , , Nt��e� Nt��f O
��f O
��e� Nt��e�      D  , , QX��e� QX��f Q���f Q���e� QX��e�      D  , , T<��e� T<��f T���f T���e� T<��e�      D  , , K���f� K���gX L&��gX L&��f� K���f�      D  , , Nt��f� Nt��gX O
��gX O
��f� Nt��f�      D  , , G:��^� G:��_G G���_G G���^� G:��^�      D  , , J��^� J��_G J���_G J���^� J��^�      D  , , M��^� M��_G M���_G M���^� M��^�      D  , , E���[� E���\6 F^��\6 F^��[� E���[�      D  , , H���[� H���\6 IB��\6 IB��[� H���[�      D  , , K���[� K���\6 L&��\6 L&��[� K���[�      D  , , Nt��[� Nt��\6 O
��\6 O
��[� Nt��[�      D  , , QX��[� QX��\6 Q���\6 Q���[� QX��[�      D  , , T<��[� T<��\6 T���\6 T���[� T<��[�      D  , , W ��[� W ��\6 W���\6 W���[� W ��[�      D  , , Z��[� Z��\6 Z���\6 Z���[� Z��[�      D  , , \���[� \���\6 ]~��\6 ]~��[� \���[�      D  , , QX��f� QX��gX Q���gX Q���f� QX��f�      D  , , T<��f� T<��gX T���gX T���f� T<��f�      D  , , QX��h QX��h� Q���h� Q���h QX��h      D  , , W ��f� W ��gX W���gX W���f� W ��f�      D  , , QX��Z` QX��Z� Q���Z� Q���Z` QX��Z`      D  , , QX��P` QX��P� Q���P� Q���P` QX��P`      D  , , QX��R� QX��Sv Q���Sv Q���R� QX��R�      D  , , QX��W� QX��Xv Q���Xv Q���W� QX��W�      D  , , QX��O  QX��O� Q���O� Q���O  QX��O       D  , , QX��T  QX��T� Q���T� Q���T  QX��T       D  , , QX��M� QX��Nv Q���Nv Q���M� QX��M�      D  , , QX��U` QX��U� Q���U� Q���U` QX��U`      D  , , QX��Y  QX��Y� Q���Y� Q���Y  QX��Y       D  , , QX��V� QX��W6 Q���W6 Q���V� QX��V�      D  , , QX��L� QX��M6 Q���M6 Q���L� QX��L�      D  , , QX��Q� QX��R6 Q���R6 Q���Q� QX��Q�      D  , , T<��W� T<��Xv T���Xv T���W� T<��W�      D  , , W ��Z` W ��Z� W���Z� W���Z` W ��Z`      D  , , W ��V� W ��W6 W���W6 W���V� W ��V�      D  , , W ��W� W ��Xv W���Xv W���W� W ��W�      D  , , Z��W� Z��Xv Z���Xv Z���W� Z��W�      D  , , \���W� \���Xv ]~��Xv ]~��W� \���W�      D  , , Z��Z` Z��Z� Z���Z� Z���Z` Z��Z`      D  , , T<��T  T<��T� T���T� T���T  T<��T       D  , , \���U` \���U� ]~��U� ]~��U` \���U`      D  , , W ��T  W ��T� W���T� W���T  W ��T       D  , , Z��T  Z��T� Z���T� Z���T  Z��T       D  , , \���T  \���T� ]~��T� ]~��T  \���T       D  , , Z��V� Z��W6 Z���W6 Z���V� Z��V�      D  , , \���Z` \���Z� ]~��Z� ]~��Z` \���Z`      D  , , T<��U` T<��U� T���U� T���U` T<��U`      D  , , W ��U` W ��U� W���U� W���U` W ��U`      D  , , \���V� \���W6 ]~��W6 ]~��V� \���V�      D  , , T<��Y  T<��Y� T���Y� T���Y  T<��Y       D  , , W ��Y  W ��Y� W���Y� W���Y  W ��Y       D  , , Z��Y  Z��Y� Z���Y� Z���Y  Z��Y       D  , , \���Y  \���Y� ]~��Y� ]~��Y  \���Y       D  , , T<��V� T<��W6 T���W6 T���V� T<��V�      D  , , Z��U` Z��U� Z���U� Z���U` Z��U`      D  , , T<��Z` T<��Z� T���Z� T���Z` T<��Z`      D  , , H���W� H���Xv IB��Xv IB��W� H���W�      D  , , E���U` E���U� F^��U� F^��U` E���U`      D  , , H���U` H���U� IB��U� IB��U` H���U`      D  , , K���U` K���U� L&��U� L&��U` K���U`      D  , , Nt��U` Nt��U� O
��U� O
��U` Nt��U`      D  , , K���W� K���Xv L&��Xv L&��W� K���W�      D  , , E���T  E���T� F^��T� F^��T  E���T       D  , , H���T  H���T� IB��T� IB��T  H���T       D  , , E���Y  E���Y� F^��Y� F^��Y  E���Y       D  , , H���Y  H���Y� IB��Y� IB��Y  H���Y       D  , , K���Y  K���Y� L&��Y� L&��Y  K���Y       D  , , Nt��Y  Nt��Y� O
��Y� O
��Y  Nt��Y       D  , , K���T  K���T� L&��T� L&��T  K���T       D  , , Nt��T  Nt��T� O
��T� O
��T  Nt��T       D  , , Nt��W� Nt��Xv O
��Xv O
��W� Nt��W�      D  , , H���Z` H���Z� IB��Z� IB��Z` H���Z`      D  , , K���Z` K���Z� L&��Z� L&��Z` K���Z`      D  , , E���V� E���W6 F^��W6 F^��V� E���V�      D  , , H���V� H���W6 IB��W6 IB��V� H���V�      D  , , K���V� K���W6 L&��W6 L&��V� K���V�      D  , , Nt��V� Nt��W6 O
��W6 O
��V� Nt��V�      D  , , Nt��Z` Nt��Z� O
��Z� O
��Z` Nt��Z`      D  , , E���Z` E���Z� F^��Z� F^��Z` E���Z`      D  , , E���W� E���Xv F^��Xv F^��W� E���W�      D  , , E���M� E���Nv F^��Nv F^��M� E���M�      D  , , H���M� H���Nv IB��Nv IB��M� H���M�      D  , , K���M� K���Nv L&��Nv L&��M� K���M�      D  , , Nt��M� Nt��Nv O
��Nv O
��M� Nt��M�      D  , , Nt��O  Nt��O� O
��O� O
��O  Nt��O       D  , , Nt��R� Nt��Sv O
��Sv O
��R� Nt��R�      D  , , E���P` E���P� F^��P� F^��P` E���P`      D  , , H���P` H���P� IB��P� IB��P` H���P`      D  , , K���P` K���P� L&��P� L&��P` K���P`      D  , , E���Q� E���R6 F^��R6 F^��Q� E���Q�      D  , , H���Q� H���R6 IB��R6 IB��Q� H���Q�      D  , , K���Q� K���R6 L&��R6 L&��Q� K���Q�      D  , , Nt��Q� Nt��R6 O
��R6 O
��Q� Nt��Q�      D  , , Nt��P` Nt��P� O
��P� O
��P` Nt��P`      D  , , E���R� E���Sv F^��Sv F^��R� E���R�      D  , , H���R� H���Sv IB��Sv IB��R� H���R�      D  , , K���R� K���Sv L&��Sv L&��R� K���R�      D  , , E���O  E���O� F^��O� F^��O  E���O       D  , , E���L� E���M6 F^��M6 F^��L� E���L�      D  , , H���L� H���M6 IB��M6 IB��L� H���L�      D  , , K���L� K���M6 L&��M6 L&��L� K���L�      D  , , Nt��L� Nt��M6 O
��M6 O
��L� Nt��L�      D  , , H���O  H���O� IB��O� IB��O  H���O       D  , , K���O  K���O� L&��O� L&��O  K���O       D  , , Z��O  Z��O� Z���O� Z���O  Z��O       D  , , T<��M� T<��Nv T���Nv T���M� T<��M�      D  , , W ��M� W ��Nv W���Nv W���M� W ��M�      D  , , Z��M� Z��Nv Z���Nv Z���M� Z��M�      D  , , \���M� \���Nv ]~��Nv ]~��M� \���M�      D  , , \���O  \���O� ]~��O� ]~��O  \���O       D  , , \���R� \���Sv ]~��Sv ]~��R� \���R�      D  , , \���Q� \���R6 ]~��R6 ]~��Q� \���Q�      D  , , T<��Q� T<��R6 T���R6 T���Q� T<��Q�      D  , , W ��Q� W ��R6 W���R6 W���Q� W ��Q�      D  , , Z��Q� Z��R6 Z���R6 Z���Q� Z��Q�      D  , , T<��P` T<��P� T���P� T���P` T<��P`      D  , , W ��P` W ��P� W���P� W���P` W ��P`      D  , , Z��P` Z��P� Z���P� Z���P` Z��P`      D  , , \���P` \���P� ]~��P� ]~��P` \���P`      D  , , T<��R� T<��Sv T���Sv T���R� T<��R�      D  , , W ��R� W ��Sv W���Sv W���R� W ��R�      D  , , Z��R� Z��Sv Z���Sv Z���R� Z��R�      D  , , T<��O  T<��O� T���O� T���O  T<��O       D  , , T<��L� T<��M6 T���M6 T���L� T<��L�      D  , , W ��L� W ��M6 W���M6 W���L� W ��L�      D  , , Z��L� Z��M6 Z���M6 Z���L� Z��L�      D  , , \���L� \���M6 ]~��M6 ]~��L� \���L�      D  , , W ��O  W ��O� W���O� W���O  W ��O       D  , , _���Q� _���R6 `b��R6 `b��Q� _���Q�      D  , , b���Q� b���R6 cF��R6 cF��Q� b���Q�      D  , , e���Q� e���R6 f*��R6 f*��Q� e���Q�      D  , , hx��Q� hx��R6 i��R6 i��Q� hx��Q�      D  , , k\��Q� k\��R6 k���R6 k���Q� k\��Q�      D  , , n@��Q� n@��R6 n���R6 n���Q� n@��Q�      D  , , _���O  _���O� `b��O� `b��O  _���O       D  , , b���O  b���O� cF��O� cF��O  b���O       D  , , e���O  e���O� f*��O� f*��O  e���O       D  , , hx��O  hx��O� i��O� i��O  hx��O       D  , , k\��O  k\��O� k���O� k���O  k\��O       D  , , n@��O  n@��O� n���O� n���O  n@��O       D  , , q$��O  q$��O� q���O� q���O  q$��O       D  , , t��O  t��O� t���O� t���O  t��O       D  , , q$��Q� q$��R6 q���R6 q���Q� q$��Q�      D  , , t��Q� t��R6 t���R6 t���Q� t��Q�      D  , , k\��R� k\��Sv k���Sv k���R� k\��R�      D  , , _���Y  _���Y� `b��Y� `b��Y  _���Y       D  , , _���W� _���Xv `b��Xv `b��W� _���W�      D  , , b���W� b���Xv cF��Xv cF��W� b���W�      D  , , e���W� e���Xv f*��Xv f*��W� e���W�      D  , , hx��W� hx��Xv i��Xv i��W� hx��W�      D  , , k\��W� k\��Xv k���Xv k���W� k\��W�      D  , , n@��W� n@��Xv n���Xv n���W� n@��W�      D  , , q$��W� q$��Xv q���Xv q���W� q$��W�      D  , , t��W� t��Xv t���Xv t���W� t��W�      D  , , b���Y  b���Y� cF��Y� cF��Y  b���Y       D  , , e���Y  e���Y� f*��Y� f*��Y  e���Y       D  , , hx��Y  hx��Y� i��Y� i��Y  hx��Y       D  , , k\��Y  k\��Y� k���Y� k���Y  k\��Y       D  , , n@��Y  n@��Y� n���Y� n���Y  n@��Y       D  , , q$��Y  q$��Y� q���Y� q���Y  q$��Y       D  , , t��Y  t��Y� t���Y� t���Y  t��Y       D  , , n@��R� n@��Sv n���Sv n���R� n@��R�      D  , , q$��R� q$��Sv q���Sv q���R� q$��R�      D  , , t��R� t��Sv t���Sv t���R� t��R�      D  , , k\��U` k\��U� k���U� k���U` k\��U`      D  , , n@��U` n@��U� n���U� n���U` n@��U`      D  , , q$��U` q$��U� q���U� q���U` q$��U`      D  , , t��U` t��U� t���U� t���U` t��U`      D  , , _���V� _���W6 `b��W6 `b��V� _���V�      D  , , _���M� _���Nv `b��Nv `b��M� _���M�      D  , , b���M� b���Nv cF��Nv cF��M� b���M�      D  , , e���M� e���Nv f*��Nv f*��M� e���M�      D  , , hx��M� hx��Nv i��Nv i��M� hx��M�      D  , , k\��M� k\��Nv k���Nv k���M� k\��M�      D  , , n@��M� n@��Nv n���Nv n���M� n@��M�      D  , , q$��M� q$��Nv q���Nv q���M� q$��M�      D  , , t��M� t��Nv t���Nv t���M� t��M�      D  , , b���V� b���W6 cF��W6 cF��V� b���V�      D  , , e���V� e���W6 f*��W6 f*��V� e���V�      D  , , hx��V� hx��W6 i��W6 i��V� hx��V�      D  , , k\��V� k\��W6 k���W6 k���V� k\��V�      D  , , n@��V� n@��W6 n���W6 n���V� n@��V�      D  , , _���T  _���T� `b��T� `b��T  _���T       D  , , b���T  b���T� cF��T� cF��T  b���T       D  , , e���T  e���T� f*��T� f*��T  e���T       D  , , _���Z` _���Z� `b��Z� `b��Z` _���Z`      D  , , b���Z` b���Z� cF��Z� cF��Z` b���Z`      D  , , _���P` _���P� `b��P� `b��P` _���P`      D  , , b���P` b���P� cF��P� cF��P` b���P`      D  , , e���P` e���P� f*��P� f*��P` e���P`      D  , , hx��P` hx��P� i��P� i��P` hx��P`      D  , , k\��P` k\��P� k���P� k���P` k\��P`      D  , , n@��P` n@��P� n���P� n���P` n@��P`      D  , , q$��P` q$��P� q���P� q���P` q$��P`      D  , , t��P` t��P� t���P� t���P` t��P`      D  , , e���Z` e���Z� f*��Z� f*��Z` e���Z`      D  , , hx��Z` hx��Z� i��Z� i��Z` hx��Z`      D  , , k\��Z` k\��Z� k���Z� k���Z` k\��Z`      D  , , n@��Z` n@��Z� n���Z� n���Z` n@��Z`      D  , , q$��Z` q$��Z� q���Z� q���Z` q$��Z`      D  , , t��Z` t��Z� t���Z� t���Z` t��Z`      D  , , hx��T  hx��T� i��T� i��T  hx��T       D  , , k\��T  k\��T� k���T� k���T  k\��T       D  , , n@��T  n@��T� n���T� n���T  n@��T       D  , , q$��T  q$��T� q���T� q���T  q$��T       D  , , t��T  t��T� t���T� t���T  t��T       D  , , q$��V� q$��W6 q���W6 q���V� q$��V�      D  , , t��V� t��W6 t���W6 t���V� t��V�      D  , , _���U` _���U� `b��U� `b��U` _���U`      D  , , b���U` b���U� cF��U� cF��U` b���U`      D  , , e���U` e���U� f*��U� f*��U` e���U`      D  , , hx��U` hx��U� i��U� i��U` hx��U`      D  , , _���R� _���Sv `b��Sv `b��R� _���R�      D  , , b���R� b���Sv cF��Sv cF��R� b���R�      D  , , e���R� e���Sv f*��Sv f*��R� e���R�      D  , , _���L� _���M6 `b��M6 `b��L� _���L�      D  , , b���L� b���M6 cF��M6 cF��L� b���L�      D  , , e���L� e���M6 f*��M6 f*��L� e���L�      D  , , hx��L� hx��M6 i��M6 i��L� hx��L�      D  , , k\��L� k\��M6 k���M6 k���L� k\��L�      D  , , n@��L� n@��M6 n���M6 n���L� n@��L�      D  , , q$��L� q$��M6 q���M6 q���L� q$��L�      D  , , t��L� t��M6 t���M6 t���L� t��L�      D  , , hx��R� hx��Sv i��Sv i��R� hx��R�      D  , , y���iB y���i� zf��i� zf��iB y���iB      D  , , |���iB |���i� }J��i� }J��iB |���iB      D  , , ���iB ���i� �.��i� �.��iB ���iB      D  , , �|��iB �|��i� ���i� ���iB �|��iB      D  , , �`��iB �`��i� ����i� ����iB �`��iB      D  , , �D��iB �D��i� ����i� ����iB �D��iB      D  , , �(��iB �(��i� ����i� ����iB �(��iB      D  , , ���iB ���i� ����i� ����iB ���iB      D  , , ����iB ����i� ����i� ����iB ����iB      D  , , ����iB ����i� �j��i� �j��iB ����iB      D  , , ����iB ����i� �N��i� �N��iB ����iB      D  , , ����iB ����i� �2��i� �2��iB ����iB      D  , , ����iB ����i� ���i� ���iB ����iB      D  , , �d��iB �d��i� ����i� ����iB �d��iB      D  , , �H��iB �H��i� ����i� ����iB �H��iB      D  , , �,��iB �,��i� ����i� ����iB �,��iB      D  , , ���iB ���i� ����i� ����iB ���iB      D  , , ����iB ����i� ����i� ����iB ����iB      D  , , ����iB ����i� �n��i� �n��iB ����iB      D  , , ����iB ����i� �R��i� �R��iB ����iB      D  , , ����iB ����i� �6��i� �6��iB ����iB      D  , , ����iB ����i� ���i� ���iB ����iB      D  , , �h��iB �h��i� ����i� ����iB �h��iB      D  , , �L��iB �L��i� ����i� ����iB �L��iB      D  , , �0��iB �0��i� ����i� ����iB �0��iB      D  , , ���iB ���i� ª��i� ª��iB ���iB      D  , , ����iB ����i� Ŏ��i� Ŏ��iB ����iB      D  , , ����iB ����i� �r��i� �r��iB ����iB      D  , , ����iB ����i� �V��i� �V��iB ����iB      D  , , ͤ��iB ͤ��i� �:��i� �:��iB ͤ��iB      D  , , ���ij ���j  Ӟ��j  Ӟ��ij ���ij      D  , , �m��ij �m��j  ���j  ���ij �m��ij      D  , , ����i) ����i� �}��i� �}��i) ����i)      D  , , ����r ����r� ����r� ����r ����r      D  , , ����r ����r� �n��r� �n��r ����r      D  , , ����r ����r� �R��r� �R��r ����r      D  , , ����r ����r� �6��r� �6��r ����r      D  , , ����r ����r� ���r� ���r ����r      D  , , �h��r �h��r� ����r� ����r �h��r      D  , , �L��r �L��r� ����r� ����r �L��r      D  , , �0��r �0��r� ����r� ����r �0��r      D  , , ���r ���r� ª��r� ª��r ���r      D  , , ����r ����r� Ŏ��r� Ŏ��r ����r      D  , , ����r ����r� �r��r� �r��r ����r      D  , , ����r ����r� �V��r� �V��r ����r      D  , , ͤ��r ͤ��r� �:��r� �:��r ͤ��r      D  , , ����k� ����lX ����lX ����k� ����k�      D  , , ����k� ����lX �n��lX �n��k� ����k�      D  , , ����k� ����lX �R��lX �R��k� ����k�      D  , , ����k� ����lX �6��lX �6��k� ����k�      D  , , ����k� ����lX ���lX ���k� ����k�      D  , , �h��k� �h��lX ����lX ����k� �h��k�      D  , , �L��k� �L��lX ����lX ����k� �L��k�      D  , , �0��k� �0��lX ����lX ����k� �0��k�      D  , , ���k� ���lX ª��lX ª��k� ���k�      D  , , ����k� ����lX Ŏ��lX Ŏ��k� ����k�      D  , , ����k� ����lX �r��lX �r��k� ����k�      D  , , ����k� ����lX �V��lX �V��k� ����k�      D  , , ͤ��k� ͤ��lX �:��lX �:��k� ͤ��k�      D  , , ����j� ����k ����k ����j� ����j�      D  , , ����j� ����k �n��k �n��j� ����j�      D  , , ����j� ����k �R��k �R��j� ����j�      D  , , ����j� ����k �6��k �6��j� ����j�      D  , , ����j� ����k ���k ���j� ����j�      D  , , �h��j� �h��k ����k ����j� �h��j�      D  , , �L��j� �L��k ����k ����j� �L��j�      D  , , �0��j� �0��k ����k ����j� �0��j�      D  , , ���j� ���k ª��k ª��j� ���j�      D  , , ����j� ����k Ŏ��k Ŏ��j� ����j�      D  , , ����j� ����k �r��k �r��j� ����j�      D  , , ����j� ����k �V��k �V��j� ����j�      D  , , ͤ��j� ͤ��k �:��k �:��j� ͤ��j�      D  , , ����p� ����qX ����qX ����p� ����p�      D  , , ����p� ����qX �n��qX �n��p� ����p�      D  , , ����p� ����qX �R��qX �R��p� ����p�      D  , , ����p� ����qX �6��qX �6��p� ����p�      D  , , ����p� ����qX ���qX ���p� ����p�      D  , , �h��p� �h��qX ����qX ����p� �h��p�      D  , , �L��p� �L��qX ����qX ����p� �L��p�      D  , , �0��p� �0��qX ����qX ����p� �0��p�      D  , , ���p� ���qX ª��qX ª��p� ���p�      D  , , ����p� ����qX Ŏ��qX Ŏ��p� ����p�      D  , , ����p� ����qX �r��qX �r��p� ����p�      D  , , ����p� ����qX �V��qX �V��p� ����p�      D  , , ����o� ����p ����p ����o� ����o�      D  , , ����o� ����p �n��p �n��o� ����o�      D  , , ����o� ����p �R��p �R��o� ����o�      D  , , ����o� ����p �6��p �6��o� ����o�      D  , , ����o� ����p ���p ���o� ����o�      D  , , �h��o� �h��p ����p ����o� �h��o�      D  , , �L��o� �L��p ����p ����o� �L��o�      D  , , �0��o� �0��p ����p ����o� �0��o�      D  , , ���o� ���p ª��p ª��o� ���o�      D  , , ����o� ����p Ŏ��p Ŏ��o� ����o�      D  , , ����o� ����p �r��p �r��o� ����o�      D  , , ����o� ����p �V��p �V��o� ����o�      D  , , ͤ��o� ͤ��p �:��p �:��o� ͤ��o�      D  , , �0��m �0��m� ����m� ����m �0��m      D  , , ���m ���m� ª��m� ª��m ���m      D  , , ����m ����m� Ŏ��m� Ŏ��m ����m      D  , , ����m ����m� �r��m� �r��m ����m      D  , , ����m ����m� �V��m� �V��m ����m      D  , , ͤ��m ͤ��m� �:��m� �:��m ͤ��m      D  , , ͤ��p� ͤ��qX �:��qX �:��p� ͤ��p�      D  , , ����nB ����n� ����n� ����nB ����nB      D  , , ����nB ����n� �n��n� �n��nB ����nB      D  , , ����nB ����n� �R��n� �R��nB ����nB      D  , , ����m ����m� ����m� ����m ����m      D  , , ����m ����m� �n��m� �n��m ����m      D  , , ����m ����m� �R��m� �R��m ����m      D  , , ����m ����m� �6��m� �6��m ����m      D  , , ����m ����m� ���m� ���m ����m      D  , , �h��m �h��m� ����m� ����m �h��m      D  , , �L��m �L��m� ����m� ����m �L��m      D  , , ����nB ����n� �6��n� �6��nB ����nB      D  , , ����nB ����n� ���n� ���nB ����nB      D  , , �h��nB �h��n� ����n� ����nB �h��nB      D  , , �L��nB �L��n� ����n� ����nB �L��nB      D  , , �0��nB �0��n� ����n� ����nB �0��nB      D  , , ���nB ���n� ª��n� ª��nB ���nB      D  , , ����nB ����n� Ŏ��n� Ŏ��nB ����nB      D  , , ����nB ����n� �r��n� �r��nB ����nB      D  , , ����nB ����n� �V��n� �V��nB ����nB      D  , , ͤ��nB ͤ��n� �:��n� �:��nB ͤ��nB      D  , , �D��j� �D��k ����k ����j� �D��j�      D  , , �(��j� �(��k ����k ����j� �(��j�      D  , , ���j� ���k ����k ����j� ���j�      D  , , ���o� ���p ����p ����o� ���o�      D  , , |���j� |���k }J��k }J��j� |���j�      D  , , y���p� y���qX zf��qX zf��p� y���p�      D  , , |���p� |���qX }J��qX }J��p� |���p�      D  , , ���j� ���k �.��k �.��j� ���j�      D  , , y���nB y���n� zf��n� zf��nB y���nB      D  , , |���nB |���n� }J��n� }J��nB |���nB      D  , , ���nB ���n� �.��n� �.��nB ���nB      D  , , �|��nB �|��n� ���n� ���nB �|��nB      D  , , �`��nB �`��n� ����n� ����nB �`��nB      D  , , y���r y���r� zf��r� zf��r y���r      D  , , |���r |���r� }J��r� }J��r |���r      D  , , ���r ���r� �.��r� �.��r ���r      D  , , �|��r �|��r� ���r� ���r �|��r      D  , , �`��r �`��r� ����r� ����r �`��r      D  , , �D��r �D��r� ����r� ����r �D��r      D  , , ���p� ���qX �.��qX �.��p� ���p�      D  , , y���o� y���p zf��p zf��o� y���o�      D  , , |���o� |���p }J��p }J��o� |���o�      D  , , ���o� ���p �.��p �.��o� ���o�      D  , , �|��o� �|��p ���p ���o� �|��o�      D  , , �`��o� �`��p ����p ����o� �`��o�      D  , , �D��o� �D��p ����p ����o� �D��o�      D  , , �(��o� �(��p ����p ����o� �(��o�      D  , , �|��p� �|��qX ���qX ���p� �|��p�      D  , , �`��p� �`��qX ����qX ����p� �`��p�      D  , , �D��p� �D��qX ����qX ����p� �D��p�      D  , , �(��p� �(��qX ����qX ����p� �(��p�      D  , , ���p� ���qX ����qX ����p� ���p�      D  , , �(��r �(��r� ����r� ����r �(��r      D  , , ���r ���r� ����r� ����r ���r      D  , , �D��nB �D��n� ����n� ����nB �D��nB      D  , , �(��nB �(��n� ����n� ����nB �(��nB      D  , , ���nB ���n� ����n� ����nB ���nB      D  , , y���k� y���lX zf��lX zf��k� y���k�      D  , , |���k� |���lX }J��lX }J��k� |���k�      D  , , y���m y���m� zf��m� zf��m y���m      D  , , |���m |���m� }J��m� }J��m |���m      D  , , y���j� y���k zf��k zf��j� y���j�      D  , , ���m ���m� �.��m� �.��m ���m      D  , , �|��m �|��m� ���m� ���m �|��m      D  , , �`��m �`��m� ����m� ����m �`��m      D  , , �D��m �D��m� ����m� ����m �D��m      D  , , �(��m �(��m� ����m� ����m �(��m      D  , , ���m ���m� ����m� ����m ���m      D  , , ���k� ���lX �.��lX �.��k� ���k�      D  , , �|��k� �|��lX ���lX ���k� �|��k�      D  , , �`��k� �`��lX ����lX ����k� �`��k�      D  , , �D��k� �D��lX ����lX ����k� �D��k�      D  , , �(��k� �(��lX ����lX ����k� �(��k�      D  , , ���k� ���lX ����lX ����k� ���k�      D  , , �|��j� �|��k ���k ���j� �|��j�      D  , , �`��j� �`��k ����k ����j� �`��j�      D  , , ����o� ����p �2��p �2��o� ����o�      D  , , ����o� ����p ���p ���o� ����o�      D  , , ���p� ���qX ����qX ����p� ���p�      D  , , �d��o� �d��p ����p ����o� �d��o�      D  , , �H��o� �H��p ����p ����o� �H��o�      D  , , �,��o� �,��p ����p ����o� �,��o�      D  , , ���o� ���p ����p ����o� ���o�      D  , , ����p� ����qX ����qX ����p� ����p�      D  , , ����p� ����qX �j��qX �j��p� ����p�      D  , , ����p� ����qX �N��qX �N��p� ����p�      D  , , ����p� ����qX �2��qX �2��p� ����p�      D  , , �H��j� �H��k ����k ����j� �H��j�      D  , , �,��j� �,��k ����k ����j� �,��j�      D  , , ���j� ���k ����k ����j� ���j�      D  , , ����j� ����k �j��k �j��j� ����j�      D  , , ����j� ����k �N��k �N��j� ����j�      D  , , ����nB ����n� ����n� ����nB ����nB      D  , , ����nB ����n� �j��n� �j��nB ����nB      D  , , ����nB ����n� �N��n� �N��nB ����nB      D  , , ����nB ����n� �2��n� �2��nB ����nB      D  , , ����nB ����n� ���n� ���nB ����nB      D  , , �d��nB �d��n� ����n� ����nB �d��nB      D  , , �H��nB �H��n� ����n� ����nB �H��nB      D  , , �,��nB �,��n� ����n� ����nB �,��nB      D  , , ���nB ���n� ����n� ����nB ���nB      D  , , ����p� ����qX ���qX ���p� ����p�      D  , , ����j� ����k �2��k �2��j� ����j�      D  , , ����j� ����k ���k ���j� ����j�      D  , , �d��j� �d��k ����k ����j� �d��j�      D  , , ����j� ����k ����k ����j� ����j�      D  , , ����o� ����p ����p ����o� ����o�      D  , , ����o� ����p �j��p �j��o� ����o�      D  , , ����o� ����p �N��p �N��o� ����o�      D  , , �d��p� �d��qX ����qX ����p� �d��p�      D  , , �H��p� �H��qX ����qX ����p� �H��p�      D  , , �,��p� �,��qX ����qX ����p� �,��p�      D  , , ����r ����r� ����r� ����r ����r      D  , , ����m ����m� ����m� ����m ����m      D  , , ����m ����m� �j��m� �j��m ����m      D  , , ����m ����m� �N��m� �N��m ����m      D  , , ����m ����m� �2��m� �2��m ����m      D  , , ����m ����m� ���m� ���m ����m      D  , , �d��m �d��m� ����m� ����m �d��m      D  , , �H��m �H��m� ����m� ����m �H��m      D  , , �,��m �,��m� ����m� ����m �,��m      D  , , ���m ���m� ����m� ����m ���m      D  , , ����r ����r� �j��r� �j��r ����r      D  , , ����r ����r� �N��r� �N��r ����r      D  , , ����r ����r� �2��r� �2��r ����r      D  , , ����r ����r� ���r� ���r ����r      D  , , �d��r �d��r� ����r� ����r �d��r      D  , , �H��r �H��r� ����r� ����r �H��r      D  , , ����k� ����lX ����lX ����k� ����k�      D  , , ����k� ����lX �j��lX �j��k� ����k�      D  , , ����k� ����lX �N��lX �N��k� ����k�      D  , , ����k� ����lX �2��lX �2��k� ����k�      D  , , ����k� ����lX ���lX ���k� ����k�      D  , , �d��k� �d��lX ����lX ����k� �d��k�      D  , , �H��k� �H��lX ����lX ����k� �H��k�      D  , , �,��k� �,��lX ����lX ����k� �,��k�      D  , , ���k� ���lX ����lX ����k� ���k�      D  , , �,��r �,��r� ����r� ����r �,��r      D  , , ���r ���r� ����r� ����r ���r      D  , , �b��_� �b��`� ����`� ����_� �b��_�      D  , , �F��_� �F��`� ����`� ����_� �F��_�      D  , , �*��_� �*��`� ����`� ����_� �*��_�      D  , , ���f� ���gX ����gX ����f� ���f�      D  , , �d��h �d��h� ����h� ����h �d��h      D  , , �H��h �H��h� ����h� ����h �H��h      D  , , �,��h �,��h� ����h� ����h �,��h      D  , , ���h ���h� ����h� ����h ���h      D  , , ����e� ����f ����f ����e� ����e�      D  , , ����e� ����f �j��f �j��e� ����e�      D  , , ����e� ����f �N��f �N��e� ����e�      D  , , ����e� ����f �2��f �2��e� ����e�      D  , , ����e� ����f ���f ���e� ����e�      D  , , ����c ����c� ����c� ����c ����c      D  , , ����c ����c� �j��c� �j��c ����c      D  , , ����c ����c� �N��c� �N��c ����c      D  , , ����c ����c� �2��c� �2��c ����c      D  , , ����c ����c� ���c� ���c ����c      D  , , �d��c �d��c� ����c� ����c �d��c      D  , , �H��c �H��c� ����c� ����c �H��c      D  , , �,��c �,��c� ����c� ����c �,��c      D  , , ���c ���c� ����c� ����c ���c      D  , , ����h ����h� ����h� ����h ����h      D  , , ����h ����h� �j��h� �j��h ����h      D  , , ����h ����h� �N��h� �N��h ����h      D  , , ����h ����h� �2��h� �2��h ����h      D  , , ����h ����h� ���h� ���h ����h      D  , , ����f� ����gX ����gX ����f� ����f�      D  , , ����f� ����gX �j��gX �j��f� ����f�      D  , , ����f� ����gX �N��gX �N��f� ����f�      D  , , ����f� ����gX �2��gX �2��f� ����f�      D  , , �d��e� �d��f ����f ����e� �d��e�      D  , , �H��e� �H��f ����f ����e� �H��e�      D  , , �,��e� �,��f ����f ����e� �,��e�      D  , , ���e� ���f ����f ����e� ���e�      D  , , ����[� ����\6 ����\6 ����[� ����[�      D  , , ����[� ����\6 �j��\6 �j��[� ����[�      D  , , ����[� ����\6 �N��\6 �N��[� ����[�      D  , , ����[� ����\6 �2��\6 �2��[� ����[�      D  , , ����[� ����\6 ���\6 ���[� ����[�      D  , , �d��[� �d��\6 ����\6 ����[� �d��[�      D  , , �H��[� �H��\6 ����\6 ����[� �H��[�      D  , , �,��[� �,��\6 ����\6 ����[� �,��[�      D  , , ���[� ���\6 ����\6 ����[� ���[�      D  , , ����f� ����gX ���gX ���f� ����f�      D  , , �d��f� �d��gX ����gX ����f� �d��f�      D  , , �H��f� �H��gX ����gX ����f� �H��f�      D  , , �,��f� �,��gX ����gX ����f� �,��f�      D  , , ���_� ���`� ����`� ����_� ���_�      D  , , ����_� ����`� ����`� ����_� ����_�      D  , , ����_� ����`� �l��`� �l��_� ����_�      D  , , ����_� ����`� �P��`� �P��_� ����_�      D  , , ����dB ����d� ����d� ����dB ����dB      D  , , ����dB ����d� �j��d� �j��dB ����dB      D  , , ����dB ����d� �N��d� �N��dB ����dB      D  , , ����dB ����d� �2��d� �2��dB ����dB      D  , , ����dB ����d� ���d� ���dB ����dB      D  , , �d��dB �d��d� ����d� ����dB �d��dB      D  , , �H��dB �H��d� ����d� ����dB �H��dB      D  , , �,��dB �,��d� ����d� ����dB �,��dB      D  , , ���dB ���d� ����d� ����dB ���dB      D  , , �b��^� �b��_G ����_G ����^� �b��^�      D  , , �F��^� �F��_G ����_G ����^� �F��^�      D  , , �*��^� �*��_G ����_G ����^� �*��^�      D  , , ���^� ���_G ����_G ����^� ���^�      D  , , ����^� ����_G ����_G ����^� ����^�      D  , , ����^� ����_G �l��_G �l��^� ����^�      D  , , ����^� ����_G �P��_G �P��^� ����^�      D  , , ����^� ����_G �4��_G �4��^� ����^�      D  , , ����_� ����`� �4��`� �4��_� ����_�      D  , , �|��c �|��c� ���c� ���c �|��c      D  , , �`��c �`��c� ����c� ����c �`��c      D  , , �D��c �D��c� ����c� ����c �D��c      D  , , �(��c �(��c� ����c� ����c �(��c      D  , , y���[� y���\6 zf��\6 zf��[� y���[�      D  , , |���[� |���\6 }J��\6 }J��[� |���[�      D  , , ���[� ���\6 �.��\6 �.��[� ���[�      D  , , �|��[� �|��\6 ���\6 ���[� �|��[�      D  , , �`��[� �`��\6 ����\6 ����[� �`��[�      D  , , �D��[� �D��\6 ����\6 ����[� �D��[�      D  , , �(��[� �(��\6 ����\6 ����[� �(��[�      D  , , ���[� ���\6 ����\6 ����[� ���[�      D  , , ���c ���c� ����c� ����c ���c      D  , , �~��_� �~��`� ���`� ���_� �~��_�      D  , , ~&��_� ~&��`� ~���`� ~���_� ~&��_�      D  , , y���e� y���f zf��f zf��e� y���e�      D  , , |���e� |���f }J��f }J��e� |���e�      D  , , ���e� ���f �.��f �.��e� ���e�      D  , , �|��e� �|��f ���f ���e� �|��e�      D  , , �`��e� �`��f ����f ����e� �`��e�      D  , , �D��e� �D��f ����f ����e� �D��e�      D  , , �(��e� �(��f ����f ����e� �(��e�      D  , , y���h y���h� zf��h� zf��h y���h      D  , , |���h |���h� }J��h� }J��h |���h      D  , , ���h ���h� ����h� ����h ���h      D  , , y���dB y���d� zf��d� zf��dB y���dB      D  , , |���dB |���d� }J��d� }J��dB |���dB      D  , , ���dB ���d� �.��d� �.��dB ���dB      D  , , �|��dB �|��d� ���d� ���dB �|��dB      D  , , �`��dB �`��d� ����d� ����dB �`��dB      D  , , �D��dB �D��d� ����d� ����dB �D��dB      D  , , �(��dB �(��d� ����d� ����dB �(��dB      D  , , x^��_� x^��`� x���`� x���_� x^��_�      D  , , {B��_� {B��`� {���`� {���_� {B��_�      D  , , ���e� ���f ����f ����e� ���e�      D  , , �
��_� �
��`� ����`� ����_� �
��_�      D  , , ����_� ����`� ����`� ����_� ����_�      D  , , ����_� ����`� �h��`� �h��_� ����_�      D  , , ���dB ���d� ����d� ����dB ���dB      D  , , ����_� ����`� �L��`� �L��_� ����_�      D  , , y���f� y���gX zf��gX zf��f� y���f�      D  , , |���f� |���gX }J��gX }J��f� |���f�      D  , , ���f� ���gX �.��gX �.��f� ���f�      D  , , ���h ���h� �.��h� �.��h ���h      D  , , �|��h �|��h� ���h� ���h �|��h      D  , , �`��h �`��h� ����h� ����h �`��h      D  , , �D��h �D��h� ����h� ����h �D��h      D  , , �(��h �(��h� ����h� ����h �(��h      D  , , x^��^� x^��_G x���_G x���^� x^��^�      D  , , {B��^� {B��_G {���_G {���^� {B��^�      D  , , ~&��^� ~&��_G ~���_G ~���^� ~&��^�      D  , , �
��^� �
��_G ����_G ����^� �
��^�      D  , , ����^� ����_G ����_G ����^� ����^�      D  , , ����^� ����_G �h��_G �h��^� ����^�      D  , , ����^� ����_G �L��_G �L��^� ����^�      D  , , ����^� ����_G �0��_G �0��^� ����^�      D  , , �~��^� �~��_G ���_G ���^� �~��^�      D  , , �|��f� �|��gX ���gX ���f� �|��f�      D  , , �`��f� �`��gX ����gX ����f� �`��f�      D  , , �D��f� �D��gX ����gX ����f� �D��f�      D  , , �(��f� �(��gX ����gX ����f� �(��f�      D  , , ���f� ���gX ����gX ����f� ���f�      D  , , ����_� ����`� �0��`� �0��_� ����_�      D  , , y���c y���c� zf��c� zf��c y���c      D  , , |���c |���c� }J��c� }J��c |���c      D  , , ���c ���c� �.��c� �.��c ���c      D  , , �D��P` �D��P� ����P� ����P` �D��P`      D  , , �(��P` �(��P� ����P� ����P` �(��P`      D  , , ���P` ���P� ����P� ����P` ���P`      D  , , ���R� ���Sv ����Sv ����R� ���R�      D  , , y���Y  y���Y� zf��Y� zf��Y  y���Y       D  , , |���Y  |���Y� }J��Y� }J��Y  |���Y       D  , , ���Y  ���Y� �.��Y� �.��Y  ���Y       D  , , �|��Y  �|��Y� ���Y� ���Y  �|��Y       D  , , �`��Y  �`��Y� ����Y� ����Y  �`��Y       D  , , �D��Y  �D��Y� ����Y� ����Y  �D��Y       D  , , �(��Y  �(��Y� ����Y� ����Y  �(��Y       D  , , ���Y  ���Y� ����Y� ����Y  ���Y       D  , , y���W� y���Xv zf��Xv zf��W� y���W�      D  , , y���V� y���W6 zf��W6 zf��V� y���V�      D  , , |���V� |���W6 }J��W6 }J��V� |���V�      D  , , ���V� ���W6 �.��W6 �.��V� ���V�      D  , , �|��V� �|��W6 ���W6 ���V� �|��V�      D  , , �`��V� �`��W6 ����W6 ����V� �`��V�      D  , , �D��V� �D��W6 ����W6 ����V� �D��V�      D  , , �(��V� �(��W6 ����W6 ����V� �(��V�      D  , , ���V� ���W6 ����W6 ����V� ���V�      D  , , y���O  y���O� zf��O� zf��O  y���O       D  , , |���O  |���O� }J��O� }J��O  |���O       D  , , ���O  ���O� �.��O� �.��O  ���O       D  , , �|��O  �|��O� ���O� ���O  �|��O       D  , , �`��O  �`��O� ����O� ����O  �`��O       D  , , �D��O  �D��O� ����O� ����O  �D��O       D  , , �(��O  �(��O� ����O� ����O  �(��O       D  , , ���O  ���O� ����O� ����O  ���O       D  , , |���W� |���Xv }J��Xv }J��W� |���W�      D  , , ���W� ���Xv �.��Xv �.��W� ���W�      D  , , �|��W� �|��Xv ���Xv ���W� �|��W�      D  , , �`��W� �`��Xv ����Xv ����W� �`��W�      D  , , �D��W� �D��Xv ����Xv ����W� �D��W�      D  , , �(��W� �(��Xv ����Xv ����W� �(��W�      D  , , ���W� ���Xv ����Xv ����W� ���W�      D  , , |���T  |���T� }J��T� }J��T  |���T       D  , , ���T  ���T� �.��T� �.��T  ���T       D  , , �|��T  �|��T� ���T� ���T  �|��T       D  , , �`��T  �`��T� ����T� ����T  �`��T       D  , , �D��T  �D��T� ����T� ����T  �D��T       D  , , �(��T  �(��T� ����T� ����T  �(��T       D  , , ���T  ���T� ����T� ����T  ���T       D  , , y���T  y���T� zf��T� zf��T  y���T       D  , , y���R� y���Sv zf��Sv zf��R� y���R�      D  , , |���R� |���Sv }J��Sv }J��R� |���R�      D  , , y���Q� y���R6 zf��R6 zf��Q� y���Q�      D  , , |���Q� |���R6 }J��R6 }J��Q� |���Q�      D  , , ���Q� ���R6 �.��R6 �.��Q� ���Q�      D  , , �|��Q� �|��R6 ���R6 ���Q� �|��Q�      D  , , �`��Q� �`��R6 ����R6 ����Q� �`��Q�      D  , , �D��Q� �D��R6 ����R6 ����Q� �D��Q�      D  , , �(��Q� �(��R6 ����R6 ����Q� �(��Q�      D  , , ���Q� ���R6 ����R6 ����Q� ���Q�      D  , , ���R� ���Sv �.��Sv �.��R� ���R�      D  , , �|��R� �|��Sv ���Sv ���R� �|��R�      D  , , �`��R� �`��Sv ����Sv ����R� �`��R�      D  , , �D��R� �D��Sv ����Sv ����R� �D��R�      D  , , �(��R� �(��Sv ����Sv ����R� �(��R�      D  , , y���P` y���P� zf��P� zf��P` y���P`      D  , , y���M� y���Nv zf��Nv zf��M� y���M�      D  , , |���M� |���Nv }J��Nv }J��M� |���M�      D  , , ���M� ���Nv �.��Nv �.��M� ���M�      D  , , �|��M� �|��Nv ���Nv ���M� �|��M�      D  , , �`��M� �`��Nv ����Nv ����M� �`��M�      D  , , �D��M� �D��Nv ����Nv ����M� �D��M�      D  , , �(��M� �(��Nv ����Nv ����M� �(��M�      D  , , ���M� ���Nv ����Nv ����M� ���M�      D  , , |���P` |���P� }J��P� }J��P` |���P`      D  , , ���P` ���P� �.��P� �.��P` ���P`      D  , , �|��P` �|��P� ���P� ���P` �|��P`      D  , , y���U` y���U� zf��U� zf��U` y���U`      D  , , |���U` |���U� }J��U� }J��U` |���U`      D  , , ���U` ���U� �.��U� �.��U` ���U`      D  , , �|��U` �|��U� ���U� ���U` �|��U`      D  , , �`��U` �`��U� ����U� ����U` �`��U`      D  , , �D��U` �D��U� ����U� ����U` �D��U`      D  , , �(��U` �(��U� ����U� ����U` �(��U`      D  , , ���U` ���U� ����U� ����U` ���U`      D  , , �`��P` �`��P� ����P� ����P` �`��P`      D  , , y���Z` y���Z� zf��Z� zf��Z` y���Z`      D  , , |���Z` |���Z� }J��Z� }J��Z` |���Z`      D  , , ���Z` ���Z� �.��Z� �.��Z` ���Z`      D  , , �|��Z` �|��Z� ���Z� ���Z` �|��Z`      D  , , �`��Z` �`��Z� ����Z� ����Z` �`��Z`      D  , , �D��Z` �D��Z� ����Z� ����Z` �D��Z`      D  , , �(��Z` �(��Z� ����Z� ����Z` �(��Z`      D  , , ���Z` ���Z� ����Z� ����Z` ���Z`      D  , , y���L� y���M6 zf��M6 zf��L� y���L�      D  , , |���L� |���M6 }J��M6 }J��L� |���L�      D  , , ���L� ���M6 �.��M6 �.��L� ���L�      D  , , �|��L� �|��M6 ���M6 ���L� �|��L�      D  , , �`��L� �`��M6 ����M6 ����L� �`��L�      D  , , �D��L� �D��M6 ����M6 ����L� �D��L�      D  , , �(��L� �(��M6 ����M6 ����L� �(��L�      D  , , ���L� ���M6 ����M6 ����L� ���L�      D  , , ����V� ����W6 ���W6 ���V� ����V�      D  , , ����Q� ����R6 ���R6 ���Q� ����Q�      D  , , ����Y  ����Y� ���Y� ���Y  ����Y       D  , , ����P` ����P� ���P� ���P` ����P`      D  , , ����T  ����T� ���T� ���T  ����T       D  , , ����M� ����Nv ���Nv ���M� ����M�      D  , , ����W� ����Xv ���Xv ���W� ����W�      D  , , ����R� ����Sv ���Sv ���R� ����R�      D  , , ����U` ����U� ���U� ���U` ����U`      D  , , ����O  ����O� ���O� ���O  ����O       D  , , ����Z` ����Z� ���Z� ���Z` ����Z`      D  , , ����L� ����M6 ���M6 ���L� ����L�      D  , , �H��Y  �H��Y� ����Y� ����Y  �H��Y       D  , , ���V� ���W6 ����W6 ����V� ���V�      D  , , �d��T  �d��T� ����T� ����T  �d��T       D  , , �H��T  �H��T� ����T� ����T  �H��T       D  , , �,��T  �,��T� ����T� ����T  �,��T       D  , , �,��W� �,��Xv ����Xv ����W� �,��W�      D  , , ���W� ���Xv ����Xv ����W� ���W�      D  , , �d��W� �d��Xv ����Xv ����W� �d��W�      D  , , �H��W� �H��Xv ����Xv ����W� �H��W�      D  , , �,��Y  �,��Y� ����Y� ����Y  �,��Y       D  , , ���Y  ���Y� ����Y� ����Y  ���Y       D  , , �d��V� �d��W6 ����W6 ����V� �d��V�      D  , , �H��V� �H��W6 ����W6 ����V� �H��V�      D  , , �d��U` �d��U� ����U� ����U` �d��U`      D  , , �H��U` �H��U� ����U� ����U` �H��U`      D  , , �,��U` �,��U� ����U� ����U` �,��U`      D  , , ���U` ���U� ����U� ����U` ���U`      D  , , ���T  ���T� ����T� ����T  ���T       D  , , �d��Y  �d��Y� ����Y� ����Y  �d��Y       D  , , �d��Z` �d��Z� ����Z� ����Z` �d��Z`      D  , , �H��Z` �H��Z� ����Z� ����Z` �H��Z`      D  , , �,��Z` �,��Z� ����Z� ����Z` �,��Z`      D  , , ���Z` ���Z� ����Z� ����Z` ���Z`      D  , , �,��V� �,��W6 ����W6 ����V� �,��V�      D  , , ����U` ����U� ����U� ����U` ����U`      D  , , ����U` ����U� �j��U� �j��U` ����U`      D  , , ����U` ����U� �N��U� �N��U` ����U`      D  , , ����U` ����U� �2��U� �2��U` ����U`      D  , , ����Y  ����Y� �2��Y� �2��Y  ����Y       D  , , ����W� ����Xv ����Xv ����W� ����W�      D  , , ����W� ����Xv �j��Xv �j��W� ����W�      D  , , ����W� ����Xv �N��Xv �N��W� ����W�      D  , , ����Y  ����Y� ����Y� ����Y  ����Y       D  , , ����W� ����Xv �2��Xv �2��W� ����W�      D  , , ����Z` ����Z� ����Z� ����Z` ����Z`      D  , , ����Z` ����Z� �j��Z� �j��Z` ����Z`      D  , , ����Z` ����Z� �N��Z� �N��Z` ����Z`      D  , , ����Z` ����Z� �2��Z� �2��Z` ����Z`      D  , , ����T  ����T� �j��T� �j��T  ����T       D  , , ����T  ����T� �N��T� �N��T  ����T       D  , , ����T  ����T� �2��T� �2��T  ����T       D  , , ����Y  ����Y� �j��Y� �j��Y  ����Y       D  , , ����T  ����T� ����T� ����T  ����T       D  , , ����V� ����W6 ����W6 ����V� ����V�      D  , , ����V� ����W6 �j��W6 �j��V� ����V�      D  , , ����V� ����W6 �N��W6 �N��V� ����V�      D  , , ����V� ����W6 �2��W6 �2��V� ����V�      D  , , ����Y  ����Y� �N��Y� �N��Y  ����Y       D  , , ����Q� ����R6 �j��R6 �j��Q� ����Q�      D  , , ����O  ����O� ����O� ����O  ����O       D  , , ����O  ����O� �j��O� �j��O  ����O       D  , , ����O  ����O� �N��O� �N��O  ����O       D  , , ����O  ����O� �2��O� �2��O  ����O       D  , , ����R� ����Sv ����Sv ����R� ����R�      D  , , ����R� ����Sv �j��Sv �j��R� ����R�      D  , , ����Q� ����R6 �N��R6 �N��Q� ����Q�      D  , , ����Q� ����R6 �2��R6 �2��Q� ����Q�      D  , , ����R� ����Sv �N��Sv �N��R� ����R�      D  , , ����R� ����Sv �2��Sv �2��R� ����R�      D  , , ����Q� ����R6 ����R6 ����Q� ����Q�      D  , , ����M� ����Nv ����Nv ����M� ����M�      D  , , ����M� ����Nv �j��Nv �j��M� ����M�      D  , , ����M� ����Nv �N��Nv �N��M� ����M�      D  , , ����M� ����Nv �2��Nv �2��M� ����M�      D  , , ����P` ����P� ����P� ����P` ����P`      D  , , ����P` ����P� �j��P� �j��P` ����P`      D  , , ����P` ����P� �N��P� �N��P` ����P`      D  , , ����L� ����M6 ����M6 ����L� ����L�      D  , , ����L� ����M6 �j��M6 �j��L� ����L�      D  , , ����L� ����M6 �N��M6 �N��L� ����L�      D  , , ����L� ����M6 �2��M6 �2��L� ����L�      D  , , ����P` ����P� �2��P� �2��P` ����P`      D  , , �d��Q� �d��R6 ����R6 ����Q� �d��Q�      D  , , �d��P` �d��P� ����P� ����P` �d��P`      D  , , �H��P` �H��P� ����P� ����P` �H��P`      D  , , �,��P` �,��P� ����P� ����P` �,��P`      D  , , ���P` ���P� ����P� ����P` ���P`      D  , , �d��R� �d��Sv ����Sv ����R� �d��R�      D  , , �H��R� �H��Sv ����Sv ����R� �H��R�      D  , , �d��O  �d��O� ����O� ����O  �d��O       D  , , �H��O  �H��O� ����O� ����O  �H��O       D  , , �,��O  �,��O� ����O� ����O  �,��O       D  , , ���O  ���O� ����O� ����O  ���O       D  , , �,��R� �,��Sv ����Sv ����R� �,��R�      D  , , ���R� ���Sv ����Sv ����R� ���R�      D  , , �d��M� �d��Nv ����Nv ����M� �d��M�      D  , , �H��M� �H��Nv ����Nv ����M� �H��M�      D  , , �,��M� �,��Nv ����Nv ����M� �,��M�      D  , , ���M� ���Nv ����Nv ����M� ���M�      D  , , �H��Q� �H��R6 ����R6 ����Q� �H��Q�      D  , , �,��Q� �,��R6 ����R6 ����Q� �,��Q�      D  , , ���Q� ���R6 ����R6 ����Q� ���Q�      D  , , �d��L� �d��M6 ����M6 ����L� �d��L�      D  , , �H��L� �H��M6 ����M6 ����L� �H��L�      D  , , �,��L� �,��M6 ����M6 ����L� �,��L�      D  , , ���L� ���M6 ����M6 ����L� ���L�      D  , , ���f� ���gX ª��gX ª��f� ���f�      D  , , ���W� ���Xv ª��Xv ª��W� ���W�      D  , , ���V� ���W6 ª��W6 ª��V� ���V�      D  , , ���T  ���T� ª��T� ª��T  ���T       D  , , ���P` ���P� ª��P� ª��P` ���P`      D  , , ���[� ���\6 ª��\6 ª��[� ���[�      D  , , ���e� ���f ª��f ª��e� ���e�      D  , , ���Z` ���Z� ª��Z� ª��Z` ���Z`      D  , , ���O  ���O� ª��O� ª��O  ���O       D  , , ���Y  ���Y� ª��Y� ª��Y  ���Y       D  , , ���R� ���Sv ª��Sv ª��R� ���R�      D  , , ���U` ���U� ª��U� ª��U` ���U`      D  , , ���M� ���Nv ª��Nv ª��M� ���M�      D  , , ���c ���c� ª��c� ª��c ���c      D  , , ���dB ���d� ª��d� ª��dB ���dB      D  , , ���h ���h� ª��h� ª��h ���h      D  , , ���Q� ���R6 ª��R6 ª��Q� ���Q�      D  , , ���L� ���M6 ª��M6 ª��L� ���L�      D  , , ����[� ����\6 Ŏ��\6 Ŏ��[� ����[�      D  , , ����[� ����\6 �r��\6 �r��[� ����[�      D  , , ����[� ����\6 �V��\6 �V��[� ����[�      D  , , ͤ��[� ͤ��\6 �:��\6 �:��[� ͤ��[�      D  , , ���[� ���\@ Ӟ��\@ Ӟ��[� ���[�      D  , , �m��[� �m��\@ ���\@ ���[� �m��[�      D  , , ����[i ����[� �}��[� �}��[i ����[i      D  , , �j��_� �j��`� � ��`� � ��_� �j��_�      D  , , ���_j ���`  Ӟ��`  Ӟ��_j ���_j      D  , , �m��_j �m��`  ���`  ���_j �m��_j      D  , , ���\� ���]� Ӟ��]� Ӟ��\� ���\�      D  , , �m��\� �m��]� ���]� ���\� �m��\�      D  , , ����\� ����]? �}��]? �}��\� ����\�      D  , , �N��_� �N��`� ����`� ����_� �N��_�      D  , , ����f� ����gX �V��gX �V��f� ����f�      D  , , ����e� ����f Ŏ��f Ŏ��e� ����e�      D  , , ����e� ����f �r��f �r��e� ����e�      D  , , ����e� ����f �V��f �V��e� ����e�      D  , , ���a� ���b� Ӟ��b� Ӟ��a� ���a�      D  , , �2��_� �2��`� ����`� ����_� �2��_�      D  , , ����`i ����`� �}��`� �}��`i ����`i      D  , , ͤ��f� ͤ��gX �:��gX �:��f� ͤ��f�      D  , , �m��^* �m��^� ���^� ���^* �m��^*      D  , , �m��a� �m��b� ���b� ���a� �m��a�      D  , , ����a� ����b? �}��b? �}��a� ����a�      D  , , ͤ��e� ͤ��f �:��f �:��e� ͤ��e�      D  , , ���e� ���f@ Ӟ��f@ Ӟ��e� ���e�      D  , , �m��e� �m��f@ ���f@ ���e� �m��e�      D  , , ����ei ����e� �}��e� �}��ei ����ei      D  , , ����]� ����^ �}��^ �}��]� ����]�      D  , , ���^* ���^� Ӟ��^� Ӟ��^* ���^*      D  , , ���f� ���g� Ӟ��g� Ӟ��f� ���f�      D  , , Æ��^� Æ��_G ���_G ���^� Æ��^�      D  , , �j��^� �j��_G � ��_G � ��^� �j��^�      D  , , �N��^� �N��_G ����_G ����^� �N��^�      D  , , �2��^� �2��_G ����_G ����^� �2��^�      D  , , ����_) ����_� �}��_� �}��_) ����_)      D  , , �m��f� �m��g� ���g� ���f� �m��f�      D  , , ���`� ���a@ Ӟ��a@ Ӟ��`� ���`�      D  , , �m��`� �m��a@ ���a@ ���`� �m��`�      D  , , ����f� ����g? �}��g? �}��f� ����f�      D  , , ����c ����c� Ŏ��c� Ŏ��c ����c      D  , , ����c ����c� �r��c� �r��c ����c      D  , , ����c ����c� �V��c� �V��c ����c      D  , , ͤ��c ͤ��c� �:��c� �:��c ͤ��c      D  , , ���c* ���c� Ӟ��c� Ӟ��c* ���c*      D  , , �m��c* �m��c� ���c� ���c* �m��c*      D  , , ����b� ����c �}��c �}��b� ����b�      D  , , ����g� ����h �}��h �}��g� ����g�      D  , , ����dB ����d� Ŏ��d� Ŏ��dB ����dB      D  , , ����dB ����d� �r��d� �r��dB ����dB      D  , , ����dB ����d� �V��d� �V��dB ����dB      D  , , ͤ��dB ͤ��d� �:��d� �:��dB ͤ��dB      D  , , ���dj ���e  Ӟ��e  Ӟ��dj ���dj      D  , , �m��dj �m��e  ���e  ���dj �m��dj      D  , , ����d) ����d� �}��d� �}��d) ����d)      D  , , ����f� ����gX Ŏ��gX Ŏ��f� ����f�      D  , , ����h ����h� Ŏ��h� Ŏ��h ����h      D  , , ����h ����h� �r��h� �r��h ����h      D  , , ����h ����h� �V��h� �V��h ����h      D  , , ͤ��h ͤ��h� �:��h� �:��h ͤ��h      D  , , ���h* ���h� Ӟ��h� Ӟ��h* ���h*      D  , , �m��h* �m��h� ���h� ���h* �m��h*      D  , , Æ��_� Æ��`� ���`� ���_� Æ��_�      D  , , ����f� ����gX �r��gX �r��f� ����f�      D  , , ����^� ����_G �T��_G �T��^� ����^�      D  , , �0��[� �0��\6 ����\6 ����[� �0��[�      D  , , �h��f� �h��gX ����gX ����f� �h��f�      D  , , �L��f� �L��gX ����gX ����f� �L��f�      D  , , ����_� ����`� ���`� ���_� ����_�      D  , , �f��_� �f��`� ����`� ����_� �f��_�      D  , , �J��_� �J��`� ����`� ����_� �J��_�      D  , , �0��f� �0��gX ����gX ����f� �0��f�      D  , , �.��_� �.��`� ����`� ����_� �.��_�      D  , , ����h ����h� ���h� ���h ����h      D  , , �h��h �h��h� ����h� ����h �h��h      D  , , �L��h �L��h� ����h� ����h �L��h      D  , , �0��h �0��h� ����h� ����h �0��h      D  , , ���_� ���`� ����`� ����_� ���_�      D  , , ����^� ����_G �8��_G �8��^� ����^�      D  , , ����_� ����`� ����`� ����_� ����_�      D  , , ����_� ����`� �p��`� �p��_� ����_�      D  , , ����_� ����`� �T��`� �T��_� ����_�      D  , , ����_� ����`� �8��`� �8��_� ����_�      D  , , ����e� ����f ����f ����e� ����e�      D  , , ����dB ����d� ���d� ���dB ����dB      D  , , ����c ����c� ����c� ����c ����c      D  , , ����c ����c� �n��c� �n��c ����c      D  , , ����dB ����d� ����d� ����dB ����dB      D  , , ����dB ����d� �n��d� �n��dB ����dB      D  , , ����e� ����f �n��f �n��e� ����e�      D  , , ����c ����c� �R��c� �R��c ����c      D  , , ����c ����c� �6��c� �6��c ����c      D  , , ����c ����c� ���c� ���c ����c      D  , , �h��c �h��c� ����c� ����c �h��c      D  , , �L��c �L��c� ����c� ����c �L��c      D  , , �0��c �0��c� ����c� ����c �0��c      D  , , ����e� ����f �R��f �R��e� ����e�      D  , , ����e� ����f �6��f �6��e� ����e�      D  , , ����e� ����f ���f ���e� ����e�      D  , , �h��e� �h��f ����f ����e� �h��e�      D  , , �L��e� �L��f ����f ����e� �L��e�      D  , , �0��e� �0��f ����f ����e� �0��e�      D  , , ����dB ����d� �R��d� �R��dB ����dB      D  , , ����dB ����d� �6��d� �6��dB ����dB      D  , , �h��dB �h��d� ����d� ����dB �h��dB      D  , , �L��dB �L��d� ����d� ����dB �L��dB      D  , , �0��dB �0��d� ����d� ����dB �0��dB      D  , , ����[� ����\6 ����\6 ����[� ����[�      D  , , ����[� ����\6 �n��\6 �n��[� ����[�      D  , , ����[� ����\6 �R��\6 �R��[� ����[�      D  , , ����[� ����\6 �6��\6 �6��[� ����[�      D  , , ����h ����h� �n��h� �n��h ����h      D  , , ����[� ����\6 ���\6 ���[� ����[�      D  , , �h��[� �h��\6 ����\6 ����[� �h��[�      D  , , ����h ����h� ����h� ����h ����h      D  , , ����h ����h� �R��h� �R��h ����h      D  , , ����h ����h� �6��h� �6��h ����h      D  , , ����^� ����_G ���_G ���^� ����^�      D  , , �f��^� �f��_G ����_G ����^� �f��^�      D  , , �J��^� �J��_G ����_G ����^� �J��^�      D  , , �L��[� �L��\6 ����\6 ����[� �L��[�      D  , , �.��^� �.��_G ����_G ����^� �.��^�      D  , , ���^� ���_G ����_G ����^� ���^�      D  , , ����^� ����_G ����_G ����^� ����^�      D  , , ����f� ����gX ����gX ����f� ����f�      D  , , ����f� ����gX �n��gX �n��f� ����f�      D  , , ����f� ����gX �R��gX �R��f� ����f�      D  , , ����f� ����gX �6��gX �6��f� ����f�      D  , , ����f� ����gX ���gX ���f� ����f�      D  , , ����^� ����_G �p��_G �p��^� ����^�      D  , , ����V� ����W6 ���W6 ���V� ����V�      D  , , ����U` ����U� ����U� ����U` ����U`      D  , , ����U` ����U� �n��U� �n��U` ����U`      D  , , ����U` ����U� �R��U� �R��U` ����U`      D  , , ����U` ����U� �6��U� �6��U` ����U`      D  , , ����U` ����U� ���U� ���U` ����U`      D  , , �h��U` �h��U� ����U� ����U` �h��U`      D  , , �L��U` �L��U� ����U� ����U` �L��U`      D  , , �0��U` �0��U� ����U� ����U` �0��U`      D  , , �L��W� �L��Xv ����Xv ����W� �L��W�      D  , , �h��V� �h��W6 ����W6 ����V� �h��V�      D  , , ����P` ����P� ����P� ����P` ����P`      D  , , �L��Z` �L��Z� ����Z� ����Z` �L��Z`      D  , , �0��Z` �0��Z� ����Z� ����Z` �0��Z`      D  , , ����P` ����P� �n��P� �n��P` ����P`      D  , , ����P` ����P� �R��P� �R��P` ����P`      D  , , ����P` ����P� �6��P� �6��P` ����P`      D  , , ����P` ����P� ���P� ���P` ����P`      D  , , �h��P` �h��P� ����P� ����P` �h��P`      D  , , ����M� ����Nv ����Nv ����M� ����M�      D  , , ����M� ����Nv �n��Nv �n��M� ����M�      D  , , ����M� ����Nv �R��Nv �R��M� ����M�      D  , , ����M� ����Nv �6��Nv �6��M� ����M�      D  , , ����M� ����Nv ���Nv ���M� ����M�      D  , , �h��M� �h��Nv ����Nv ����M� �h��M�      D  , , �L��M� �L��Nv ����Nv ����M� �L��M�      D  , , �0��M� �0��Nv ����Nv ����M� �0��M�      D  , , �L��P` �L��P� ����P� ����P` �L��P`      D  , , �0��P` �0��P� ����P� ����P` �0��P`      D  , , ����O  ����O� ����O� ����O  ����O       D  , , ����O  ����O� �n��O� �n��O  ����O       D  , , ����O  ����O� �R��O� �R��O  ����O       D  , , ����O  ����O� �6��O� �6��O  ����O       D  , , ����O  ����O� ���O� ���O  ����O       D  , , �h��O  �h��O� ����O� ����O  �h��O       D  , , �L��O  �L��O� ����O� ����O  �L��O       D  , , �0��O  �0��O� ����O� ����O  �0��O       D  , , �L��V� �L��W6 ����W6 ����V� �L��V�      D  , , �0��V� �0��W6 ����W6 ����V� �0��V�      D  , , �0��W� �0��Xv ����Xv ����W� �0��W�      D  , , ����T  ����T� ����T� ����T  ����T       D  , , ����T  ����T� �n��T� �n��T  ����T       D  , , ����T  ����T� �R��T� �R��T  ����T       D  , , ����Y  ����Y� ����Y� ����Y  ����Y       D  , , ����Y  ����Y� �n��Y� �n��Y  ����Y       D  , , ����Y  ����Y� �R��Y� �R��Y  ����Y       D  , , ����Y  ����Y� �6��Y� �6��Y  ����Y       D  , , ����Y  ����Y� ���Y� ���Y  ����Y       D  , , �h��Y  �h��Y� ����Y� ����Y  �h��Y       D  , , ����T  ����T� �6��T� �6��T  ����T       D  , , ����T  ����T� ���T� ���T  ����T       D  , , �h��T  �h��T� ����T� ����T  �h��T       D  , , �L��T  �L��T� ����T� ����T  �L��T       D  , , �0��T  �0��T� ����T� ����T  �0��T       D  , , �h��W� �h��Xv ����Xv ����W� �h��W�      D  , , �L��Y  �L��Y� ����Y� ����Y  �L��Y       D  , , �0��Y  �0��Y� ����Y� ����Y  �0��Y       D  , , ����V� ����W6 ����W6 ����V� ����V�      D  , , ����R� ����Sv ����Sv ����R� ����R�      D  , , ����R� ����Sv �n��Sv �n��R� ����R�      D  , , ����R� ����Sv �R��Sv �R��R� ����R�      D  , , ����R� ����Sv �6��Sv �6��R� ����R�      D  , , ����R� ����Sv ���Sv ���R� ����R�      D  , , ����W� ����Xv ����Xv ����W� ����W�      D  , , ����W� ����Xv �n��Xv �n��W� ����W�      D  , , ����Q� ����R6 ����R6 ����Q� ����Q�      D  , , ����Q� ����R6 �n��R6 �n��Q� ����Q�      D  , , ����Q� ����R6 �R��R6 �R��Q� ����Q�      D  , , ����Q� ����R6 �6��R6 �6��Q� ����Q�      D  , , ����Z` ����Z� ����Z� ����Z` ����Z`      D  , , ����Z` ����Z� �n��Z� �n��Z` ����Z`      D  , , ����Z` ����Z� �R��Z� �R��Z` ����Z`      D  , , ����Z` ����Z� �6��Z� �6��Z` ����Z`      D  , , ����Z` ����Z� ���Z� ���Z` ����Z`      D  , , ����Q� ����R6 ���R6 ���Q� ����Q�      D  , , �h��Q� �h��R6 ����R6 ����Q� �h��Q�      D  , , �L��Q� �L��R6 ����R6 ����Q� �L��Q�      D  , , �0��Q� �0��R6 ����R6 ����Q� �0��Q�      D  , , �h��R� �h��Sv ����Sv ����R� �h��R�      D  , , ����W� ����Xv �R��Xv �R��W� ����W�      D  , , ����W� ����Xv �6��Xv �6��W� ����W�      D  , , ����W� ����Xv ���Xv ���W� ����W�      D  , , �L��R� �L��Sv ����Sv ����R� �L��R�      D  , , �0��R� �0��Sv ����Sv ����R� �0��R�      D  , , ����V� ����W6 �n��W6 �n��V� ����V�      D  , , ����V� ����W6 �R��W6 �R��V� ����V�      D  , , �h��Z` �h��Z� ����Z� ����Z` �h��Z`      D  , , ����L� ����M6 ����M6 ����L� ����L�      D  , , ����L� ����M6 �n��M6 �n��L� ����L�      D  , , ����L� ����M6 �R��M6 �R��L� ����L�      D  , , ����L� ����M6 �6��M6 �6��L� ����L�      D  , , ����L� ����M6 ���M6 ���L� ����L�      D  , , �h��L� �h��M6 ����M6 ����L� �h��L�      D  , , �L��L� �L��M6 ����M6 ����L� �L��L�      D  , , �0��L� �0��M6 ����M6 ����L� �0��L�      D  , , ����V� ����W6 �6��W6 �6��V� ����V�      D  , , ����Z) ����Z� �}��Z� �}��Z) ����Z)      D  , , ����Y  ����Y� Ŏ��Y� Ŏ��Y  ����Y       D  , , ����V� ����W6 Ŏ��W6 Ŏ��V� ����V�      D  , , ����P` ����P� Ŏ��P� Ŏ��P` ����P`      D  , , ����P` ����P� �r��P� �r��P` ����P`      D  , , ����O  ����O� Ŏ��O� Ŏ��O  ����O       D  , , ����O  ����O� �r��O� �r��O  ����O       D  , , ����O  ����O� �V��O� �V��O  ����O       D  , , ͤ��O  ͤ��O� �:��O� �:��O  ͤ��O       D  , , ����P` ����P� �V��P� �V��P` ����P`      D  , , ͤ��P` ͤ��P� �:��P� �:��P` ͤ��P`      D  , , ����R� ����Sv Ŏ��Sv Ŏ��R� ����R�      D  , , ����R� ����Sv �r��Sv �r��R� ����R�      D  , , ����R� ����Sv �V��Sv �V��R� ����R�      D  , , ����M� ����Nv Ŏ��Nv Ŏ��M� ����M�      D  , , ����M� ����Nv �r��Nv �r��M� ����M�      D  , , ����M� ����Nv �V��Nv �V��M� ����M�      D  , , ͤ��M� ͤ��Nv �:��Nv �:��M� ͤ��M�      D  , , ͤ��R� ͤ��Sv �:��Sv �:��R� ͤ��R�      D  , , ����Y  ����Y� �r��Y� �r��Y  ����Y       D  , , ����Y  ����Y� �V��Y� �V��Y  ����Y       D  , , ͤ��Y  ͤ��Y� �:��Y� �:��Y  ͤ��Y       D  , , ����Z` ����Z� Ŏ��Z� Ŏ��Z` ����Z`      D  , , ����Z` ����Z� �r��Z� �r��Z` ����Z`      D  , , ����Z` ����Z� �V��Z� �V��Z` ����Z`      D  , , ͤ��Z` ͤ��Z� �:��Z� �:��Z` ͤ��Z`      D  , , ����Q� ����R6 Ŏ��R6 Ŏ��Q� ����Q�      D  , , ����Q� ����R6 �r��R6 �r��Q� ����Q�      D  , , ����Q� ����R6 �V��R6 �V��Q� ����Q�      D  , , ͤ��Q� ͤ��R6 �:��R6 �:��Q� ͤ��Q�      D  , , ����T  ����T� Ŏ��T� Ŏ��T  ����T       D  , , ���Zj ���[  Ӟ��[  Ӟ��Zj ���Zj      D  , , �m��Zj �m��[  ���[  ���Zj �m��Zj      D  , , ����T  ����T� �r��T� �r��T  ����T       D  , , ����T  ����T� �V��T� �V��T  ����T       D  , , ͤ��T  ͤ��T� �:��T� �:��T  ͤ��T       D  , , ����V� ����W6 �r��W6 �r��V� ����V�      D  , , ����V� ����W6 �V��W6 �V��V� ����V�      D  , , ͤ��V� ͤ��W6 �:��W6 �:��V� ͤ��V�      D  , , ����U` ����U� Ŏ��U� Ŏ��U` ����U`      D  , , ����U` ����U� �r��U� �r��U` ����U`      D  , , ����U` ����U� �V��U� �V��U` ����U`      D  , , ͤ��U` ͤ��U� �:��U� �:��U` ͤ��U`      D  , , ����W� ����Xv Ŏ��Xv Ŏ��W� ����W�      D  , , ����W� ����Xv �r��Xv �r��W� ����W�      D  , , ����W� ����Xv �V��Xv �V��W� ����W�      D  , , ͤ��W� ͤ��Xv �:��Xv �:��W� ͤ��W�      D  , , ����L� ����M6 Ŏ��M6 Ŏ��L� ����L�      D  , , ����L� ����M6 �r��M6 �r��L� ����L�      D  , , ����L� ����M6 �V��M6 �V��L� ����L�      D  , , ͤ��L� ͤ��M6 �:��M6 �:��L� ͤ��L�      E  , , ���qq ���r9 S��r9 S��qq ���qq      E  , , ���o� ���p� S��p� S��o� ���o�      E  , , ���nQ ���o S��o S��nQ ���nQ      E  , , ���l� ���m� S��m� S��l� ���l�      E  , , ���k1 ���k� S��k� S��k1 ���k1      E  , , ���i� ���ji S��ji S��i� ���i�      E  , , ���h ���h� S��h� S��h ���h      E  , , ���f� ���gI S��gI S��f� ���f�      E  , , ���d� ���e� S��e� S��d� ���d�      E  , , ���ca ���d) S��d) S��ca ���ca      E  , , ���[ ���[� S��[� S��[ ���[      E  , , ���Y ���ZG S��ZG S��Y ���Y      E  , , ���W� ���X� S��X� S��W� ���W�      E  , , ���V_ ���W' S��W' S��V_ ���V_      E  , , ���T� ���U� S��U� S��T� ���T�      E  , , ���S? ���T S��T S��S? ���S?      E  , , ���Q� ���Rw S��Rw S��Q� ���Q�      E  , , ���P ���P� S��P� S��P ���P      E  , , ���N� ���OW S��OW S��N� ���N�      E  , , ���L� ���M� S��M� S��L� ���L�      E  , , ��  2� ��  3� ��  3� ��  2� ��  2�      E  , , ��  1V ��  2 ��  2 ��  1V ��  1V      E  , , ��  /� ��  0� ��  0� ��  /� ��  /�      E  , , ��  .6 ��  .� ��  .� ��  .6 ��  .6      E  , , ��  ,� ��  -n ��  -n ��  ,� ��  ,�      E  , , ��  + ��  +� ��  +� ��  + ��  +      E  , , ��  )� ��  *N ��  *N ��  )� ��  )�      E  , , ��  "� ��  #Z ��  #Z ��  "� ��  "�      E  , , ��  ! ��  !� ��  !� ��  ! ��  !      E  , , ��  r ��   : ��   : ��  r ��  r      E  , , ��  � ��  � ��  � ��  � ��  �      E  , , ��  R ��   ��   ��  R ��  R      E  , , ��  � ��  � ��  � ��  � ��  �      E  , , ��  2 ��  � ��  � ��  2 ��  2      E  , , ŉ  1V ŉ  2 �Q  2 �Q  1V ŉ  1V      E  , , �%  1V �%  2 ��  2 ��  1V �%  1V      E  , , ��  1V ��  2 ω  2 ω  1V ��  1V      E  , , ŉ  /� ŉ  0� �Q  0� �Q  /� ŉ  /�      E  , , �%  /� �%  0� ��  0� ��  /� �%  /�      E  , , ��  /� ��  0� ω  0� ω  /� ��  /�      E  , , ŉ  .6 ŉ  .� �Q  .� �Q  .6 ŉ  .6      E  , , �%  .6 �%  .� ��  .� ��  .6 �%  .6      E  , , ��  .6 ��  .� ω  .� ω  .6 ��  .6      E  , , ŉ  ,� ŉ  -n �Q  -n �Q  ,� ŉ  ,�      E  , , �%  ,� �%  -n ��  -n ��  ,� �%  ,�      E  , , ��  ,� ��  -n ω  -n ω  ,� ��  ,�      E  , , ŉ  + ŉ  +� �Q  +� �Q  + ŉ  +      E  , , �%  + �%  +� ��  +� ��  + �%  +      E  , , ��  + ��  +� ω  +� ω  + ��  +      E  , , ŉ  2� ŉ  3� �Q  3� �Q  2� ŉ  2�      E  , , ŉ  )� ŉ  *N �Q  *N �Q  )� ŉ  )�      E  , , �%  )� �%  *N ��  *N ��  )� �%  )�      E  , , ��  )� ��  *N ω  *N ω  )� ��  )�      E  , , �%  2� �%  3� ��  3� ��  2� �%  2�      E  , , ��  2� ��  3� ω  3� ω  2� ��  2�      E  , , �Q  /� �Q  0� �  0� �  /� �Q  /�      E  , , �Q  2� �Q  3� �  3� �  2� �Q  2�      E  , , �}  ,� �}  -n �E  -n �E  ,� �}  ,�      E  , , �  ,� �  -n ��  -n ��  ,� �  ,�      E  , , ��  ,� ��  -n �}  -n �}  ,� ��  ,�      E  , , �Q  ,� �Q  -n �  -n �  ,� �Q  ,�      E  , , ��  ,� ��  -n ��  -n ��  ,� ��  ,�      E  , , ��  /� ��  0� ��  0� ��  /� ��  /�      E  , , ��  1V ��  2 ��  2 ��  1V ��  1V      E  , , �  2� �  3� ��  3� ��  2� �  2�      E  , , ��  2� ��  3� ��  3� ��  2� ��  2�      E  , , �}  + �}  +� �E  +� �E  + �}  +      E  , , �  + �  +� ��  +� ��  + �  +      E  , , ��  + ��  +� �}  +� �}  + ��  +      E  , , �Q  + �Q  +� �  +� �  + �Q  +      E  , , ��  + ��  +� ��  +� ��  + ��  +      E  , , �}  /� �}  0� �E  0� �E  /� �}  /�      E  , , ��  2� ��  3� �}  3� �}  2� ��  2�      E  , , �}  .6 �}  .� �E  .� �E  .6 �}  .6      E  , , �  .6 �  .� ��  .� ��  .6 �  .6      E  , , �}  )� �}  *N �E  *N �E  )� �}  )�      E  , , �  )� �  *N ��  *N ��  )� �  )�      E  , , ��  )� ��  *N �}  *N �}  )� ��  )�      E  , , �Q  )� �Q  *N �  *N �  )� �Q  )�      E  , , ��  )� ��  *N ��  *N ��  )� ��  )�      E  , , ��  .6 ��  .� �}  .� �}  .6 ��  .6      E  , , �Q  .6 �Q  .� �  .� �  .6 �Q  .6      E  , , ��  .6 ��  .� ��  .� ��  .6 ��  .6      E  , , �  /� �  0� ��  0� ��  /� �  /�      E  , , ��  /� ��  0� �}  0� �}  /� ��  /�      E  , , �}  2� �}  3� �E  3� �E  2� �}  2�      E  , , �}  1V �}  2 �E  2 �E  1V �}  1V      E  , , �  1V �  2 ��  2 ��  1V �  1V      E  , , ��  1V ��  2 �}  2 �}  1V ��  1V      E  , , �Q  1V �Q  2 �  2 �  1V �Q  1V      E  , , �}  ! �}  !� �E  !� �E  ! �}  !      E  , , �  ! �  !� ��  !� ��  ! �  !      E  , , ��  ! ��  !� �}  !� �}  ! ��  !      E  , , �Q  ! �Q  !� �  !� �  ! �Q  !      E  , , ��  ! ��  !� ��  !� ��  ! ��  !      E  , , �  "� �  #Z ��  #Z ��  "� �  "�      E  , , �}  r �}   : �E   : �E  r �}  r      E  , , �  r �   : ��   : ��  r �  r      E  , , ��  r ��   : �}   : �}  r ��  r      E  , , �Q  r �Q   : �   : �  r �Q  r      E  , , ��  r ��   : ��   : ��  r ��  r      E  , , ��  "� ��  #Z �}  #Z �}  "� ��  "�      E  , , �}  � �}  � �E  � �E  � �}  �      E  , , �  � �  � ��  � ��  � �  �      E  , , ��  � ��  � �}  � �}  � ��  �      E  , , �Q  � �Q  � �  � �  � �Q  �      E  , , ��  � ��  � ��  � ��  � ��  �      E  , , �Q  "� �Q  #Z �  #Z �  "� �Q  "�      E  , , �}  R �}   �E   �E  R �}  R      E  , , �  R �   ��   ��  R �  R      E  , , ��  R ��   �}   �}  R ��  R      E  , , �Q  R �Q   �   �  R �Q  R      E  , , ��  R ��   ��   ��  R ��  R      E  , , ��  "� ��  #Z ��  #Z ��  "� ��  "�      E  , , �}  � �}  � �E  � �E  � �}  �      E  , , �  � �  � ��  � ��  � �  �      E  , , ��  � ��  � �}  � �}  � ��  �      E  , , �Q  � �Q  � �  � �  � �Q  �      E  , , ��  � ��  � ��  � ��  � ��  �      E  , , �}  "� �}  #Z �E  #Z �E  "� �}  "�      E  , , �}  2 �}  � �E  � �E  2 �}  2      E  , , �  2 �  � ��  � ��  2 �  2      E  , , ��  2 ��  � �}  � �}  2 ��  2      E  , , �Q  2 �Q  � �  � �  2 �Q  2      E  , , ��  2 ��  � ��  � ��  2 ��  2      E  , , ŉ  R ŉ   �Q   �Q  R ŉ  R      E  , , �%  R �%   ��   ��  R �%  R      E  , , ��  R ��   ω   ω  R ��  R      E  , , ŉ  ! ŉ  !� �Q  !� �Q  ! ŉ  !      E  , , �%  ! �%  !� ��  !� ��  ! �%  !      E  , , ��  ! ��  !� ω  !� ω  ! ��  !      E  , , ŉ  � ŉ  � �Q  � �Q  � ŉ  �      E  , , �%  � �%  � ��  � ��  � �%  �      E  , , ��  � ��  � ω  � ω  � ��  �      E  , , ŉ  � ŉ  � �Q  � �Q  � ŉ  �      E  , , �%  � �%  � ��  � ��  � �%  �      E  , , ��  � ��  � ω  � ω  � ��  �      E  , , ŉ  r ŉ   : �Q   : �Q  r ŉ  r      E  , , �%  r �%   : ��   : ��  r �%  r      E  , , ��  r ��   : ω   : ω  r ��  r      E  , , ŉ  "� ŉ  #Z �Q  #Z �Q  "� ŉ  "�      E  , , �%  "� �%  #Z ��  #Z ��  "� �%  "�      E  , , ��  "� ��  #Z ω  #Z ω  "� ��  "�      E  , , ŉ  2 ŉ  � �Q  � �Q  2 ŉ  2      E  , , �%  2 �%  � ��  � ��  2 �%  2      E  , , ��  2 ��  � ω  � ω  2 ��  2      E  , , �  + �  +� ��  +� ��  + �  +      E  , , ��  + ��  +� �q  +� �q  + ��  +      E  , , �E  + �E  +� �  +� �  + �E  +      E  , , �  .6 �  .� ��  .� ��  .6 �  .6      E  , , ��  .6 ��  .� �q  .� �q  .6 ��  .6      E  , , �E  .6 �E  .� �  .� �  .6 �E  .6      E  , , y�  r y�   : zf   : zf  r y�  r      E  , , ~:  r ~:   :    :   r ~:  r      E  , , �q  r �q   : �9   : �9  r �q  r      E  , , �  r �   : ��   : ��  r �  r      E  , , ��  r ��   : �q   : �q  r ��  r      E  , , �E  r �E   : �   : �  r �E  r      E  , , y�  /� y�  0� zf  0� zf  /� y�  /�      E  , , ~:  /� ~:  0�   0�   /� ~:  /�      E  , , �q  /� �q  0� �9  0� �9  /� �q  /�      E  , , �  /� �  0� ��  0� ��  /� �  /�      E  , , ��  /� ��  0� �q  0� �q  /� ��  /�      E  , , �E  /� �E  0� �  0� �  /� �E  /�      E  , , y�  )� y�  *N zf  *N zf  )� y�  )�      E  , , ~:  )� ~:  *N   *N   )� ~:  )�      E  , , �q  )� �q  *N �9  *N �9  )� �q  )�      E  , , y�  � y�  � zf  � zf  � y�  �      E  , , ~:  � ~:  �   �   � ~:  �      E  , , �q  � �q  � �9  � �9  � �q  �      E  , , �  � �  � ��  � ��  � �  �      E  , , ��  � ��  � �q  � �q  � ��  �      E  , , �E  � �E  � �  � �  � �E  �      E  , , �  )� �  *N ��  *N ��  )� �  )�      E  , , ��  )� ��  *N �q  *N �q  )� ��  )�      E  , , �E  )� �E  *N �  *N �  )� �E  )�      E  , , �  2� �  3� ��  3� ��  2� �  2�      E  , , ��  2� ��  3� �q  3� �q  2� ��  2�      E  , , �E  2� �E  3� �  3� �  2� �E  2�      E  , , y�  ,� y�  -n zf  -n zf  ,� y�  ,�      E  , , ~:  ,� ~:  -n   -n   ,� ~:  ,�      E  , , �q  ,� �q  -n �9  -n �9  ,� �q  ,�      E  , , y�  R y�   zf   zf  R y�  R      E  , , ~:  R ~:        R ~:  R      E  , , �q  R �q   �9   �9  R �q  R      E  , , �  R �   ��   ��  R �  R      E  , , ��  R ��   �q   �q  R ��  R      E  , , �E  R �E   �   �  R �E  R      E  , , �  ,� �  -n ��  -n ��  ,� �  ,�      E  , , ��  ,� ��  -n �q  -n �q  ,� ��  ,�      E  , , �E  ,� �E  -n �  -n �  ,� �E  ,�      E  , , y�  "� y�  #Z zf  #Z zf  "� y�  "�      E  , , ~:  "� ~:  #Z   #Z   "� ~:  "�      E  , , �q  "� �q  #Z �9  #Z �9  "� �q  "�      E  , , �  "� �  #Z ��  #Z ��  "� �  "�      E  , , ��  "� ��  #Z �q  #Z �q  "� ��  "�      E  , , �E  "� �E  #Z �  #Z �  "� �E  "�      E  , , y�  � y�  � zf  � zf  � y�  �      E  , , ~:  � ~:  �   �   � ~:  �      E  , , �q  � �q  � �9  � �9  � �q  �      E  , , �  � �  � ��  � ��  � �  �      E  , , ��  � ��  � �q  � �q  � ��  �      E  , , �E  � �E  � �  � �  � �E  �      E  , , y�  1V y�  2 zf  2 zf  1V y�  1V      E  , , ~:  1V ~:  2   2   1V ~:  1V      E  , , �q  1V �q  2 �9  2 �9  1V �q  1V      E  , , �  1V �  2 ��  2 ��  1V �  1V      E  , , ��  1V ��  2 �q  2 �q  1V ��  1V      E  , , �E  1V �E  2 �  2 �  1V �E  1V      E  , , y�  .6 y�  .� zf  .� zf  .6 y�  .6      E  , , ~:  .6 ~:  .�   .�   .6 ~:  .6      E  , , �q  .6 �q  .� �9  .� �9  .6 �q  .6      E  , , y�  2 y�  � zf  � zf  2 y�  2      E  , , ~:  2 ~:  �   �   2 ~:  2      E  , , �q  2 �q  � �9  � �9  2 �q  2      E  , , �  2 �  � ��  � ��  2 �  2      E  , , ��  2 ��  � �q  � �q  2 ��  2      E  , , �E  2 �E  � �  � �  2 �E  2      E  , , y�  ! y�  !� zf  !� zf  ! y�  !      E  , , ~:  ! ~:  !�   !�   ! ~:  !      E  , , �q  ! �q  !� �9  !� �9  ! �q  !      E  , , �  ! �  !� ��  !� ��  ! �  !      E  , , ��  ! ��  !� �q  !� �q  ! ��  !      E  , , �E  ! �E  !� �  !� �  ! �E  !      E  , , y�  + y�  +� zf  +� zf  + y�  +      E  , , ~:  + ~:  +�   +�   + ~:  +      E  , , �q  + �q  +� �9  +� �9  + �q  +      E  , , y�  2� y�  3� zf  3� zf  2� y�  2�      E  , , ~:  2� ~:  3�   3�   2� ~:  2�      E  , , �q  2� �q  3� �9  3� �9  2� �q  2�      E  , , b�  /� b�  0� cZ  0� cZ  /� b�  /�      E  , , b�  ,� b�  -n cZ  -n cZ  ,� b�  ,�      E  , , g.  ,� g.  -n g�  -n g�  ,� g.  ,�      E  , , k�  ,� k�  -n l�  -n l�  ,� k�  ,�      E  , , pf  ,� pf  -n q.  -n q.  ,� pf  ,�      E  , , u  ,� u  -n u�  -n u�  ,� u  ,�      E  , , g.  /� g.  0� g�  0� g�  /� g.  /�      E  , , k�  /� k�  0� l�  0� l�  /� k�  /�      E  , , pf  /� pf  0� q.  0� q.  /� pf  /�      E  , , u  /� u  0� u�  0� u�  /� u  /�      E  , , pf  1V pf  2 q.  2 q.  1V pf  1V      E  , , u  1V u  2 u�  2 u�  1V u  1V      E  , , b�  + b�  +� cZ  +� cZ  + b�  +      E  , , g.  + g.  +� g�  +� g�  + g.  +      E  , , k�  + k�  +� l�  +� l�  + k�  +      E  , , pf  + pf  +� q.  +� q.  + pf  +      E  , , u  + u  +� u�  +� u�  + u  +      E  , , b�  1V b�  2 cZ  2 cZ  1V b�  1V      E  , , b�  )� b�  *N cZ  *N cZ  )� b�  )�      E  , , g.  )� g.  *N g�  *N g�  )� g.  )�      E  , , k�  )� k�  *N l�  *N l�  )� k�  )�      E  , , pf  )� pf  *N q.  *N q.  )� pf  )�      E  , , u  )� u  *N u�  *N u�  )� u  )�      E  , , b�  .6 b�  .� cZ  .� cZ  .6 b�  .6      E  , , g.  .6 g.  .� g�  .� g�  .6 g.  .6      E  , , k�  .6 k�  .� l�  .� l�  .6 k�  .6      E  , , pf  .6 pf  .� q.  .� q.  .6 pf  .6      E  , , u  .6 u  .� u�  .� u�  .6 u  .6      E  , , g.  1V g.  2 g�  2 g�  1V g.  1V      E  , , k�  1V k�  2 l�  2 l�  1V k�  1V      E  , , b�  2� b�  3� cZ  3� cZ  2� b�  2�      E  , , g.  2� g.  3� g�  3� g�  2� g.  2�      E  , , k�  2� k�  3� l�  3� l�  2� k�  2�      E  , , pf  2� pf  3� q.  3� q.  2� pf  2�      E  , , u  2� u  3� u�  3� u�  2� u  2�      E  , , ]�  /� ]�  0� ^�  0� ^�  /� ]�  /�      E  , , K�  /� K�  0� LN  0� LN  /� K�  /�      E  , , T�  1V T�  2 U�  2 U�  1V T�  1V      E  , , YZ  1V YZ  2 Z"  2 Z"  1V YZ  1V      E  , , ]�  1V ]�  2 ^�  2 ^�  1V ]�  1V      E  , , F�  ,� F�  -n G�  -n G�  ,� F�  ,�      E  , , F�  .6 F�  .� G�  .� G�  .6 F�  .6      E  , , K�  .6 K�  .� LN  .� LN  .6 K�  .6      E  , , P"  .6 P"  .� P�  .� P�  .6 P"  .6      E  , , T�  .6 T�  .� U�  .� U�  .6 T�  .6      E  , , YZ  .6 YZ  .� Z"  .� Z"  .6 YZ  .6      E  , , F�  )� F�  *N G�  *N G�  )� F�  )�      E  , , K�  )� K�  *N LN  *N LN  )� K�  )�      E  , , P"  )� P"  *N P�  *N P�  )� P"  )�      E  , , T�  )� T�  *N U�  *N U�  )� T�  )�      E  , , YZ  )� YZ  *N Z"  *N Z"  )� YZ  )�      E  , , ]�  )� ]�  *N ^�  *N ^�  )� ]�  )�      E  , , K�  ,� K�  -n LN  -n LN  ,� K�  ,�      E  , , P"  ,� P"  -n P�  -n P�  ,� P"  ,�      E  , , T�  ,� T�  -n U�  -n U�  ,� T�  ,�      E  , , YZ  ,� YZ  -n Z"  -n Z"  ,� YZ  ,�      E  , , ]�  ,� ]�  -n ^�  -n ^�  ,� ]�  ,�      E  , , ]�  .6 ]�  .� ^�  .� ^�  .6 ]�  .6      E  , , F�  1V F�  2 G�  2 G�  1V F�  1V      E  , , K�  1V K�  2 LN  2 LN  1V K�  1V      E  , , P"  1V P"  2 P�  2 P�  1V P"  1V      E  , , F�  + F�  +� G�  +� G�  + F�  +      E  , , K�  + K�  +� LN  +� LN  + K�  +      E  , , P"  + P"  +� P�  +� P�  + P"  +      E  , , T�  + T�  +� U�  +� U�  + T�  +      E  , , F�  /� F�  0� G�  0� G�  /� F�  /�      E  , , F�  2� F�  3� G�  3� G�  2� F�  2�      E  , , K�  2� K�  3� LN  3� LN  2� K�  2�      E  , , P"  2� P"  3� P�  3� P�  2� P"  2�      E  , , T�  2� T�  3� U�  3� U�  2� T�  2�      E  , , YZ  2� YZ  3� Z"  3� Z"  2� YZ  2�      E  , , ]�  2� ]�  3� ^�  3� ^�  2� ]�  2�      E  , , YZ  + YZ  +� Z"  +� Z"  + YZ  +      E  , , ]�  + ]�  +� ^�  +� ^�  + ]�  +      E  , , P"  /� P"  0� P�  0� P�  /� P"  /�      E  , , T�  /� T�  0� U�  0� U�  /� T�  /�      E  , , YZ  /� YZ  0� Z"  0� Z"  /� YZ  /�      E  , , K�  � K�  � LN  � LN  � K�  �      E  , , P"  � P"  � P�  � P�  � P"  �      E  , , T�  � T�  � U�  � U�  � T�  �      E  , , YZ  � YZ  � Z"  � Z"  � YZ  �      E  , , ]�  � ]�  � ^�  � ^�  � ]�  �      E  , , K�  � K�  � LN  � LN  � K�  �      E  , , P"  � P"  � P�  � P�  � P"  �      E  , , T�  � T�  � U�  � U�  � T�  �      E  , , YZ  � YZ  � Z"  � Z"  � YZ  �      E  , , ]�  � ]�  � ^�  � ^�  � ]�  �      E  , , F�  ! F�  !� G�  !� G�  ! F�  !      E  , , K�  ! K�  !� LN  !� LN  ! K�  !      E  , , P"  ! P"  !� P�  !� P�  ! P"  !      E  , , T�  ! T�  !� U�  !� U�  ! T�  !      E  , , YZ  ! YZ  !� Z"  !� Z"  ! YZ  !      E  , , ]�  ! ]�  !� ^�  !� ^�  ! ]�  !      E  , , T�  "� T�  #Z U�  #Z U�  "� T�  "�      E  , , YZ  "� YZ  #Z Z"  #Z Z"  "� YZ  "�      E  , , F�  r F�   : G�   : G�  r F�  r      E  , , F�  2 F�  � G�  � G�  2 F�  2      E  , , K�  2 K�  � LN  � LN  2 K�  2      E  , , P"  2 P"  � P�  � P�  2 P"  2      E  , , T�  2 T�  � U�  � U�  2 T�  2      E  , , YZ  2 YZ  � Z"  � Z"  2 YZ  2      E  , , ]�  2 ]�  � ^�  � ^�  2 ]�  2      E  , , K�  r K�   : LN   : LN  r K�  r      E  , , P"  r P"   : P�   : P�  r P"  r      E  , , T�  r T�   : U�   : U�  r T�  r      E  , , YZ  r YZ   : Z"   : Z"  r YZ  r      E  , , ]�  r ]�   : ^�   : ^�  r ]�  r      E  , , F�  R F�   G�   G�  R F�  R      E  , , K�  R K�   LN   LN  R K�  R      E  , , P"  R P"   P�   P�  R P"  R      E  , , T�  R T�   U�   U�  R T�  R      E  , , YZ  R YZ   Z"   Z"  R YZ  R      E  , , ]�  R ]�   ^�   ^�  R ]�  R      E  , , ]�  "� ]�  #Z ^�  #Z ^�  "� ]�  "�      E  , , F�  "� F�  #Z G�  #Z G�  "� F�  "�      E  , , K�  "� K�  #Z LN  #Z LN  "� K�  "�      E  , , P"  "� P"  #Z P�  #Z P�  "� P"  "�      E  , , F�  � F�  � G�  � G�  � F�  �      E  , , F�  � F�  � G�  � G�  � F�  �      E  , , pf  � pf  � q.  � q.  � pf  �      E  , , u  � u  � u�  � u�  � u  �      E  , , b�  R b�   cZ   cZ  R b�  R      E  , , g.  R g.   g�   g�  R g.  R      E  , , k�  R k�   l�   l�  R k�  R      E  , , pf  R pf   q.   q.  R pf  R      E  , , u  R u   u�   u�  R u  R      E  , , b�  r b�   : cZ   : cZ  r b�  r      E  , , g.  r g.   : g�   : g�  r g.  r      E  , , k�  r k�   : l�   : l�  r k�  r      E  , , pf  r pf   : q.   : q.  r pf  r      E  , , u  r u   : u�   : u�  r u  r      E  , , b�  "� b�  #Z cZ  #Z cZ  "� b�  "�      E  , , b�  2 b�  � cZ  � cZ  2 b�  2      E  , , g.  2 g.  � g�  � g�  2 g.  2      E  , , k�  2 k�  � l�  � l�  2 k�  2      E  , , pf  2 pf  � q.  � q.  2 pf  2      E  , , u  2 u  � u�  � u�  2 u  2      E  , , g.  "� g.  #Z g�  #Z g�  "� g.  "�      E  , , k�  "� k�  #Z l�  #Z l�  "� k�  "�      E  , , pf  "� pf  #Z q.  #Z q.  "� pf  "�      E  , , u  "� u  #Z u�  #Z u�  "� u  "�      E  , , b�  ! b�  !� cZ  !� cZ  ! b�  !      E  , , b�  � b�  � cZ  � cZ  � b�  �      E  , , g.  � g.  � g�  � g�  � g.  �      E  , , k�  � k�  � l�  � l�  � k�  �      E  , , pf  � pf  � q.  � q.  � pf  �      E  , , u  � u  � u�  � u�  � u  �      E  , , g.  ! g.  !� g�  !� g�  ! g.  !      E  , , k�  ! k�  !� l�  !� l�  ! k�  !      E  , , pf  ! pf  !� q.  !� q.  ! pf  !      E  , , u  ! u  !� u�  !� u�  ! u  !      E  , , b�  � b�  � cZ  � cZ  � b�  �      E  , , g.  � g.  � g�  � g�  � g.  �      E  , , k�  � k�  � l�  � l�  � k�  �      E  , , �  � �  � o  � o  � �  �      E  , , C  � C  �   �   � C  �      E  , , �  � �  �  �  �  �  � �  �      E  , , ${  � ${  � %C  � %C  � ${  �      E  , , )  � )  � )�  � )�  � )  �      E  , , -�  � -�  � .{  � .{  � -�  �      E  , , -�  ,� -�  -n .{  -n .{  ,� -�  ,�      E  , , �  ,� �  -n o  -n o  ,� �  ,�      E  , , C  ,� C  -n   -n   ,� C  ,�      E  , , �  ,� �  -n  �  -n  �  ,� �  ,�      E  , , �  ! �  !� o  !� o  ! �  !      E  , , C  ! C  !�   !�   ! C  !      E  , , �  ! �  !�  �  !�  �  ! �  !      E  , , ${  ! ${  !� %C  !� %C  ! ${  !      E  , , )  ! )  !� )�  !� )�  ! )  !      E  , , -�  ! -�  !� .{  !� .{  ! -�  !      E  , , C  1V C  2   2   1V C  1V      E  , , -�  )� -�  *N .{  *N .{  )� -�  )�      E  , , �  1V �  2  �  2  �  1V �  1V      E  , , ${  1V ${  2 %C  2 %C  1V ${  1V      E  , , )  1V )  2 )�  2 )�  1V )  1V      E  , , -�  1V -�  2 .{  2 .{  1V -�  1V      E  , , ${  ,� ${  -n %C  -n %C  ,� ${  ,�      E  , , �  1V �  2 o  2 o  1V �  1V      E  , , �  r �   : o   : o  r �  r      E  , , �  + �  +� o  +� o  + �  +      E  , , C  + C  +�   +�   + C  +      E  , , �  .6 �  .� o  .� o  .6 �  .6      E  , , �  R �   o   o  R �  R      E  , , C  R C        R C  R      E  , , �  R �    �    �  R �  R      E  , , ${  R ${   %C   %C  R ${  R      E  , , �  2 �  � o  � o  2 �  2      E  , , C  2 C  �   �   2 C  2      E  , , �  2 �  �  �  �  �  2 �  2      E  , , ${  2 ${  � %C  � %C  2 ${  2      E  , , )  2 )  � )�  � )�  2 )  2      E  , , -�  2 -�  � .{  � .{  2 -�  2      E  , , )  R )   )�   )�  R )  R      E  , , -�  R -�   .{   .{  R -�  R      E  , , �  + �  +�  �  +�  �  + �  +      E  , , ${  + ${  +� %C  +� %C  + ${  +      E  , , )  + )  +� )�  +� )�  + )  +      E  , , -�  + -�  +� .{  +� .{  + -�  +      E  , , C  r C   :    :   r C  r      E  , , �  � �  � o  � o  � �  �      E  , , C  � C  �   �   � C  �      E  , , �  � �  �  �  �  �  � �  �      E  , , ${  � ${  � %C  � %C  � ${  �      E  , , )  � )  � )�  � )�  � )  �      E  , , -�  � -�  � .{  � .{  � -�  �      E  , , C  .6 C  .�   .�   .6 C  .6      E  , , �  .6 �  .�  �  .�  �  .6 �  .6      E  , , ${  .6 ${  .� %C  .� %C  .6 ${  .6      E  , , �  /� �  0� o  0� o  /� �  /�      E  , , C  /� C  0�   0�   /� C  /�      E  , , �  /� �  0�  �  0�  �  /� �  /�      E  , , ${  /� ${  0� %C  0� %C  /� ${  /�      E  , , )  /� )  0� )�  0� )�  /� )  /�      E  , , -�  /� -�  0� .{  0� .{  /� -�  /�      E  , , )  .6 )  .� )�  .� )�  .6 )  .6      E  , , �  "� �  #Z o  #Z o  "� �  "�      E  , , C  "� C  #Z   #Z   "� C  "�      E  , , �  "� �  #Z  �  #Z  �  "� �  "�      E  , , �  2� �  3� o  3� o  2� �  2�      E  , , C  2� C  3�   3�   2� C  2�      E  , , �  2� �  3�  �  3�  �  2� �  2�      E  , , ${  2� ${  3� %C  3� %C  2� ${  2�      E  , , )  2� )  3� )�  3� )�  2� )  2�      E  , , -�  2� -�  3� .{  3� .{  2� -�  2�      E  , , -�  .6 -�  .� .{  .� .{  .6 -�  .6      E  , , �  r �   :  �   :  �  r �  r      E  , , ${  r ${   : %C   : %C  r ${  r      E  , , )  r )   : )�   : )�  r )  r      E  , , -�  r -�   : .{   : .{  r -�  r      E  , , )  ,� )  -n )�  -n )�  ,� )  ,�      E  , , �  )� �  *N o  *N o  )� �  )�      E  , , C  )� C  *N   *N   )� C  )�      E  , , �  )� �  *N  �  *N  �  )� �  )�      E  , , ${  )� ${  *N %C  *N %C  )� ${  )�      E  , , )  )� )  *N )�  *N )�  )� )  )�      E  , , ${  "� ${  #Z %C  #Z %C  "� ${  "�      E  , , )  "� )  #Z )�  #Z )�  "� )  "�      E  , , -�  "� -�  #Z .{  #Z .{  "� -�  "�      E  , ,  �c  �  �c  �  �+  �  �+  �  �c  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  ��  �  ��  �  c  �  c  �  ��  �      E  , , 7  � 7  � �  � �  � 7  �      E  , , �  � �  � 	�  � 	�  � �  �      E  , , o  � o  � 7  � 7  � o  �      E  , ,   �   � �  � �  �   �      E  , ,  ��  !  ��  !�  c  !�  c  !  ��  !      E  , , 7  ! 7  !� �  !� �  ! 7  !      E  , , �  ! �  !� 	�  !� 	�  ! �  !      E  , , o  ! o  !� 7  !� 7  ! o  !      E  , ,   !   !� �  !� �  !   !      E  , , 7  /� 7  0� �  0� �  /� 7  /�      E  , ,  �c  �  �c  �  �+  �  �+  �  �c  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  ��  �  ��  �  c  �  c  �  ��  �      E  , , 7  � 7  � �  � �  � 7  �      E  , , �  � �  � 	�  � 	�  � �  �      E  , , o  � o  � 7  � 7  � o  �      E  , ,   �   � �  � �  �   �      E  , , �  /� �  0� 	�  0� 	�  /� �  /�      E  , , o  /� o  0� 7  0� 7  /� o  /�      E  , ,   /�   0� �  0� �  /�   /�      E  , ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      E  , ,  ��  2�  ��  3�  c  3�  c  2�  ��  2�      E  , , 7  2� 7  3� �  3� �  2� 7  2�      E  , ,  �c  1V  �c  2  �+  2  �+  1V  �c  1V      E  , ,  ��  1V  ��  2  ��  2  ��  1V  ��  1V      E  , ,  ��  1V  ��  2  c  2  c  1V  ��  1V      E  , , 7  1V 7  2 �  2 �  1V 7  1V      E  , , �  1V �  2 	�  2 	�  1V �  1V      E  , , o  1V o  2 7  2 7  1V o  1V      E  , ,   1V   2 �  2 �  1V   1V      E  , , �  2� �  3� 	�  3� 	�  2� �  2�      E  , ,  �c  .6  �c  .�  �+  .�  �+  .6  �c  .6      E  , ,  ��  .6  ��  .�  ��  .�  ��  .6  ��  .6      E  , ,  �c  "�  �c  #Z  �+  #Z  �+  "�  �c  "�      E  , ,  ��  "�  ��  #Z  ��  #Z  ��  "�  ��  "�      E  , ,  ��  "�  ��  #Z  c  #Z  c  "�  ��  "�      E  , ,  �c  2  �c  �  �+  �  �+  2  �c  2      E  , ,  ��  2  ��  �  ��  �  ��  2  ��  2      E  , ,  ��  2  ��  �  c  �  c  2  ��  2      E  , , 7  2 7  � �  � �  2 7  2      E  , , �  2 �  � 	�  � 	�  2 �  2      E  , , o  2 o  � 7  � 7  2 o  2      E  , ,   2   � �  � �  2   2      E  , , 7  "� 7  #Z �  #Z �  "� 7  "�      E  , , �  "� �  #Z 	�  #Z 	�  "� �  "�      E  , , o  "� o  #Z 7  #Z 7  "� o  "�      E  , ,   "�   #Z �  #Z �  "�   "�      E  , ,  ��  .6  ��  .�  c  .�  c  .6  ��  .6      E  , , 7  .6 7  .� �  .� �  .6 7  .6      E  , , �  .6 �  .� 	�  .� 	�  .6 �  .6      E  , , o  .6 o  .� 7  .� 7  .6 o  .6      E  , ,   .6   .� �  .� �  .6   .6      E  , , o  2� o  3� 7  3� 7  2� o  2�      E  , ,   2�   3� �  3� �  2�   2�      E  , ,  �c  2�  �c  3�  �+  3�  �+  2�  �c  2�      E  , ,  �c  r  �c   :  �+   :  �+  r  �c  r      E  , ,  �c  R  �c    �+    �+  R  �c  R      E  , ,  ��  R  ��    ��    ��  R  ��  R      E  , ,  ��  R  ��    c    c  R  ��  R      E  , , 7  R 7   �   �  R 7  R      E  , , �  R �   	�   	�  R �  R      E  , , o  R o   7   7  R o  R      E  , ,   R    �   �  R   R      E  , ,  ��  r  ��   :  ��   :  ��  r  ��  r      E  , ,  ��  r  ��   :  c   :  c  r  ��  r      E  , , 7  r 7   : �   : �  r 7  r      E  , , �  r �   : 	�   : 	�  r �  r      E  , , o  r o   : 7   : 7  r o  r      E  , ,   r    : �   : �  r   r      E  , ,  �c  /�  �c  0�  �+  0�  �+  /�  �c  /�      E  , ,  �c  ,�  �c  -n  �+  -n  �+  ,�  �c  ,�      E  , ,  �c  )�  �c  *N  �+  *N  �+  )�  �c  )�      E  , ,  ��  )�  ��  *N  ��  *N  ��  )�  ��  )�      E  , ,  ��  )�  ��  *N  c  *N  c  )�  ��  )�      E  , , 7  )� 7  *N �  *N �  )� 7  )�      E  , , �  )� �  *N 	�  *N 	�  )� �  )�      E  , , o  )� o  *N 7  *N 7  )� o  )�      E  , ,   )�   *N �  *N �  )�   )�      E  , ,  ��  ,�  ��  -n  ��  -n  ��  ,�  ��  ,�      E  , ,  ��  ,�  ��  -n  c  -n  c  ,�  ��  ,�      E  , , 7  ,� 7  -n �  -n �  ,� 7  ,�      E  , ,  �c  +  �c  +�  �+  +�  �+  +  �c  +      E  , ,  ��  +  ��  +�  ��  +�  ��  +  ��  +      E  , ,  ��  +  ��  +�  c  +�  c  +  ��  +      E  , , 7  + 7  +� �  +� �  + 7  +      E  , , �  + �  +� 	�  +� 	�  + �  +      E  , , o  + o  +� 7  +� 7  + o  +      E  , ,   +   +� �  +� �  +   +      E  , , �  ,� �  -n 	�  -n 	�  ,� �  ,�      E  , , o  ,� o  -n 7  -n 7  ,� o  ,�      E  , ,   ,�   -n �  -n �  ,�   ,�      E  , ,  ��  /�  ��  0�  ��  0�  ��  /�  ��  /�      E  , ,  ��  /�  ��  0�  c  0�  c  /�  ��  /�      E  , ,  �c  !  �c  !�  �+  !�  �+  !  �c  !      E  , ,  ��  !  ��  !�  ��  !�  ��  !  ��  !      E  , ,  ��  �  ��  V  Ϗ  V  Ϗ  �  ��  �      E  , ,  �  �  �  �  ��  �  ��  �  �  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  �W  �  �W  �  �  �  �  �  �W  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  ŏ  �  ŏ  �  �W  �  �W  �  ŏ  �      E  , ,  �+  �  �+  �  ��  �  ��  �  �+  �      E  , ,  ��  �  ��  �  Ϗ  �  Ϗ  �  ��  �      E  , ,  �  n  �  6  ��  6  ��  n  �  n      E  , ,  ��  n  ��  6  ��  6  ��  n  ��  n      E  , ,  �W  n  �W  6  �  6  �  n  �W  n      E  , ,  ��  n  ��  6  ��  6  ��  n  ��  n      E  , ,  ŏ  n  ŏ  6  �W  6  �W  n  ŏ  n      E  , ,  �+  n  �+  6  ��  6  ��  n  �+  n      E  , ,  ��  n  ��  6  Ϗ  6  Ϗ  n  ��  n      E  , ,  �  �  �  �  ��  �  ��  �  �  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  �W  �  �W  �  �  �  �  �  �W  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  ŏ  �  ŏ  �  �W  �  �W  �  ŏ  �      E  , ,  �+  �  �+  �  ��  �  ��  �  �+  �      E  , ,  ��  �  ��  �  Ϗ  �  Ϗ  �  ��  �      E  , ,  �  N  �    ��    ��  N  �  N      E  , ,  ��  N  ��    ��    ��  N  ��  N      E  , ,  �W  N  �W    �    �  N  �W  N      E  , ,  ��  N  ��    ��    ��  N  ��  N      E  , ,  ŏ  N  ŏ    �W    �W  N  ŏ  N      E  , ,  �+  N  �+    ��    ��  N  �+  N      E  , ,  ��  N  ��    Ϗ    Ϗ  N  ��  N      E  , ,  �  Z  �  "  ��  "  ��  Z  �  Z      E  , ,  ��  Z  ��  "  ��  "  ��  Z  ��  Z      E  , ,  �W  Z  �W  "  �  "  �  Z  �W  Z      E  , ,  ��  Z  ��  "  ��  "  ��  Z  ��  Z      E  , ,  ŏ  Z  ŏ  "  �W  "  �W  Z  ŏ  Z      E  , ,  �+  Z  �+  "  ��  "  ��  Z  �+  Z      E  , ,  ��  Z  ��  "  Ϗ  "  Ϗ  Z  ��  Z      E  , ,  �  �  �  �  ��  �  ��  �  �  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  �W  �  �W  �  �  �  �  �  �W  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  ŏ  �  ŏ  �  �W  �  �W  �  ŏ  �      E  , ,  �+  �  �+  �  ��  �  ��  �  �+  �      E  , ,  ��  �  ��  �  Ϗ  �  Ϗ  �  ��  �      E  , ,  �  :  �    ��    ��  :  �  :      E  , ,  ��  :  ��    ��    ��  :  ��  :      E  , ,  �W  :  �W    �    �  :  �W  :      E  , ,  ��  :  ��    ��    ��  :  ��  :      E  , ,  ŏ  :  ŏ    �W    �W  :  ŏ  :      E  , ,  �+  :  �+    ��    ��  :  �+  :      E  , ,  ��  :  ��    Ϗ    Ϗ  :  ��  :      E  , ,  �   �  �  r  ��  r  ��   �  �   �      E  , ,  ��   �  ��  r  ��  r  ��   �  ��   �      E  , ,  �W   �  �W  r  �  r  �   �  �W   �      E  , ,  ��   �  ��  r  ��  r  ��   �  ��   �      E  , ,  ŏ   �  ŏ  r  �W  r  �W   �  ŏ   �      E  , ,  �+   �  �+  r  ��  r  ��   �  �+   �      E  , ,  ��   �  ��  r  Ϗ  r  Ϗ   �  ��   �      E  , ,  ����  �����  ������  �����  ����      E  , ,  �����  ������  ������  �����  �����      E  , ,  �W���  �W����  �����  ����  �W���      E  , ,  �����  ������  ������  �����  �����      E  , ,  ŏ���  ŏ����  �W����  �W���  ŏ���      E  , ,  �+���  �+����  ������  �����  �+���      E  , ,  �����  ������  Ϗ����  Ϗ���  �����      E  , ,  �����  ����R  �����R  ������  �����      E  , ,  ������  �����R  �����R  ������  ������      E  , ,  �W����  �W���R  ����R  �����  �W����      E  , ,  ������  �����R  �����R  ������  ������      E  , ,  ŏ����  ŏ���R  �W���R  �W����  ŏ����      E  , ,  �+����  �+���R  �����R  ������  �+����      E  , ,  ������  �����R  Ϗ���R  Ϗ����  ������      E  , ,  �����  �����  ������  ������  �����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �W����  �W����  �����  �����  �W����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ŏ����  ŏ����  �W����  �W����  ŏ����      E  , ,  �+����  �+����  ������  ������  �+����      E  , ,  ������  ������  Ϗ����  Ϗ����  ������      E  , ,  �  �  �  v  ��  v  ��  �  �  �      E  , ,  ��  �  ��  v  ��  v  ��  �  ��  �      E  , ,  �W  �  �W  v  �  v  �  �  �W  �      E  , ,  ��  �  ��  v  ��  v  ��  �  ��  �      E  , ,  ŏ  �  ŏ  v  �W  v  �W  �  ŏ  �      E  , ,  �+  �  �+  v  ��  v  ��  �  �+  �      E  , ,  ��  �  ��  v  Ϗ  v  Ϗ  �  ��  �      E  , ,  �    �  �  ��  �  ��    �        E  , ,  ��    ��  �  ��  �  ��    ��        E  , ,  �W    �W  �  �  �  �    �W        E  , ,  ��    ��  �  ��  �  ��    ��        E  , ,  ŏ    ŏ  �  �W  �  �W    ŏ        E  , ,  �+    �+  �  ��  �  ��    �+        E  , ,  ��    ��  �  Ϗ  �  Ϗ    ��        E  , ,  �  �  �  V  ��  V  ��  �  �  �      E  , ,  ��  �  ��  V  ��  V  ��  �  ��  �      E  , ,  �W  �  �W  V  �  V  �  �  �W  �      E  , ,  ��  �  ��  V  ��  V  ��  �  ��  �      E  , ,  ŏ  �  ŏ  V  �W  V  �W  �  ŏ  �      E  , ,  �+  �  �+  V  ��  V  ��  �  �+  �      E  , ,  m�    m�  �  n�  �  n�    m�        E  , ,  r�    r�  �  s_  �  s_    r�        E  , ,  w3    w3  �  w�  �  w�    w3        E  , ,  {�    {�  �  |�  �  |�    {�        E  , ,  `'  �  `'  �  `�  �  `�  �  `'  �      E  , ,  d�  �  d�  �  e�  �  e�  �  d�  �      E  , ,  i_  �  i_  �  j'  �  j'  �  i_  �      E  , ,  m�  �  m�  �  n�  �  n�  �  m�  �      E  , ,  r�  �  r�  �  s_  �  s_  �  r�  �      E  , ,  w3  �  w3  �  w�  �  w�  �  w3  �      E  , ,  {�  �  {�  �  |�  �  |�  �  {�  �      E  , ,  `'  N  `'    `�    `�  N  `'  N      E  , ,  d�  N  d�    e�    e�  N  d�  N      E  , ,  i_  N  i_    j'    j'  N  i_  N      E  , ,  m�  N  m�    n�    n�  N  m�  N      E  , ,  r�  N  r�    s_    s_  N  r�  N      E  , ,  w3  N  w3    w�    w�  N  w3  N      E  , ,  {�  N  {�    |�    |�  N  {�  N      E  , ,  `'  Z  `'  "  `�  "  `�  Z  `'  Z      E  , ,  d�  Z  d�  "  e�  "  e�  Z  d�  Z      E  , ,  i_  Z  i_  "  j'  "  j'  Z  i_  Z      E  , ,  m�  Z  m�  "  n�  "  n�  Z  m�  Z      E  , ,  r�  Z  r�  "  s_  "  s_  Z  r�  Z      E  , ,  w3  Z  w3  "  w�  "  w�  Z  w3  Z      E  , ,  {�  Z  {�  "  |�  "  |�  Z  {�  Z      E  , ,  `'  �  `'  V  `�  V  `�  �  `'  �      E  , ,  d�  �  d�  V  e�  V  e�  �  d�  �      E  , ,  i_  �  i_  V  j'  V  j'  �  i_  �      E  , ,  m�  �  m�  V  n�  V  n�  �  m�  �      E  , ,  r�  �  r�  V  s_  V  s_  �  r�  �      E  , ,  w3  �  w3  V  w�  V  w�  �  w3  �      E  , ,  `'  �  `'  �  `�  �  `�  �  `'  �      E  , ,  d�  �  d�  �  e�  �  e�  �  d�  �      E  , ,  i_  �  i_  �  j'  �  j'  �  i_  �      E  , ,  m�  �  m�  �  n�  �  n�  �  m�  �      E  , ,  r�  �  r�  �  s_  �  s_  �  r�  �      E  , ,  w3  �  w3  �  w�  �  w�  �  w3  �      E  , ,  {�  �  {�  �  |�  �  |�  �  {�  �      E  , ,  {�  �  {�  V  |�  V  |�  �  {�  �      E  , ,  `'  :  `'    `�    `�  :  `'  :      E  , ,  d�  :  d�    e�    e�  :  d�  :      E  , ,  i_  :  i_    j'    j'  :  i_  :      E  , ,  m�  :  m�    n�    n�  :  m�  :      E  , ,  r�  :  r�    s_    s_  :  r�  :      E  , ,  w3  :  w3    w�    w�  :  w3  :      E  , ,  {�  :  {�    |�    |�  :  {�  :      E  , ,  `'   �  `'  r  `�  r  `�   �  `'   �      E  , ,  d�   �  d�  r  e�  r  e�   �  d�   �      E  , ,  i_   �  i_  r  j'  r  j'   �  i_   �      E  , ,  m�   �  m�  r  n�  r  n�   �  m�   �      E  , ,  r�   �  r�  r  s_  r  s_   �  r�   �      E  , ,  w3   �  w3  r  w�  r  w�   �  w3   �      E  , ,  {�   �  {�  r  |�  r  |�   �  {�   �      E  , ,  `'  �  `'  v  `�  v  `�  �  `'  �      E  , ,  d�  �  d�  v  e�  v  e�  �  d�  �      E  , ,  i_  �  i_  v  j'  v  j'  �  i_  �      E  , ,  `'  �  `'  �  `�  �  `�  �  `'  �      E  , ,  d�  �  d�  �  e�  �  e�  �  d�  �      E  , ,  `'���  `'����  `�����  `����  `'���      E  , ,  d����  d�����  e�����  e����  d����      E  , ,  i_���  i_����  j'����  j'���  i_���      E  , ,  m����  m�����  n�����  n����  m����      E  , ,  r����  r�����  s_����  s_���  r����      E  , ,  w3���  w3����  w�����  w����  w3���      E  , ,  {����  {�����  |�����  |����  {����      E  , ,  i_  �  i_  �  j'  �  j'  �  i_  �      E  , ,  m�  �  m�  �  n�  �  n�  �  m�  �      E  , ,  r�  �  r�  �  s_  �  s_  �  r�  �      E  , ,  w3  �  w3  �  w�  �  w�  �  w3  �      E  , ,  {�  �  {�  �  |�  �  |�  �  {�  �      E  , ,  `'����  `'���R  `����R  `�����  `'����      E  , ,  d�����  d����R  e����R  e�����  d�����      E  , ,  i_����  i_���R  j'���R  j'����  i_����      E  , ,  m�����  m����R  n����R  n�����  m�����      E  , ,  r�����  r����R  s_���R  s_����  r�����      E  , ,  w3����  w3���R  w����R  w�����  w3����      E  , ,  {�����  {����R  |����R  |�����  {�����      E  , ,  `'����  `'����  `�����  `�����  `'����      E  , ,  d�����  d�����  e�����  e�����  d�����      E  , ,  i_����  i_����  j'����  j'����  i_����      E  , ,  m�����  m�����  n�����  n�����  m�����      E  , ,  r�����  r�����  s_����  s_����  r�����      E  , ,  w3����  w3����  w�����  w�����  w3����      E  , ,  {�����  {�����  |�����  |�����  {�����      E  , ,  m�  �  m�  v  n�  v  n�  �  m�  �      E  , ,  r�  �  r�  v  s_  v  s_  �  r�  �      E  , ,  w3  �  w3  v  w�  v  w�  �  w3  �      E  , ,  {�  �  {�  v  |�  v  |�  �  {�  �      E  , ,  `'    `'  �  `�  �  `�    `'        E  , ,  d�    d�  �  e�  �  e�    d�        E  , ,  i_    i_  �  j'  �  j'    i_        E  , ,  `'  n  `'  6  `�  6  `�  n  `'  n      E  , ,  d�  n  d�  6  e�  6  e�  n  d�  n      E  , ,  i_  n  i_  6  j'  6  j'  n  i_  n      E  , ,  m�  n  m�  6  n�  6  n�  n  m�  n      E  , ,  r�  n  r�  6  s_  6  s_  n  r�  n      E  , ,  w3  n  w3  6  w�  6  w�  n  w3  n      E  , ,  {�  n  {�  6  |�  6  |�  n  {�  n      E  , ,  �  N  �    ��    ��  N  �  N      E  , ,  �  �  �  V  ��  V  ��  �  �  �      E  , ,  ��  �  ��  V  �w  V  �w  �  ��  �      E  , ,  �K  �  �K  V  �  V  �  �  �K  �      E  , ,  ��  �  ��  V  ��  V  ��  �  ��  �      E  , ,  ��  �  ��  V  �K  V  �K  �  ��  �      E  , ,  ��  �  ��  v  �w  v  �w  �  ��  �      E  , ,  �K  �  �K  v  �  v  �  �  �K  �      E  , ,  ��  N  ��    �w    �w  N  ��  N      E  , ,  �K  N  �K    �    �  N  �K  N      E  , ,  ��  N  ��    ��    ��  N  ��  N      E  , ,  ��  N  ��    �K    �K  N  ��  N      E  , ,  ��    ��  �  �K  �  �K    ��        E  , ,  ��  �  ��  v  ��  v  ��  �  ��  �      E  , ,  ��  �  ��  v  �K  v  �K  �  ��  �      E  , ,  �  �  �  �  ��  �  ��  �  �  �      E  , ,  ��  �  ��  �  �w  �  �w  �  ��  �      E  , ,  �K  �  �K  �  �  �  �  �  �K  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  ��  �  ��  �  �K  �  �K  �  ��  �      E  , ,  �  �  �  v  ��  v  ��  �  �  �      E  , ,  �  �  �  �  ��  �  ��  �  �  �      E  , ,  ��  �  ��  �  �w  �  �w  �  ��  �      E  , ,  �K  �  �K  �  �  �  �  �  �K  �      E  , ,  �    �  �  ��  �  ��    �        E  , ,  ��    ��  �  �w  �  �w    ��        E  , ,  �K    �K  �  �  �  �    �K        E  , ,  ��    ��  �  ��  �  ��    ��        E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  ��  �  ��  �  �K  �  �K  �  ��  �      E  , ,  �  n  �  6  ��  6  ��  n  �  n      E  , ,  ��  n  ��  6  �w  6  �w  n  ��  n      E  , ,  �K  n  �K  6  �  6  �  n  �K  n      E  , ,  ��  n  ��  6  ��  6  ��  n  ��  n      E  , ,  ��  n  ��  6  �K  6  �K  n  ��  n      E  , ,  �w  �  �w  �  �?  �  �?  �  �w  �      E  , ,  �  �  �  V  ��  V  ��  �  �  �      E  , ,  ��  �  ��  V  �k  V  �k  �  ��  �      E  , ,  �?  �  �?  V  �  V  �  �  �?  �      E  , ,  ��  �  ��  V  ��  V  ��  �  ��  �      E  , ,  �w  �  �w  V  �?  V  �?  �  �w  �      E  , ,  �k  �  �k  �  �3  �  �3  �  �k  �      E  , ,  �  �  �  �  ��  �  ��  �  �  �      E  , ,  �k  N  �k    �3    �3  N  �k  N      E  , ,  �?    �?  �  �  �  �    �?        E  , ,  ��  �  ��  �  �k  �  �k  �  ��  �      E  , ,  �?  �  �?  �  �  �  �  �  �?  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  �w  �  �w  �  �?  �  �?  �  �w  �      E  , ,  �  N  �    ��    ��  N  �  N      E  , ,  ��  N  ��    �k    �k  N  ��  N      E  , ,  �?  N  �?    �    �  N  �?  N      E  , ,  ��    ��  �  ��  �  ��    ��        E  , ,  �w    �w  �  �?  �  �?    �w        E  , ,  ��  N  ��    ��    ��  N  ��  N      E  , ,  �w  N  �w    �?    �?  N  �w  N      E  , ,  �k  �  �k  v  �3  v  �3  �  �k  �      E  , ,  �  �  �  v  ��  v  ��  �  �  �      E  , ,  �    �  �  ��  �  ��    �        E  , ,  �?  �  �?  �  �  �  �  �  �?  �      E  , ,  �k  �  �k  V  �3  V  �3  �  �k  �      E  , ,  ��    ��  �  �k  �  �k    ��        E  , ,  �k    �k  �  �3  �  �3    �k        E  , ,  �k  �  �k  �  �3  �  �3  �  �k  �      E  , ,  �  �  �  �  ��  �  ��  �  �  �      E  , ,  ��  �  ��  �  �k  �  �k  �  ��  �      E  , ,  �k  n  �k  6  �3  6  �3  n  �k  n      E  , ,  �  n  �  6  ��  6  ��  n  �  n      E  , ,  ��  n  ��  6  �k  6  �k  n  ��  n      E  , ,  �?  n  �?  6  �  6  �  n  �?  n      E  , ,  ��  n  ��  6  ��  6  ��  n  ��  n      E  , ,  �w  n  �w  6  �?  6  �?  n  �w  n      E  , ,  ��  �  ��  v  �k  v  �k  �  ��  �      E  , ,  �?  �  �?  v  �  v  �  �  �?  �      E  , ,  ��  �  ��  v  ��  v  ��  �  ��  �      E  , ,  �w  �  �w  v  �?  v  �?  �  �w  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  �   �  �  r  ��  r  ��   �  �   �      E  , ,  ��   �  ��  r  �k  r  �k   �  ��   �      E  , ,  �?   �  �?  r  �  r  �   �  �?   �      E  , ,  ��   �  ��  r  ��  r  ��   �  ��   �      E  , ,  �w   �  �w  r  �?  r  �?   �  �w   �      E  , ,  ��  :  ��    �k    �k  :  ��  :      E  , ,  �k  Z  �k  "  �3  "  �3  Z  �k  Z      E  , ,  �k���  �k����  �3����  �3���  �k���      E  , ,  ����  �����  ������  �����  ����      E  , ,  �����  ������  �k����  �k���  �����      E  , ,  �?���  �?����  �����  ����  �?���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �k����  �k����  �3����  �3����  �k����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ������  ������  �k����  �k����  ������      E  , ,  �?����  �?����  �����  �����  �?����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �w����  �w����  �?����  �?����  �w����      E  , ,  �w���  �w����  �?����  �?���  �w���      E  , ,  �  Z  �  "  ��  "  ��  Z  �  Z      E  , ,  ��  Z  ��  "  �k  "  �k  Z  ��  Z      E  , ,  �?  Z  �?  "  �  "  �  Z  �?  Z      E  , ,  ��  Z  ��  "  ��  "  ��  Z  ��  Z      E  , ,  �w  Z  �w  "  �?  "  �?  Z  �w  Z      E  , ,  �?  :  �?    �    �  :  �?  :      E  , ,  �k  �  �k  �  �3  �  �3  �  �k  �      E  , ,  �  �  �  �  ��  �  ��  �  �  �      E  , ,  ��  �  ��  �  �k  �  �k  �  ��  �      E  , ,  �?  �  �?  �  �  �  �  �  �?  �      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  �w  �  �w  �  �?  �  �?  �  �w  �      E  , ,  ��  :  ��    ��    ��  :  ��  :      E  , ,  �w  :  �w    �?    �?  :  �w  :      E  , ,  �k  :  �k    �3    �3  :  �k  :      E  , ,  �k����  �k���R  �3���R  �3����  �k����      E  , ,  �����  ����R  �����R  ������  �����      E  , ,  ������  �����R  �k���R  �k����  ������      E  , ,  �?����  �?���R  ����R  �����  �?����      E  , ,  ������  �����R  �����R  ������  ������      E  , ,  �w����  �w���R  �?���R  �?����  �w����      E  , ,  �  :  �    ��    ��  :  �  :      E  , ,  �k   �  �k  r  �3  r  �3   �  �k   �      E  , ,  ��  :  ��    ��    ��  :  ��  :      E  , ,  �   �  �  r  ��  r  ��   �  �   �      E  , ,  ����  �����  ������  �����  ����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ������  ������  �w����  �w����  ������      E  , ,  �K����  �K����  �����  �����  �K����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �K����  �K����  ������      E  , ,  �����  ������  �w����  �w���  �����      E  , ,  �K���  �K����  �����  ����  �K���      E  , ,  �����  ����R  �����R  ������  �����      E  , ,  ������  �����R  �w���R  �w����  ������      E  , ,  �K����  �K���R  ����R  �����  �K����      E  , ,  ������  �����R  �����R  ������  ������      E  , ,  ������  �����R  �K���R  �K����  ������      E  , ,  �����  ������  ������  �����  �����      E  , ,  �����  ������  �K����  �K���  �����      E  , ,  ��   �  ��  r  �w  r  �w   �  ��   �      E  , ,  �K   �  �K  r  �  r  �   �  �K   �      E  , ,  ��   �  ��  r  ��  r  ��   �  ��   �      E  , ,  ��   �  ��  r  �K  r  �K   �  ��   �      E  , ,  �  �  �  �  ��  �  ��  �  �  �      E  , ,  ��  �  ��  �  �w  �  �w  �  ��  �      E  , ,  �K  �  �K  �  �  �  �  �  �K  �      E  , ,  ��  :  ��    �K    �K  :  ��  :      E  , ,  ��  �  ��  �  ��  �  ��  �  ��  �      E  , ,  ��  �  ��  �  �K  �  �K  �  ��  �      E  , ,  �  Z  �  "  ��  "  ��  Z  �  Z      E  , ,  ��  Z  ��  "  �w  "  �w  Z  ��  Z      E  , ,  �K  Z  �K  "  �  "  �  Z  �K  Z      E  , ,  ��  Z  ��  "  ��  "  ��  Z  ��  Z      E  , ,  ��  Z  ��  "  �K  "  �K  Z  ��  Z      E  , ,  �  :  �    ��    ��  :  �  :      E  , ,  ��  :  ��    �w    �w  :  ��  :      E  , ,  �K  :  �K    �    �  :  �K  :      E  , ,  �k���  �k����  �3����  �3���  �k���      E  , ,  ����  �����  ������  �����  ����      E  , ,  �����  ������  �k����  �k���  �����      E  , ,  �?���  �?����  �����  ����  �?���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �w���  �w����  �?����  �?���  �w���      E  , ,  ����  �����  ������  �����  ����      E  , ,  �����  ������  �w����  �w���  �����      E  , ,  �K���  �K����  �����  ����  �K���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �����  ������  �K����  �K���  �����      E  , ,  �k���  �k���L  �3���L  �3���  �k���      E  , ,  ����  ����L  �����L  �����  ����      E  , ,  �����  �����L  �k���L  �k���  �����      E  , ,  �?���  �?���L  ����L  ����  �?���      E  , ,  �����  �����L  �����L  �����  �����      E  , ,  �w���  �w���L  �?���L  �?���  �w���      E  , ,  ����  ����L  �����L  �����  ����      E  , ,  �����  �����L  �w���L  �w���  �����      E  , ,  �K���  �K���L  ����L  ����  �K���      E  , ,  �����  �����L  �����L  �����  �����      E  , ,  �����  �����L  �K���L  �K���  �����      E  , ,  �k����  �k���  �3���  �3����  �k����      E  , ,  �����  ����  �����  ������  �����      E  , ,  ������  �����  �k���  �k����  ������      E  , ,  �?����  �?���  ����  �����  �?����      E  , ,  ������  �����  �����  ������  ������      E  , ,  �w����  �w���  �?���  �?����  �w����      E  , ,  �����  ����  �����  ������  �����      E  , ,  ������  �����  �w���  �w����  ������      E  , ,  �K����  �K���  ����  �����  �K����      E  , ,  ������  �����  �����  ������  ������      E  , ,  ������  �����  �K���  �K����  ������      E  , ,  �k���d  �k���,  �3���,  �3���d  �k���d      E  , ,  ����d  ����,  �����,  �����d  ����d      E  , ,  �����d  �����,  �k���,  �k���d  �����d      E  , ,  �?���d  �?���,  ����,  ����d  �?���d      E  , ,  �����d  �����,  �����,  �����d  �����d      E  , ,  �w���d  �w���,  �?���,  �?���d  �w���d      E  , ,  ����d  ����,  �����,  �����d  ����d      E  , ,  �����d  �����,  �w���,  �w���d  �����d      E  , ,  �K���d  �K���,  ����,  ����d  �K���d      E  , ,  �����d  �����,  �����,  �����d  �����d      E  , ,  �����d  �����,  �K���,  �K���d  �����d      E  , ,  �k����  �k���  �3���  �3����  �k����      E  , ,  �����  ����  �����  ������  �����      E  , ,  ������  �����  �k���  �k����  ������      E  , ,  �?����  �?���  ����  �����  �?����      E  , ,  ������  �����  �����  ������  ������      E  , ,  �w����  �w���  �?���  �?����  �w����      E  , ,  �����  ����  �����  ������  �����      E  , ,  ������  �����  �w���  �w����  ������      E  , ,  �K����  �K���  ����  �����  �K����      E  , ,  ������  �����  �����  ������  ������      E  , ,  ������  �����  �K���  �K����  ������      E  , ,  �k���D  �k���  �3���  �3���D  �k���D      E  , ,  ����D  ����  �����  �����D  ����D      E  , ,  �����D  �����  �k���  �k���D  �����D      E  , ,  �?���D  �?���  ����  ����D  �?���D      E  , ,  �����D  �����  �����  �����D  �����D      E  , ,  �w���D  �w���  �?���  �?���D  �w���D      E  , ,  ����D  ����  �����  �����D  ����D      E  , ,  �����D  �����  �w���  �w���D  �����D      E  , ,  �K���D  �K���  ����  ����D  �K���D      E  , ,  �����D  �����  �����  �����D  �����D      E  , ,  �����D  �����  �K���  �K���D  �����D      E  , ,  �k���P  �k���  �3���  �3���P  �k���P      E  , ,  ����P  ����  �����  �����P  ����P      E  , ,  �����P  �����  �k���  �k���P  �����P      E  , ,  �?���P  �?���  ����  ����P  �?���P      E  , ,  �����P  �����  �����  �����P  �����P      E  , ,  �w���P  �w���  �?���  �?���P  �w���P      E  , ,  ����P  ����  �����  �����P  ����P      E  , ,  �����P  �����  �w���  �w���P  �����P      E  , ,  �K���P  �K���  ����  ����P  �K���P      E  , ,  �����P  �����  �����  �����P  �����P      E  , ,  �����P  �����  �K���  �K���P  �����P      E  , ,  �k���  �k���l  �3���l  �3���  �k���      E  , ,  ����  ����l  �����l  �����  ����      E  , ,  �����  �����l  �k���l  �k���  �����      E  , ,  �?���  �?���l  ����l  ����  �?���      E  , ,  �����  �����l  �����l  �����  �����      E  , ,  �w���  �w���l  �?���l  �?���  �w���      E  , ,  ����  ����l  �����l  �����  ����      E  , ,  �����  �����l  �w���l  �w���  �����      E  , ,  �K���  �K���l  ����l  ����  �K���      E  , ,  �����  �����l  �����l  �����  �����      E  , ,  �����  �����l  �K���l  �K���  �����      E  , ,  `'���D  `'���  `����  `����D  `'���D      E  , ,  d����D  d����  e����  e����D  d����D      E  , ,  i_���D  i_���  j'���  j'���D  i_���D      E  , ,  m����D  m����  n����  n����D  m����D      E  , ,  r����D  r����  s_���  s_���D  r����D      E  , ,  w3���D  w3���  w����  w����D  w3���D      E  , ,  {����D  {����  |����  |����D  {����D      E  , ,  m����d  m����,  n����,  n����d  m����d      E  , ,  r����d  r����,  s_���,  s_���d  r����d      E  , ,  w3���d  w3���,  w����,  w����d  w3���d      E  , ,  {����d  {����,  |����,  |����d  {����d      E  , ,  w3���  w3���L  w����L  w����  w3���      E  , ,  `'����  `'���  `����  `�����  `'����      E  , ,  d�����  d����  e����  e�����  d�����      E  , ,  i_����  i_���  j'���  j'����  i_����      E  , ,  m�����  m����  n����  n�����  m�����      E  , ,  r�����  r����  s_���  s_����  r�����      E  , ,  w3����  w3���  w����  w�����  w3����      E  , ,  `'���P  `'���  `����  `����P  `'���P      E  , ,  d����P  d����  e����  e����P  d����P      E  , ,  i_���P  i_���  j'���  j'���P  i_���P      E  , ,  m����P  m����  n����  n����P  m����P      E  , ,  r����P  r����  s_���  s_���P  r����P      E  , ,  w3���P  w3���  w����  w����P  w3���P      E  , ,  {����P  {����  |����  |����P  {����P      E  , ,  {�����  {����  |����  |�����  {�����      E  , ,  {����  {����L  |����L  |����  {����      E  , ,  m����  m�����  n�����  n����  m����      E  , ,  r����  r�����  s_����  s_���  r����      E  , ,  `'����  `'���  `����  `�����  `'����      E  , ,  d�����  d����  e����  e�����  d�����      E  , ,  i_����  i_���  j'���  j'����  i_����      E  , ,  m�����  m����  n����  n�����  m�����      E  , ,  r�����  r����  s_���  s_����  r�����      E  , ,  w3����  w3���  w����  w�����  w3����      E  , ,  {�����  {����  |����  |�����  {�����      E  , ,  `'���  `'���l  `����l  `����  `'���      E  , ,  d����  d����l  e����l  e����  d����      E  , ,  i_���  i_���l  j'���l  j'���  i_���      E  , ,  m����  m����l  n����l  n����  m����      E  , ,  r����  r����l  s_���l  s_���  r����      E  , ,  w3���  w3���l  w����l  w����  w3���      E  , ,  {����  {����l  |����l  |����  {����      E  , ,  w3���  w3����  w�����  w����  w3���      E  , ,  {����  {�����  |�����  |����  {����      E  , ,  i_���  i_����  j'����  j'���  i_���      E  , ,  `'���  `'���L  `����L  `����  `'���      E  , ,  d����  d����L  e����L  e����  d����      E  , ,  i_���  i_���L  j'���L  j'���  i_���      E  , ,  m����  m����L  n����L  n����  m����      E  , ,  r����  r����L  s_���L  s_���  r����      E  , ,  `'���d  `'���,  `����,  `����d  `'���d      E  , ,  d����d  d����,  e����,  e����d  d����d      E  , ,  i_���d  i_���,  j'���,  j'���d  i_���d      E  , ,  `'���  `'����  `�����  `����  `'���      E  , ,  d����  d�����  e�����  e����  d����      E  , ,  {���ؠ  {����h  |����h  |���ؠ  {���ؠ      E  , ,  `'���  `'����  `�����  `����  `'���      E  , ,  d����  d�����  e�����  e����  d����      E  , ,  i_���  i_����  j'����  j'���  i_���      E  , ,  m����  m�����  n�����  n����  m����      E  , ,  r����  r�����  s_����  s_���  r����      E  , ,  w3���  w3����  w�����  w����  w3���      E  , ,  {����  {�����  |�����  |����  {����      E  , ,  `'��Հ  `'���H  `����H  `���Հ  `'��Հ      E  , ,  d���Հ  d����H  e����H  e���Հ  d���Հ      E  , ,  i_��Հ  i_���H  j'���H  j'��Հ  i_��Հ      E  , ,  m���Հ  m����H  n����H  n���Հ  m���Հ      E  , ,  r���Հ  r����H  s_���H  s_��Հ  r���Հ      E  , ,  w3��Հ  w3���H  w����H  w���Հ  w3��Հ      E  , ,  {���Հ  {����H  |����H  |���Հ  {���Հ      E  , ,  `'����  `'��Ը  `���Ը  `�����  `'����      E  , ,  d�����  d���Ը  e���Ը  e�����  d�����      E  , ,  i_����  i_��Ը  j'��Ը  j'����  i_����      E  , ,  m�����  m���Ը  n���Ը  n�����  m�����      E  , ,  r�����  r���Ը  s_��Ը  s_����  r�����      E  , ,  w3����  w3��Ը  w���Ը  w�����  w3����      E  , ,  {�����  {���Ը  |���Ը  |�����  {�����      E  , ,  `;��Ś  `;���b  a���b  a��Ś  `;��Ś      E  , ,  d���Ś  d����b  e����b  e���Ś  d���Ś      E  , ,  is��Ś  is���b  j;���b  j;��Ś  is��Ś      E  , ,  n��Ś  n���b  n����b  n���Ś  n��Ś      E  , ,  r���Ś  r����b  ss���b  ss��Ś  r���Ś      E  , ,  wG��Ś  wG���b  x���b  x��Ś  wG��Ś      E  , ,  {���Ś  {����b  |����b  |���Ś  {���Ś      E  , ,  `;���
  `;����  a����  a���
  `;���
      E  , ,  d����
  d�����  e�����  e����
  d����
      E  , ,  is���
  is����  j;����  j;���
  is���
      E  , ,  n���
  n����  n�����  n����
  n���
      E  , ,  r����
  r�����  ss����  ss���
  r����
      E  , ,  wG���
  wG����  x����  x���
  wG���
      E  , ,  {����
  {�����  |�����  |����
  {����
      E  , ,  `;���z  `;���B  a���B  a���z  `;���z      E  , ,  d����z  d����B  e����B  e����z  d����z      E  , ,  is���z  is���B  j;���B  j;���z  is���z      E  , ,  n���z  n���B  n����B  n����z  n���z      E  , ,  r����z  r����B  ss���B  ss���z  r����z      E  , ,  wG���z  wG���B  x���B  x���z  wG���z      E  , ,  {����z  {����B  |����B  |����z  {����z      E  , ,  `;����  `;����  a����  a����  `;����      E  , ,  d�����  d�����  e�����  e�����  d�����      E  , ,  is����  is����  j;����  j;����  is����      E  , ,  n����  n����  n�����  n�����  n����      E  , ,  r�����  r�����  ss����  ss����  r�����      E  , ,  wG����  wG����  x����  x����  wG����      E  , ,  {�����  {�����  |�����  |�����  {�����      E  , ,  `'����  `'��܈  `���܈  `�����  `'����      E  , ,  d�����  d���܈  e���܈  e�����  d�����      E  , ,  i_����  i_��܈  j'��܈  j'����  i_����      E  , ,  m�����  m���܈  n���܈  n�����  m�����      E  , ,  r�����  r���܈  s_��܈  s_����  r�����      E  , ,  w3����  w3��܈  w���܈  w�����  w3����      E  , ,  {�����  {���܈  |���܈  |�����  {�����      E  , ,  `'���0  `'����  `�����  `����0  `'���0      E  , ,  d����0  d�����  e�����  e����0  d����0      E  , ,  i_���0  i_����  j'����  j'���0  i_���0      E  , ,  m����0  m�����  n�����  n����0  m����0      E  , ,  r����0  r�����  s_����  s_���0  r����0      E  , ,  w3���0  w3����  w�����  w����0  w3���0      E  , ,  {����0  {�����  |�����  |����0  {����0      E  , ,  `'��ؠ  `'���h  `����h  `���ؠ  `'��ؠ      E  , ,  d���ؠ  d����h  e����h  e���ؠ  d���ؠ      E  , ,  i_��ؠ  i_���h  j'���h  j'��ؠ  i_��ؠ      E  , ,  m���ؠ  m����h  n����h  n���ؠ  m���ؠ      E  , ,  r���ؠ  r����h  s_���h  s_��ؠ  r���ؠ      E  , ,  w3��ؠ  w3���h  w����h  w���ؠ  w3��ؠ      E  , ,  �����0  ������  �K����  �K���0  �����0      E  , ,  ������  ����܈  �w��܈  �w����  ������      E  , ,  �K����  �K��܈  ���܈  �����  �K����      E  , ,  ������  ����܈  ����܈  ������  ������      E  , ,  ������  ����܈  �K��܈  �K����  ������      E  , ,  �����  ���Ը  ����Ը  ������  �����      E  , ,  ������  ����Ը  �w��Ը  �w����  ������      E  , ,  �K����  �K��Ը  ���Ը  �����  �K����      E  , ,  ������  ����Ը  ����Ը  ������  ������      E  , ,  ������  ����Ը  �K��Ը  �K����  ������      E  , ,  ���ؠ  ����h  �����h  ����ؠ  ���ؠ      E  , ,  ����ؠ  �����h  �w���h  �w��ؠ  ����ؠ      E  , ,  �K��ؠ  �K���h  ����h  ���ؠ  �K��ؠ      E  , ,  ����ؠ  �����h  �����h  ����ؠ  ����ؠ      E  , ,  ����ؠ  �����h  �K���h  �K��ؠ  ����ؠ      E  , ,  �����  ���܈  ����܈  ������  �����      E  , ,  ����  �����  ������  �����  ����      E  , ,  �����  ������  �w����  �w���  �����      E  , ,  �K���  �K����  �����  ����  �K���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �����  ������  �K����  �K���  �����      E  , ,  ����0  �����  ������  �����0  ����0      E  , ,  �����0  ������  �w����  �w���0  �����0      E  , ,  �K���0  �K����  �����  ����0  �K���0      E  , ,  �����0  ������  ������  �����0  �����0      E  , ,  ���Հ  ����H  �����H  ����Հ  ���Հ      E  , ,  ����Հ  �����H  �w���H  �w��Հ  ����Հ      E  , ,  �K��Հ  �K���H  ����H  ���Հ  �K��Հ      E  , ,  ����Հ  �����H  �����H  ����Հ  ����Հ      E  , ,  ����Հ  �����H  �K���H  �K��Հ  ����Հ      E  , ,  �?����  �?��܈  ���܈  �����  �?����      E  , ,  ������  ����܈  ����܈  ������  ������      E  , ,  �w����  �w��܈  �?��܈  �?����  �w����      E  , ,  �k����  �k��Ը  �3��Ը  �3����  �k����      E  , ,  �k���0  �k����  �3����  �3���0  �k���0      E  , ,  ����0  �����  ������  �����0  ����0      E  , ,  �����0  ������  �k����  �k���0  �����0      E  , ,  �k���  �k����  �3����  �3���  �k���      E  , ,  ����  �����  ������  �����  ����      E  , ,  �����  ������  �k����  �k���  �����      E  , ,  �?���  �?����  �����  ����  �?���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �w���  �w����  �?����  �?���  �w���      E  , ,  �����  ���Ը  ����Ը  ������  �����      E  , ,  ������  ����Ը  �k��Ը  �k����  ������      E  , ,  ������  ����܈  �k��܈  �k����  ������      E  , ,  �k��ؠ  �k���h  �3���h  �3��ؠ  �k��ؠ      E  , ,  ���ؠ  ����h  �����h  ����ؠ  ���ؠ      E  , ,  �?���0  �?����  �����  ����0  �?���0      E  , ,  �����0  ������  ������  �����0  �����0      E  , ,  �w���0  �w����  �?����  �?���0  �w���0      E  , ,  ����ؠ  �����h  �k���h  �k��ؠ  ����ؠ      E  , ,  �?��ؠ  �?���h  ����h  ���ؠ  �?��ؠ      E  , ,  ����ؠ  �����h  �����h  ����ؠ  ����ؠ      E  , ,  �w��ؠ  �w���h  �?���h  �?��ؠ  �w��ؠ      E  , ,  �k��Հ  �k���H  �3���H  �3��Հ  �k��Հ      E  , ,  ���Հ  ����H  �����H  ����Հ  ���Հ      E  , ,  ����Հ  �����H  �k���H  �k��Հ  ����Հ      E  , ,  �?��Հ  �?���H  ����H  ���Հ  �?��Հ      E  , ,  ����Հ  �����H  �����H  ����Հ  ����Հ      E  , ,  �w��Հ  �w���H  �?���H  �?��Հ  �w��Հ      E  , ,  �?����  �?��Ը  ���Ը  �����  �?����      E  , ,  ������  ����Ը  ����Ը  ������  ������      E  , ,  �w����  �w��Ը  �?��Ը  �?����  �w����      E  , ,  �k����  �k��܈  �3��܈  �3����  �k����      E  , ,  �����  ���܈  ����܈  ������  �����      E  , ,  ������  ������  �����  �����  ������      E  , ,  �S����  �S����  �����  �����  �S����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �S����  �S����  ������      E  , ,  �S��Ś  �S���b  ����b  ���Ś  �S��Ś      E  , ,  ����Ś  �����b  �����b  ����Ś  ����Ś      E  , ,  ����Ś  �����b  �S���b  �S��Ś  ����Ś      E  , ,  ���Ś  ����b  �G���b  �G��Ś  ���Ś      E  , ,  ����
  �����  �G����  �G���
  ����
      E  , ,  ����z  ����B  �G���B  �G���z  ����z      E  , ,  ����z  ����B  �����B  �����z  ����z      E  , ,  �����z  �����B  ����B  ����z  �����z      E  , ,  �S���z  �S���B  ����B  ����z  �S���z      E  , ,  �����z  �����B  �����B  �����z  �����z      E  , ,  �����z  �����B  �S���B  �S���z  �����z      E  , ,  ����
  �����  ������  �����
  ����
      E  , ,  �����
  ������  �����  ����
  �����
      E  , ,  �S���
  �S����  �����  ����
  �S���
      E  , ,  �����
  ������  ������  �����
  �����
      E  , ,  �����
  ������  �S����  �S���
  �����
      E  , ,  ���Ś  ����b  �����b  ����Ś  ���Ś      E  , ,  ����Ś  �����b  ����b  ���Ś  ����Ś      E  , ,  �����  �����  �G����  �G����  �����      E  , ,  �����  �����  ������  ������  �����      E  , ,  �����z  �����B  �����B  �����z  �����z      E  , ,  �����z  �����B  �_���B  �_���z  �����z      E  , ,  ����Ś  �����b  �����b  ����Ś  ����Ś      E  , ,  �_��Ś  �_���b  �'���b  �'��Ś  �_��Ś      E  , ,  �'���
  �'����  ������  �����
  �'���
      E  , ,  �����
  ������  ������  �����
  �����
      E  , ,  �_���
  �_����  �'����  �'���
  �_���
      E  , ,  �����
  ������  ������  �����
  �����
      E  , ,  �����
  ������  �_����  �_���
  �����
      E  , ,  ����Ś  �����b  �����b  ����Ś  ����Ś      E  , ,  ����Ś  �����b  �_���b  �_��Ś  ����Ś      E  , ,  �'��Ś  �'���b  �����b  ����Ś  �'��Ś      E  , ,  �'���z  �'���B  �����B  �����z  �'���z      E  , ,  �����z  �����B  �����B  �����z  �����z      E  , ,  �_���z  �_���B  �'���B  �'���z  �_���z      E  , ,  �'����  �'����  ������  ������  �'����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �_����  �_����  �'����  �'����  �_����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �_����  �_����  ������      E  , ,  �+����  �+���  �����  ������  �+����      E  , ,  ������  �����  Ϗ���  Ϗ����  ������      E  , ,  ŏ���  ŏ���L  �W���L  �W���  ŏ���      E  , ,  �+���  �+���L  �����L  �����  �+���      E  , ,  �����  �����L  Ϗ���L  Ϗ���  �����      E  , ,  �����  �����l  �����l  �����  �����      E  , ,  �W���  �W���l  ����l  ����  �W���      E  , ,  �����  �����l  �����l  �����  �����      E  , ,  ����  �����  ������  �����  ����      E  , ,  �����  ������  ������  �����  �����      E  , ,  �����  ����  �����  ������  �����      E  , ,  ����P  ����  �����  �����P  ����P      E  , ,  �����P  �����  �����  �����P  �����P      E  , ,  �W���P  �W���  ����  ����P  �W���P      E  , ,  �����P  �����  �����  �����P  �����P      E  , ,  ŏ���P  ŏ���  �W���  �W���P  ŏ���P      E  , ,  �+���P  �+���  �����  �����P  �+���P      E  , ,  �����P  �����  Ϗ���  Ϗ���P  �����P      E  , ,  ������  �����  �����  ������  ������      E  , ,  �W����  �W���  ����  �����  �W����      E  , ,  ������  �����  �����  ������  ������      E  , ,  ŏ����  ŏ���  �W���  �W����  ŏ����      E  , ,  �+����  �+���  �����  ������  �+����      E  , ,  ������  �����  Ϗ���  Ϗ����  ������      E  , ,  �W���  �W����  �����  ����  �W���      E  , ,  �����  ������  ������  �����  �����      E  , ,  ŏ���  ŏ����  �W����  �W���  ŏ���      E  , ,  �+���  �+����  ������  �����  �+���      E  , ,  �����  ������  Ϗ����  Ϗ���  �����      E  , ,  ŏ���  ŏ���l  �W���l  �W���  ŏ���      E  , ,  �+���  �+���l  �����l  �����  �+���      E  , ,  �����  �����l  Ϗ���l  Ϗ���  �����      E  , ,  ����  ����l  �����l  �����  ����      E  , ,  ����  ����L  �����L  �����  ����      E  , ,  ����d  ����,  �����,  �����d  ����d      E  , ,  �����d  �����,  �����,  �����d  �����d      E  , ,  �W���d  �W���,  ����,  ����d  �W���d      E  , ,  �����d  �����,  �����,  �����d  �����d      E  , ,  ŏ���d  ŏ���,  �W���,  �W���d  ŏ���d      E  , ,  �+���d  �+���,  �����,  �����d  �+���d      E  , ,  �����d  �����,  Ϗ���,  Ϗ���d  �����d      E  , ,  �����  �����L  �����L  �����  �����      E  , ,  ����D  ����  �����  �����D  ����D      E  , ,  �����D  �����  �����  �����D  �����D      E  , ,  �W���D  �W���  ����  ����D  �W���D      E  , ,  �����D  �����  �����  �����D  �����D      E  , ,  ŏ���D  ŏ���  �W���  �W���D  ŏ���D      E  , ,  �+���D  �+���  �����  �����D  �+���D      E  , ,  �����D  �����  Ϗ���  Ϗ���D  �����D      E  , ,  �W���  �W���L  ����L  ����  �W���      E  , ,  �����  �����L  �����L  �����  �����      E  , ,  �����  ����  �����  ������  �����      E  , ,  ������  �����  �����  ������  ������      E  , ,  �W����  �W���  ����  �����  �W����      E  , ,  ������  �����  �����  ������  ������      E  , ,  ŏ����  ŏ���  �W���  �W����  ŏ����      E  , ,  �?��Ś  �?���b  ����b  ���Ś  �?��Ś      E  , ,  ����Ś  �����b  ϣ���b  ϣ��Ś  ����Ś      E  , ,  �W��ؠ  �W���h  ����h  ���ؠ  �W��ؠ      E  , ,  ����ؠ  �����h  �����h  ����ؠ  ����ؠ      E  , ,  ŏ��ؠ  ŏ���h  �W���h  �W��ؠ  ŏ��ؠ      E  , ,  ����  �����  ������  �����  ����      E  , ,  �����  ������  ������  �����  �����      E  , ,  �W���  �W����  �����  ����  �W���      E  , ,  �����  ������  ������  �����  �����      E  , ,  ŏ���  ŏ����  �W����  �W���  ŏ���      E  , ,  �+���  �+����  ������  �����  �+���      E  , ,  �����  ������  Ϗ����  Ϗ���  �����      E  , ,  �+��ؠ  �+���h  �����h  ����ؠ  �+��ؠ      E  , ,  ����ؠ  �����h  Ϗ���h  Ϗ��ؠ  ����ؠ      E  , ,  �����  ���܈  ����܈  ������  �����      E  , ,  ������  ����܈  ����܈  ������  ������      E  , ,  �W����  �W��܈  ���܈  �����  �W����      E  , ,  ������  ����܈  ����܈  ������  ������      E  , ,  �3���z  �3���B  �����B  �����z  �3���z      E  , ,  �����z  �����B  �����B  �����z  �����z      E  , ,  �k���z  �k���B  �3���B  �3���z  �k���z      E  , ,  ����z  ����B  �����B  �����z  ����z      E  , ,  ţ���z  ţ���B  �k���B  �k���z  ţ���z      E  , ,  �?���z  �?���B  ����B  ����z  �?���z      E  , ,  �����z  �����B  ϣ���B  ϣ���z  �����z      E  , ,  ŏ����  ŏ��܈  �W��܈  �W����  ŏ����      E  , ,  �+����  �+��܈  ����܈  ������  �+����      E  , ,  ������  ����܈  Ϗ��܈  Ϗ����  ������      E  , ,  �+����  �+��Ը  ����Ը  ������  �+����      E  , ,  ������  ����Ը  Ϗ��Ը  Ϗ����  ������      E  , ,  ������  ����Ը  ����Ը  ������  ������      E  , ,  �W����  �W��Ը  ���Ը  �����  �W����      E  , ,  ������  ����Ը  ����Ը  ������  ������      E  , ,  ŏ����  ŏ��Ը  �W��Ը  �W����  ŏ����      E  , ,  ���ؠ  ����h  �����h  ����ؠ  ���ؠ      E  , ,  ����ؠ  �����h  �����h  ����ؠ  ����ؠ      E  , ,  �3��Ś  �3���b  �����b  ����Ś  �3��Ś      E  , ,  ���Հ  ����H  �����H  ����Հ  ���Հ      E  , ,  ����Հ  �����H  �����H  ����Հ  ����Հ      E  , ,  �W��Հ  �W���H  ����H  ���Հ  �W��Հ      E  , ,  ����Հ  �����H  �����H  ����Հ  ����Հ      E  , ,  ŏ��Հ  ŏ���H  �W���H  �W��Հ  ŏ��Հ      E  , ,  �+��Հ  �+���H  �����H  ����Հ  �+��Հ      E  , ,  �3����  �3����  ������  ������  �3����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �k����  �k����  �3����  �3����  �k����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ţ����  ţ����  �k����  �k����  ţ����      E  , ,  �?����  �?����  �����  �����  �?����      E  , ,  ������  ������  ϣ����  ϣ����  ������      E  , ,  ����Հ  �����H  Ϗ���H  Ϗ��Հ  ����Հ      E  , ,  ����Ś  �����b  �����b  ����Ś  ����Ś      E  , ,  �k��Ś  �k���b  �3���b  �3��Ś  �k��Ś      E  , ,  ���Ś  ����b  �����b  ����Ś  ���Ś      E  , ,  ţ��Ś  ţ���b  �k���b  �k��Ś  ţ��Ś      E  , ,  �3���
  �3����  ������  �����
  �3���
      E  , ,  �����
  ������  ������  �����
  �����
      E  , ,  �k���
  �k����  �3����  �3���
  �k���
      E  , ,  ����
  �����  ������  �����
  ����
      E  , ,  ţ���
  ţ����  �k����  �k���
  ţ���
      E  , ,  ����0  �����  ������  �����0  ����0      E  , ,  �����0  ������  ������  �����0  �����0      E  , ,  �W���0  �W����  �����  ����0  �W���0      E  , ,  �����0  ������  ������  �����0  �����0      E  , ,  ŏ���0  ŏ����  �W����  �W���0  ŏ���0      E  , ,  �+���0  �+����  ������  �����0  �+���0      E  , ,  �����0  ������  Ϗ����  Ϗ���0  �����0      E  , ,  �?���
  �?����  �����  ����
  �?���
      E  , ,  �����
  ������  ϣ����  ϣ���
  �����
      E  , ,  �����  ���Ը  ����Ը  ������  �����      E  , ,  �k���Z  �k���"  �3���"  �3���Z  �k���Z      E  , ,  ����Z  ����"  �����"  �����Z  ����Z      E  , ,  ţ���Z  ţ���"  �k���"  �k���Z  ţ���Z      E  , ,  �?���Z  �?���"  ����"  ����Z  �?���Z      E  , ,  �����Z  �����"  ϣ���"  ϣ���Z  �����Z      E  , ,  �3����  �3����  ������  ������  �3����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �k����  �k����  �3����  �3����  �k����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ţ����  ţ����  �k����  �k����  ţ����      E  , ,  �?����  �?����  �����  �����  �?����      E  , ,  ������  ������  ϣ����  ϣ����  ������      E  , ,  �3���:  �3���  �����  �����:  �3���:      E  , ,  �����:  �����  �����  �����:  �����:      E  , ,  �k���:  �k���  �3���  �3���:  �k���:      E  , ,  ����:  ����  �����  �����:  ����:      E  , ,  ţ���:  ţ���  �k���  �k���:  ţ���:      E  , ,  �?���:  �?���  ����  ����:  �?���:      E  , ,  �����:  �����  ϣ���  ϣ���:  �����:      E  , ,  �3���F  �3���  �����  �����F  �3���F      E  , ,  �����F  �����  �����  �����F  �����F      E  , ,  �k���F  �k���  �3���  �3���F  �k���F      E  , ,  ����F  ����  �����  �����F  ����F      E  , ,  ţ���F  ţ���  �k���  �k���F  ţ���F      E  , ,  �?���F  �?���  ����  ����F  �?���F      E  , ,  �����F  �����  ϣ���  ϣ���F  �����F      E  , ,  �3����  �3���~  �����~  ������  �3����      E  , ,  ������  �����~  �����~  ������  ������      E  , ,  �k����  �k���~  �3���~  �3����  �k����      E  , ,  �����  ����~  �����~  ������  �����      E  , ,  ţ����  ţ���~  �k���~  �k����  ţ����      E  , ,  �?����  �?���~  ����~  �����  �?����      E  , ,  ������  �����~  ϣ���~  ϣ����  ������      E  , ,  �3���&  �3����  ������  �����&  �3���&      E  , ,  �����&  ������  ������  �����&  �����&      E  , ,  �k���&  �k����  �3����  �3���&  �k���&      E  , ,  ����&  �����  ������  �����&  ����&      E  , ,  ţ���&  ţ����  �k����  �k���&  ţ���&      E  , ,  �?���&  �?����  �����  ����&  �?���&      E  , ,  �����&  ������  ϣ����  ϣ���&  �����&      E  , ,  �3����  �3���^  �����^  ������  �3����      E  , ,  ������  �����^  �����^  ������  ������      E  , ,  �k����  �k���^  �3���^  �3����  �k����      E  , ,  �����  ����^  �����^  ������  �����      E  , ,  ţ����  ţ���^  �k���^  �k����  ţ����      E  , ,  �?����  �?���^  ����^  �����  �?����      E  , ,  ������  �����^  ϣ���^  ϣ����  ������      E  , ,  �3���  �3����  ������  �����  �3���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �k���  �k����  �3����  �3���  �k���      E  , ,  ����  �����  ������  �����  ����      E  , ,  ţ���  ţ����  �k����  �k���  ţ���      E  , ,  �?���  �?����  �����  ����  �?���      E  , ,  �����  ������  ϣ����  ϣ���  �����      E  , ,  �3���v  �3���>  �����>  �����v  �3���v      E  , ,  �����v  �����>  �����>  �����v  �����v      E  , ,  �k���v  �k���>  �3���>  �3���v  �k���v      E  , ,  ����v  ����>  �����>  �����v  ����v      E  , ,  ţ���v  ţ���>  �k���>  �k���v  ţ���v      E  , ,  �?���v  �?���>  ����>  ����v  �?���v      E  , ,  �����v  �����>  ϣ���>  ϣ���v  �����v      E  , ,  �3����  �3����  ������  ������  �3����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �k����  �k����  �3����  �3����  �k����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ţ����  ţ����  �k����  �k����  ţ����      E  , ,  �?����  �?����  �����  �����  �?����      E  , ,  ������  ������  ϣ����  ϣ����  ������      E  , ,  �3���Z  �3���"  �����"  �����Z  �3���Z      E  , ,  �����Z  �����"  �����"  �����Z  �����Z      E  , ,  �k����  �k���X  �3���X  �3����  �k����      E  , ,  �����  ����X  �����X  ������  �����      E  , ,  ţ����  ţ���X  �k���X  �k����  ţ����      E  , ,  �?����  �?���X  ����X  �����  �?����      E  , ,  ������  �����X  ϣ���X  ϣ����  ������      E  , ,  �3���   �3����  ������  �����   �3���       E  , ,  �����   ������  ������  �����   �����       E  , ,  �k���   �k����  �3����  �3���   �k���       E  , ,  ����   �����  ������  �����   ����       E  , ,  ţ���   ţ����  �k����  �k���   ţ���       E  , ,  �?���   �?����  �����  ����   �?���       E  , ,  �����   ������  ϣ����  ϣ���   �����       E  , ,  �3���p  �3���8  �����8  �����p  �3���p      E  , ,  �����p  �����8  �����8  �����p  �����p      E  , ,  �k���p  �k���8  �3���8  �3���p  �k���p      E  , ,  ����p  ����8  �����8  �����p  ����p      E  , ,  ţ���p  ţ���8  �k���8  �k���p  ţ���p      E  , ,  �?���p  �?���8  ����8  ����p  �?���p      E  , ,  �����p  �����8  ϣ���8  ϣ���p  �����p      E  , ,  �3����  �3����  ������  ������  �3����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �k����  �k����  �3����  �3����  �k����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ţ����  ţ����  �k����  �k����  ţ����      E  , ,  �?����  �?����  �����  �����  �?����      E  , ,  ������  ������  ϣ����  ϣ����  ������      E  , ,  �3���P  �3���  �����  �����P  �3���P      E  , ,  �����P  �����  �����  �����P  �����P      E  , ,  �k���P  �k���  �3���  �3���P  �k���P      E  , ,  ����P  ����  �����  �����P  ����P      E  , ,  ţ���P  ţ���  �k���  �k���P  ţ���P      E  , ,  �?���P  �?���  ����  ����P  �?���P      E  , ,  �����P  �����  ϣ���  ϣ���P  �����P      E  , ,  �3����  �3����  ������  ������  �3����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �k����  �k����  �3����  �3����  �k����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ţ����  ţ����  �k����  �k����  ţ����      E  , ,  �?����  �?����  �����  �����  �?����      E  , ,  ������  ������  ϣ����  ϣ����  ������      E  , ,  �3���0  �3����  ������  �����0  �3���0      E  , ,  �����0  ������  ������  �����0  �����0      E  , ,  �k���0  �k����  �3����  �3���0  �k���0      E  , ,  ����0  �����  ������  �����0  ����0      E  , ,  ţ���0  ţ����  �k����  �k���0  ţ���0      E  , ,  �?���0  �?����  �����  ����0  �?���0      E  , ,  �����0  ������  ϣ����  ϣ���0  �����0      E  , ,  �3���<  �3���  �����  �����<  �3���<      E  , ,  �����<  �����  �����  �����<  �����<      E  , ,  �k���<  �k���  �3���  �3���<  �k���<      E  , ,  ����<  ����  �����  �����<  ����<      E  , ,  ţ���<  ţ���  �k���  �k���<  ţ���<      E  , ,  �?���<  �?���  ����  ����<  �?���<      E  , ,  �����<  �����  ϣ���  ϣ���<  �����<      E  , ,  �3����  �3���t  �����t  ������  �3����      E  , ,  ������  �����t  �����t  ������  ������      E  , ,  �k����  �k���t  �3���t  �3����  �k����      E  , ,  �����  ����t  �����t  ������  �����      E  , ,  ţ����  ţ���t  �k���t  �k����  ţ����      E  , ,  �?����  �?���t  ����t  �����  �?����      E  , ,  ������  �����t  ϣ���t  ϣ����  ������      E  , ,  �3���  �3����  ������  �����  �3���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �k���  �k����  �3����  �3���  �k���      E  , ,  ����  �����  ������  �����  ����      E  , ,  ţ���  ţ����  �k����  �k���  ţ���      E  , ,  �?���  �?����  �����  ����  �?���      E  , ,  �����  ������  ϣ����  ϣ���  �����      E  , ,  �3����  �3���T  �����T  ������  �3����      E  , ,  ������  �����T  �����T  ������  ������      E  , ,  �k����  �k���T  �3���T  �3����  �k����      E  , ,  �����  ����T  �����T  ������  �����      E  , ,  ţ����  ţ���T  �k���T  �k����  ţ����      E  , ,  �?����  �?���T  ����T  �����  �?����      E  , ,  ������  �����T  ϣ���T  ϣ����  ������      E  , ,  �3����  �3����  ������  ������  �3����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �k����  �k����  �3����  �3����  �k����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ţ����  ţ����  �k����  �k����  ţ����      E  , ,  �?����  �?����  �����  �����  �?����      E  , ,  ������  ������  ϣ����  ϣ����  ������      E  , ,  �3����  �3���X  �����X  ������  �3����      E  , ,  ������  �����X  �����X  ������  ������      E  , ,  �����:  �����  �����  �����:  �����:      E  , ,  �����:  �����  �_���  �_���:  �����:      E  , ,  �'����  �'����  ������  ������  �'����      E  , ,  �'���F  �'���  �����  �����F  �'���F      E  , ,  �����F  �����  �����  �����F  �����F      E  , ,  �_���F  �_���  �'���  �'���F  �_���F      E  , ,  �����F  �����  �����  �����F  �����F      E  , ,  �����F  �����  �_���  �_���F  �����F      E  , ,  ������  ������  ������  ������  ������      E  , ,  �_����  �_����  �'����  �'����  �_����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �_����  �_����  ������      E  , ,  �'����  �'���~  �����~  ������  �'����      E  , ,  ������  �����~  �����~  ������  ������      E  , ,  �_����  �_���~  �'���~  �'����  �_����      E  , ,  ������  �����~  �����~  ������  ������      E  , ,  ������  �����~  �_���~  �_����  ������      E  , ,  �'���&  �'����  ������  �����&  �'���&      E  , ,  �����&  ������  ������  �����&  �����&      E  , ,  �_���&  �_����  �'����  �'���&  �_���&      E  , ,  �����&  ������  ������  �����&  �����&      E  , ,  �����&  ������  �_����  �_���&  �����&      E  , ,  �'���:  �'���  �����  �����:  �'���:      E  , ,  �'���Z  �'���"  �����"  �����Z  �'���Z      E  , ,  �����Z  �����"  �����"  �����Z  �����Z      E  , ,  �_���Z  �_���"  �'���"  �'���Z  �_���Z      E  , ,  �����Z  �����"  �����"  �����Z  �����Z      E  , ,  �����Z  �����"  �_���"  �_���Z  �����Z      E  , ,  �����:  �����  �����  �����:  �����:      E  , ,  �_���:  �_���  �'���  �'���:  �_���:      E  , ,  �S���F  �S���  ����  ����F  �S���F      E  , ,  �����F  �����  �����  �����F  �����F      E  , ,  �����F  �����  �S���  �S���F  �����F      E  , ,  �����  �����  ������  ������  �����      E  , ,  ������  ������  �����  �����  ������      E  , ,  ����&  �����  �G����  �G���&  ����&      E  , ,  ����&  �����  ������  �����&  ����&      E  , ,  �����&  ������  �����  ����&  �����&      E  , ,  �S���&  �S����  �����  ����&  �S���&      E  , ,  �����&  ������  ������  �����&  �����&      E  , ,  �����&  ������  �S����  �S���&  �����&      E  , ,  �S����  �S����  �����  �����  �S����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �S����  �S����  ������      E  , ,  �����  �����  �G����  �G����  �����      E  , ,  ����F  ����  �G���  �G���F  ����F      E  , ,  ����:  ����  �G���  �G���:  ����:      E  , ,  ����:  ����  �����  �����:  ����:      E  , ,  �����:  �����  ����  ����:  �����:      E  , ,  �S���:  �S���  ����  ����:  �S���:      E  , ,  �����:  �����  �����  �����:  �����:      E  , ,  �����:  �����  �S���  �S���:  �����:      E  , ,  ����F  ����  �����  �����F  ����F      E  , ,  ����Z  ����"  �G���"  �G���Z  ����Z      E  , ,  ����Z  ����"  �����"  �����Z  ����Z      E  , ,  �����Z  �����"  ����"  ����Z  �����Z      E  , ,  �S���Z  �S���"  ����"  ����Z  �S���Z      E  , ,  �����Z  �����"  �����"  �����Z  �����Z      E  , ,  �����Z  �����"  �S���"  �S���Z  �����Z      E  , ,  �����F  �����  ����  ����F  �����F      E  , ,  �����  ����~  �G���~  �G����  �����      E  , ,  �����  ����~  �����~  ������  �����      E  , ,  ������  �����~  ����~  �����  ������      E  , ,  �S����  �S���~  ����~  �����  �S����      E  , ,  ������  �����~  �����~  ������  ������      E  , ,  ������  �����~  �S���~  �S����  ������      E  , ,  �����  ������  �S����  �S���  �����      E  , ,  �����  ����^  �G���^  �G����  �����      E  , ,  �����  ����^  �����^  ������  �����      E  , ,  ������  �����^  ����^  �����  ������      E  , ,  �S����  �S���^  ����^  �����  �S����      E  , ,  ������  �����^  �����^  ������  ������      E  , ,  ������  �����^  �S���^  �S����  ������      E  , ,  ����  �����  �G����  �G���  ����      E  , ,  ����v  ����>  �G���>  �G���v  ����v      E  , ,  ����v  ����>  �����>  �����v  ����v      E  , ,  �����v  �����>  ����>  ����v  �����v      E  , ,  �S���v  �S���>  ����>  ����v  �S���v      E  , ,  �����v  �����>  �����>  �����v  �����v      E  , ,  �����v  �����>  �S���>  �S���v  �����v      E  , ,  ����  �����  ������  �����  ����      E  , ,  �����  �����  �G����  �G����  �����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ������  ������  �����  �����  ������      E  , ,  �S����  �S����  �����  �����  �S����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �S����  �S����  ������      E  , ,  �����  ������  �����  ����  �����      E  , ,  �S���  �S����  �����  ����  �S���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �_����  �_���^  �'���^  �'����  �_����      E  , ,  ������  �����^  �����^  ������  ������      E  , ,  ������  �����^  �_���^  �_����  ������      E  , ,  �����v  �����>  �����>  �����v  �����v      E  , ,  �����v  �����>  �_���>  �_���v  �����v      E  , ,  �����  ������  ������  �����  �����      E  , ,  �����  ������  �_����  �_���  �����      E  , ,  �'���  �'����  ������  �����  �'���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �_���  �_����  �'����  �'���  �_���      E  , ,  �'���v  �'���>  �����>  �����v  �'���v      E  , ,  �����v  �����>  �����>  �����v  �����v      E  , ,  �'����  �'����  ������  ������  �'����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �_����  �_����  �'����  �'����  �_����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �_����  �_����  ������      E  , ,  �_���v  �_���>  �'���>  �'���v  �_���v      E  , ,  �'����  �'���^  �����^  ������  �'����      E  , ,  ������  �����^  �����^  ������  ������      E  , ,  `;���:  `;���  a���  a���:  `;���:      E  , ,  d����:  d����  e����  e����:  d����:      E  , ,  is���:  is���  j;���  j;���:  is���:      E  , ,  `;���&  `;����  a����  a���&  `;���&      E  , ,  d����&  d�����  e�����  e����&  d����&      E  , ,  is���&  is����  j;����  j;���&  is���&      E  , ,  n���&  n����  n�����  n����&  n���&      E  , ,  r����&  r�����  ss����  ss���&  r����&      E  , ,  wG���&  wG����  x����  x���&  wG���&      E  , ,  {����&  {�����  |�����  |����&  {����&      E  , ,  d����v  d����>  e����>  e����v  d����v      E  , ,  {����F  {����  |����  |����F  {����F      E  , ,  is���v  is���>  j;���>  j;���v  is���v      E  , ,  n���v  n���>  n����>  n����v  n���v      E  , ,  r����v  r����>  ss���>  ss���v  r����v      E  , ,  `;���F  `;���  a���  a���F  `;���F      E  , ,  d����F  d����  e����  e����F  d����F      E  , ,  is���F  is���  j;���  j;���F  is���F      E  , ,  n���F  n���  n����  n����F  n���F      E  , ,  r����F  r����  ss���  ss���F  r����F      E  , ,  wG���F  wG���  x���  x���F  wG���F      E  , ,  n���:  n���  n����  n����:  n���:      E  , ,  r����:  r����  ss���  ss���:  r����:      E  , ,  wG���:  wG���  x���  x���:  wG���:      E  , ,  {����:  {����  |����  |����:  {����:      E  , ,  `;����  `;����  a����  a����  `;����      E  , ,  d�����  d�����  e�����  e�����  d�����      E  , ,  is����  is����  j;����  j;����  is����      E  , ,  `;����  `;���^  a���^  a����  `;����      E  , ,  d�����  d����^  e����^  e�����  d�����      E  , ,  is����  is���^  j;���^  j;����  is����      E  , ,  n����  n���^  n����^  n�����  n����      E  , ,  r�����  r����^  ss���^  ss����  r�����      E  , ,  wG����  wG���^  x���^  x����  wG����      E  , ,  {�����  {����^  |����^  |�����  {�����      E  , ,  n����  n����  n�����  n�����  n����      E  , ,  r�����  r�����  ss����  ss����  r�����      E  , ,  wG����  wG����  x����  x����  wG����      E  , ,  `;����  `;����  a����  a����  `;����      E  , ,  d�����  d�����  e�����  e�����  d�����      E  , ,  is����  is����  j;����  j;����  is����      E  , ,  `;����  `;���~  a���~  a����  `;����      E  , ,  d�����  d����~  e����~  e�����  d�����      E  , ,  is����  is���~  j;���~  j;����  is����      E  , ,  n����  n���~  n����~  n�����  n����      E  , ,  r�����  r����~  ss���~  ss����  r�����      E  , ,  wG����  wG���~  x���~  x����  wG����      E  , ,  {�����  {����~  |����~  |�����  {�����      E  , ,  {�����  {�����  |�����  |�����  {�����      E  , ,  wG���v  wG���>  x���>  x���v  wG���v      E  , ,  `;���Z  `;���"  a���"  a���Z  `;���Z      E  , ,  d����Z  d����"  e����"  e����Z  d����Z      E  , ,  is���Z  is���"  j;���"  j;���Z  is���Z      E  , ,  n���Z  n���"  n����"  n����Z  n���Z      E  , ,  r����Z  r����"  ss���"  ss���Z  r����Z      E  , ,  wG���Z  wG���"  x���"  x���Z  wG���Z      E  , ,  {����Z  {����"  |����"  |����Z  {����Z      E  , ,  {����v  {����>  |����>  |����v  {����v      E  , ,  r����  r�����  ss����  ss���  r����      E  , ,  wG���  wG����  x����  x���  wG���      E  , ,  {����  {�����  |�����  |����  {����      E  , ,  `;���  `;����  a����  a���  `;���      E  , ,  d����  d�����  e�����  e����  d����      E  , ,  is���  is����  j;����  j;���  is���      E  , ,  n���  n����  n�����  n����  n���      E  , ,  `;���v  `;���>  a���>  a���v  `;���v      E  , ,  n����  n����  n�����  n�����  n����      E  , ,  r�����  r�����  ss����  ss����  r�����      E  , ,  wG����  wG����  x����  x����  wG����      E  , ,  {�����  {�����  |�����  |�����  {�����      E  , ,  {����<  {����  |����  |����<  {����<      E  , ,  `;����  `;���X  a���X  a����  `;����      E  , ,  d�����  d����X  e����X  e�����  d�����      E  , ,  is����  is���X  j;���X  j;����  is����      E  , ,  n����  n���X  n����X  n�����  n����      E  , ,  r�����  r����X  ss���X  ss����  r�����      E  , ,  wG����  wG���X  x���X  x����  wG����      E  , ,  {�����  {����X  |����X  |�����  {�����      E  , ,  `;����  `;���t  a���t  a����  `;����      E  , ,  d�����  d����t  e����t  e�����  d�����      E  , ,  is����  is���t  j;���t  j;����  is����      E  , ,  n����  n���t  n����t  n�����  n����      E  , ,  r�����  r����t  ss���t  ss����  r�����      E  , ,  wG����  wG���t  x���t  x����  wG����      E  , ,  {�����  {����t  |����t  |�����  {�����      E  , ,  `;���P  `;���  a���  a���P  `;���P      E  , ,  d����P  d����  e����  e����P  d����P      E  , ,  is���P  is���  j;���  j;���P  is���P      E  , ,  n���P  n���  n����  n����P  n���P      E  , ,  r����P  r����  ss���  ss���P  r����P      E  , ,  wG���P  wG���  x���  x���P  wG���P      E  , ,  {����P  {����  |����  |����P  {����P      E  , ,  `;���  `;����  a����  a���  `;���      E  , ,  d����  d�����  e�����  e����  d����      E  , ,  is���  is����  j;����  j;���  is���      E  , ,  n���  n����  n�����  n����  n���      E  , ,  r����  r�����  ss����  ss���  r����      E  , ,  wG���  wG����  x����  x���  wG���      E  , ,  {����  {�����  |�����  |����  {����      E  , ,  `;���p  `;���8  a���8  a���p  `;���p      E  , ,  d����p  d����8  e����8  e����p  d����p      E  , ,  is���p  is���8  j;���8  j;���p  is���p      E  , ,  n���p  n���8  n����8  n����p  n���p      E  , ,  r����p  r����8  ss���8  ss���p  r����p      E  , ,  wG���p  wG���8  x���8  x���p  wG���p      E  , ,  {����p  {����8  |����8  |����p  {����p      E  , ,  `;����  `;���T  a���T  a����  `;����      E  , ,  d�����  d����T  e����T  e�����  d�����      E  , ,  is����  is���T  j;���T  j;����  is����      E  , ,  n����  n���T  n����T  n�����  n����      E  , ,  r�����  r����T  ss���T  ss����  r�����      E  , ,  wG����  wG���T  x���T  x����  wG����      E  , ,  {�����  {����T  |����T  |�����  {�����      E  , ,  `;����  `;����  a����  a����  `;����      E  , ,  d�����  d�����  e�����  e�����  d�����      E  , ,  is����  is����  j;����  j;����  is����      E  , ,  n����  n����  n�����  n�����  n����      E  , ,  r�����  r�����  ss����  ss����  r�����      E  , ,  wG����  wG����  x����  x����  wG����      E  , ,  {�����  {�����  |�����  |�����  {�����      E  , ,  `;����  `;����  a����  a����  `;����      E  , ,  d�����  d�����  e�����  e�����  d�����      E  , ,  is����  is����  j;����  j;����  is����      E  , ,  n����  n����  n�����  n�����  n����      E  , ,  r�����  r�����  ss����  ss����  r�����      E  , ,  wG����  wG����  x����  x����  wG����      E  , ,  {�����  {�����  |�����  |�����  {�����      E  , ,  `;���   `;����  a����  a���   `;���       E  , ,  d����   d�����  e�����  e����   d����       E  , ,  is���   is����  j;����  j;���   is���       E  , ,  n���   n����  n�����  n����   n���       E  , ,  r����   r�����  ss����  ss���   r����       E  , ,  wG���   wG����  x����  x���   wG���       E  , ,  {����   {�����  |�����  |����   {����       E  , ,  `;���0  `;����  a����  a���0  `;���0      E  , ,  d����0  d�����  e�����  e����0  d����0      E  , ,  is���0  is����  j;����  j;���0  is���0      E  , ,  n���0  n����  n�����  n����0  n���0      E  , ,  r����0  r�����  ss����  ss���0  r����0      E  , ,  wG���0  wG����  x����  x���0  wG���0      E  , ,  {����0  {�����  |�����  |����0  {����0      E  , ,  `;����  `;����  a����  a����  `;����      E  , ,  d�����  d�����  e�����  e�����  d�����      E  , ,  is����  is����  j;����  j;����  is����      E  , ,  n����  n����  n�����  n�����  n����      E  , ,  r�����  r�����  ss����  ss����  r�����      E  , ,  wG����  wG����  x����  x����  wG����      E  , ,  {�����  {�����  |�����  |�����  {�����      E  , ,  `;���<  `;���  a���  a���<  `;���<      E  , ,  d����<  d����  e����  e����<  d����<      E  , ,  is���<  is���  j;���  j;���<  is���<      E  , ,  n���<  n���  n����  n����<  n���<      E  , ,  r����<  r����  ss���  ss���<  r����<      E  , ,  wG���<  wG���  x���  x���<  wG���<      E  , ,  �'���P  �'���  �����  �����P  �'���P      E  , ,  �����P  �����  �����  �����P  �����P      E  , ,  �_���P  �_���  �'���  �'���P  �_���P      E  , ,  �����P  �����  �����  �����P  �����P      E  , ,  �����P  �����  �_���  �_���P  �����P      E  , ,  �'���p  �'���8  �����8  �����p  �'���p      E  , ,  �����p  �����8  �����8  �����p  �����p      E  , ,  �_���p  �_���8  �'���8  �'���p  �_���p      E  , ,  �����p  �����8  �����8  �����p  �����p      E  , ,  �����p  �����8  �_���8  �_���p  �����p      E  , ,  �'���   �'����  ������  �����   �'���       E  , ,  �����   ������  ������  �����   �����       E  , ,  �_���   �_����  �'����  �'���   �_���       E  , ,  �����   ������  ������  �����   �����       E  , ,  �����   ������  �_����  �_���   �����       E  , ,  �'����  �'����  ������  ������  �'����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �_����  �_����  �'����  �'����  �_����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �_����  �_����  ������      E  , ,  �'����  �'���X  �����X  ������  �'����      E  , ,  ������  �����X  �����X  ������  ������      E  , ,  �_����  �_���X  �'���X  �'����  �_����      E  , ,  �'����  �'����  ������  ������  �'����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �_����  �_����  �'����  �'����  �_����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �_����  �_����  ������      E  , ,  ������  �����X  �����X  ������  ������      E  , ,  ������  �����X  �_���X  �_����  ������      E  , ,  �S����  �S����  �����  �����  �S����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �S����  �S����  ������      E  , ,  �����P  �����  �S���  �S���P  �����P      E  , ,  �����p  �����8  �����8  �����p  �����p      E  , ,  �����p  �����8  �S���8  �S���p  �����p      E  , ,  �S���   �S����  �����  ����   �S���       E  , ,  �����   ������  ������  �����   �����       E  , ,  ������  �����X  �����X  ������  ������      E  , ,  ������  �����X  �S���X  �S����  ������      E  , ,  �����   ������  �S����  �S���   �����       E  , ,  ����P  ����  �G���  �G���P  ����P      E  , ,  ����P  ����  �����  �����P  ����P      E  , ,  �����  �����  �G����  �G����  �����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ������  ������  �����  �����  ������      E  , ,  �S����  �S����  �����  �����  �S����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �S����  �S����  ������      E  , ,  �����P  �����  ����  ����P  �����P      E  , ,  �S���P  �S���  ����  ����P  �S���P      E  , ,  �����P  �����  �����  �����P  �����P      E  , ,  �S����  �S���X  ����X  �����  �S����      E  , ,  �����  �����  �G����  �G����  �����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ������  ������  �����  �����  ������      E  , ,  �����  ����X  �G���X  �G����  �����      E  , ,  �����  ����X  �����X  ������  �����      E  , ,  ������  �����X  ����X  �����  ������      E  , ,  ����   �����  �G����  �G���   ����       E  , ,  ����   �����  ������  �����   ����       E  , ,  �����   ������  �����  ����   �����       E  , ,  ����p  ����8  �G���8  �G���p  ����p      E  , ,  ����p  ����8  �����8  �����p  ����p      E  , ,  �����p  �����8  ����8  ����p  �����p      E  , ,  �S���p  �S���8  ����8  ����p  �S���p      E  , ,  �����  ������  �����  ����  �����      E  , ,  �S���  �S����  �����  ����  �S���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �����  ������  �S����  �S���  �����      E  , ,  ����0  �����  �G����  �G���0  ����0      E  , ,  ����0  �����  ������  �����0  ����0      E  , ,  �����0  ������  �����  ����0  �����0      E  , ,  �S���0  �S����  �����  ����0  �S���0      E  , ,  �����  �����  �G����  �G����  �����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ������  ������  �����  �����  ������      E  , ,  �S����  �S����  �����  �����  �S����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �S����  �S����  ������      E  , ,  �����0  ������  ������  �����0  �����0      E  , ,  �����0  ������  �S����  �S���0  �����0      E  , ,  ������  �����t  ����t  �����  ������      E  , ,  �S����  �S���t  ����t  �����  �S����      E  , ,  �����  ����T  �G���T  �G����  �����      E  , ,  �����  ����T  �����T  ������  �����      E  , ,  ������  �����T  ����T  �����  ������      E  , ,  �S����  �S���T  ����T  �����  �S����      E  , ,  ������  �����T  �����T  ������  ������      E  , ,  ������  �����T  �S���T  �S����  ������      E  , ,  ������  �����t  �����t  ������  ������      E  , ,  ������  �����t  �S���t  �S����  ������      E  , ,  �����  ����t  �G���t  �G����  �����      E  , ,  �����  ����t  �����t  ������  �����      E  , ,  ����  �����  �G����  �G���  ����      E  , ,  ����  �����  ������  �����  ����      E  , ,  ����<  ����  �G���  �G���<  ����<      E  , ,  ����<  ����  �����  �����<  ����<      E  , ,  �����<  �����  ����  ����<  �����<      E  , ,  �S���<  �S���  ����  ����<  �S���<      E  , ,  �����<  �����  �����  �����<  �����<      E  , ,  �����<  �����  �S���  �S���<  �����<      E  , ,  �_����  �_����  �'����  �'����  �_����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �_����  �_����  ������      E  , ,  �'����  �'���t  �����t  ������  �'����      E  , ,  ������  �����t  �����t  ������  ������      E  , ,  �'���0  �'����  ������  �����0  �'���0      E  , ,  �����0  ������  ������  �����0  �����0      E  , ,  �_���0  �_����  �'����  �'���0  �_���0      E  , ,  �����0  ������  ������  �����0  �����0      E  , ,  �����0  ������  �_����  �_���0  �����0      E  , ,  �_����  �_���t  �'���t  �'����  �_����      E  , ,  ������  �����t  �����t  ������  ������      E  , ,  ������  �����t  �_���t  �_����  ������      E  , ,  �'���  �'����  ������  �����  �'���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �_���  �_����  �'����  �'���  �_���      E  , ,  �����  ������  ������  �����  �����      E  , ,  �����  ������  �_����  �_���  �����      E  , ,  �'���<  �'���  �����  �����<  �'���<      E  , ,  �����<  �����  �����  �����<  �����<      E  , ,  �_���<  �_���  �'���  �'���<  �_���<      E  , ,  �����<  �����  �����  �����<  �����<      E  , ,  �����<  �����  �_���  �_���<  �����<      E  , ,  �'����  �'���T  �����T  ������  �'����      E  , ,  ������  �����T  �����T  ������  ������      E  , ,  �_����  �_���T  �'���T  �'����  �_����      E  , ,  ������  �����T  �����T  ������  ������      E  , ,  ������  �����T  �_���T  �_����  ������      E  , ,  �'����  �'����  ������  ������  �'����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �����  �����  �G����  �G����  �����      E  , ,  �����  �����  ������  ������  �����      E  , ,  ������  ������  �����  �����  ������      E  , ,  �S����  �S����  �����  �����  �S����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �S����  �S����  ������      E  , ,  �'����  �'����  ������  ������  �'����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �_����  �_����  �'����  �'����  �_����      E  , ,  ������  ������  ������  ������  ������      E  , ,  ������  ������  �_����  �_����  ������      E  , ,  ����q�  ����r�  ����r�  ����q�  ����q�      E  , ,  �s��q�  �s��r�  �;��r�  �;��q�  �s��q�      E  , ,  ���q�  ���r�  ����r�  ����q�  ���q�      E  , ,  ����q�  ����r�  �s��r�  �s��q�  ����q�      E  , ,  �G��q�  �G��r�  ���r�  ���q�  �G��q�      E  , ,  �	��q�  �	��r�  ����r�  ����q�  �	��q�      E  , ,  ����q�  ����r�  �m��r�  �m��q�  ����q�      E  , ,  �A��q�  �A��r�  �	��r�  �	��q�  �A��q�      E  , ,  ����q�  ����r�  ����r�  ����q�  ����q�      E  , ,  �y��q�  �y��r�  �A��r�  �A��q�  �y��q�      E  , ,  ����p1  ����p�  ����p�  ����p1  ����p1      E  , ,  �s��p1  �s��p�  �;��p�  �;��p1  �s��p1      E  , ,  ���p1  ���p�  ����p�  ����p1  ���p1      E  , ,  ����p1  ����p�  �s��p�  �s��p1  ����p1      E  , ,  �G��p1  �G��p�  ���p�  ���p1  �G��p1      E  , ,  �	��p1  �	��p�  ����p�  ����p1  �	��p1      E  , ,  ����p1  ����p�  �m��p�  �m��p1  ����p1      E  , ,  �A��p1  �A��p�  �	��p�  �	��p1  �A��p1      E  , ,  ����p1  ����p�  ����p�  ����p1  ����p1      E  , ,  �y��p1  �y��p�  �A��p�  �A��p1  �y��p1      E  , ,  ����n�  ����oi  ����oi  ����n�  ����n�      E  , ,  �s��n�  �s��oi  �;��oi  �;��n�  �s��n�      E  , ,  ���n�  ���oi  ����oi  ����n�  ���n�      E  , ,  ����n�  ����oi  �s��oi  �s��n�  ����n�      E  , ,  �G��n�  �G��oi  ���oi  ���n�  �G��n�      E  , ,  �	��n�  �	��oi  ����oi  ����n�  �	��n�      E  , ,  ����n�  ����oi  �m��oi  �m��n�  ����n�      E  , ,  �A��n�  �A��oi  �	��oi  �	��n�  �A��n�      E  , ,  ����n�  ����oi  ����oi  ����n�  ����n�      E  , ,  �y��n�  �y��oi  �A��oi  �A��n�  �y��n�      E  , ,  ����m  ����m�  ����m�  ����m  ����m      E  , ,  �s��m  �s��m�  �;��m�  �;��m  �s��m      E  , ,  ���m  ���m�  ����m�  ����m  ���m      E  , ,  ����m  ����m�  �s��m�  �s��m  ����m      E  , ,  �G��m  �G��m�  ���m�  ���m  �G��m      E  , ,  �	��m  �	��m�  ����m�  ����m  �	��m      E  , ,  ����m  ����m�  �m��m�  �m��m  ����m      E  , ,  �A��m  �A��m�  �	��m�  �	��m  �A��m      E  , ,  ����m  ����m�  ����m�  ����m  ����m      E  , ,  �y��m  �y��m�  �A��m�  �A��m  �y��m      E  , ,  ����k�  ����lI  ����lI  ����k�  ����k�      E  , ,  �s��k�  �s��lI  �;��lI  �;��k�  �s��k�      E  , ,  ���k�  ���lI  ����lI  ����k�  ���k�      E  , ,  ����k�  ����lI  �s��lI  �s��k�  ����k�      E  , ,  �G��k�  �G��lI  ���lI  ���k�  �G��k�      E  , ,  �	��k�  �	��lI  ����lI  ����k�  �	��k�      E  , ,  ����k�  ����lI  �m��lI  �m��k�  ����k�      E  , ,  �A��k�  �A��lI  �	��lI  �	��k�  �A��k�      E  , ,  ����k�  ����lI  ����lI  ����k�  ����k�      E  , ,  �y��k�  �y��lI  �A��lI  �A��k�  �y��k�      E  , ,  ����i�  ����j�  ����j�  ����i�  ����i�      E  , ,  �s��i�  �s��j�  �;��j�  �;��i�  �s��i�      E  , ,  ���i�  ���j�  ����j�  ����i�  ���i�      E  , ,  ����i�  ����j�  �s��j�  �s��i�  ����i�      E  , ,  �G��i�  �G��j�  ���j�  ���i�  �G��i�      E  , ,  �	��i�  �	��j�  ����j�  ����i�  �	��i�      E  , ,  ����i�  ����j�  �m��j�  �m��i�  ����i�      E  , ,  �A��i�  �A��j�  �	��j�  �	��i�  �A��i�      E  , ,  ����i�  ����j�  ����j�  ����i�  ����i�      E  , ,  �y��i�  �y��j�  �A��j�  �A��i�  �y��i�      E  , ,  ����l  ����4  �G���4  �G���l  ����l      E  , ,  ����l  ����4  �����4  �����l  ����l      E  , ,  �����l  �����4  ����4  ����l  �����l      E  , ,  �S���l  �S���4  ����4  ����l  �S���l      E  , ,  �����l  �����4  �����4  �����l  �����l      E  , ,  �����l  �����4  �S���4  �S���l  �����l      E  , ,  �'���l  �'���4  �����4  �����l  �'���l      E  , ,  �����l  �����4  �����4  �����l  �����l      E  , ,  �_���l  �_���4  �'���4  �'���l  �_���l      E  , ,  �����l  �����4  �����4  �����l  �����l      E  , ,  �����l  �����4  �_���4  �_���l  �����l      E  , ,  u��n�  u��oi  u���oi  u���n�  u��n�      E  , ,  y���n�  y���oi  zg��oi  zg��n�  y���n�      E  , ,  ~;��n�  ~;��oi  ��oi  ��n�  ~;��n�      E  , ,  N���xe  N���y-  Ot��y-  Ot��xe  N���xe      E  , ,  N���v�  N���w�  Ot��w�  Ot��v�  N���v�      E  , ,  N���uE  N���v  Ot��v  Ot��uE  N���uE      E  , ,  N���s�  N���t}  Ot��t}  Ot��s�  N���s�      E  , ,  `;���l  `;���4  a���4  a���l  `;���l      E  , ,  N���p�  N���q]  Ot��q]  Ot��p�  N���p�      E  , ,  u��p1  u��p�  u���p�  u���p1  u��p1      E  , ,  r����l  r����4  ss���4  ss���l  r����l      E  , ,  u��i�  u��j�  u���j�  u���i�  u��i�      E  , ,  y���i�  y���j�  zg��j�  zg��i�  y���i�      E  , ,  ~;��i�  ~;��j�  ��j�  ��i�  ~;��i�      E  , ,  y���p1  y���p�  zg��p�  zg��p1  y���p1      E  , ,  ~;��p1  ~;��p�  ��p�  ��p1  ~;��p1      E  , ,  N���r%  N���r�  Ot��r�  Ot��r%  N���r%      E  , ,  is���l  is���4  j;���4  j;���l  is���l      E  , ,  u��m  u��m�  u���m�  u���m  u��m      E  , ,  y���m  y���m�  zg��m�  zg��m  y���m      E  , ,  ~;��m  ~;��m�  ��m�  ��m  ~;��m      E  , ,  u��q�  u��r�  u���r�  u���q�  u��q�      E  , ,  y���q�  y���r�  zg��r�  zg��q�  y���q�      E  , ,  ~;��q�  ~;��r�  ��r�  ��q�  ~;��q�      E  , ,  wG���l  wG���4  x���4  x���l  wG���l      E  , ,  {����l  {����4  |����4  |����l  {����l      E  , ,  n����  n����  n�����  n�����  n����      E  , ,  r�����  r�����  ss����  ss����  r�����      E  , ,  wG����  wG����  x����  x����  wG����      E  , ,  {�����  {�����  |�����  |�����  {�����      E  , ,  is����  is����  j;����  j;����  is����      E  , ,  N���y�  N���z�  Ot��z�  Ot��y�  N���y�      E  , ,  d����l  d����4  e����4  e����l  d����l      E  , ,  n���l  n���4  n����4  n����l  n���l      E  , ,  u��k�  u��lI  u���lI  u���k�  u��k�      E  , ,  y���k�  y���lI  zg��lI  zg��k�  y���k�      E  , ,  ~;��k�  ~;��lI  ��lI  ��k�  ~;��k�      E  , ,  `;����  `;����  a����  a����  `;����      E  , ,  d�����  d�����  e�����  e�����  d�����      E  , ,  y���^�  y���_o  zg��_o  zg��^�  y���^�      E  , ,  ~;��^�  ~;��_o  ��_o  ��^�  ~;��^�      E  , ,  u��]  u��]�  u���]�  u���]  u��]      E  , ,  y���]  y���]�  zg��]�  zg��]  y���]      E  , ,  ~;��]  ~;��]�  ��]�  ��]  ~;��]      E  , ,  u��[�  u��\O  u���\O  u���[�  u��[�      E  , ,  y���[�  y���\O  zg��\O  zg��[�  y���[�      E  , ,  ~;��[�  ~;��\O  ��\O  ��[�  ~;��[�      E  , ,  y���ha  y���i)  zg��i)  zg��ha  y���ha      E  , ,  u��Y�  u��Z�  u���Z�  u���Y�  u��Y�      E  , ,  y���Y�  y���Z�  zg��Z�  zg��Y�  y���Y�      E  , ,  ~;��Y�  ~;��Z�  ��Z�  ��Y�  ~;��Y�      E  , ,  ~;��ha  ~;��i)  ��i)  ��ha  ~;��ha      E  , ,  u��Xg  u��Y/  u���Y/  u���Xg  u��Xg      E  , ,  y���Xg  y���Y/  zg��Y/  zg��Xg  y���Xg      E  , ,  ~;��Xg  ~;��Y/  ��Y/  ��Xg  ~;��Xg      E  , ,  u��ha  u��i)  u���i)  u���ha  u��ha      E  , ,  u��a�  u��b�  u���b�  u���a�  u��a�      E  , ,  y���a�  y���b�  zg��b�  zg��a�  y���a�      E  , ,  ~;��a�  ~;��b�  ��b�  ��a�  ~;��a�      E  , ,  u��`7  u��`�  u���`�  u���`7  u��`7      E  , ,  y���`7  y���`�  zg��`�  zg��`7  y���`7      E  , ,  ~;��`7  ~;��`�  ��`�  ��`7  ~;��`7      E  , ,  u��^�  u��_o  u���_o  u���^�  u��^�      E  , ,  �	��`7  �	��`�  ����`�  ����`7  �	��`7      E  , ,  ����`7  ����`�  �m��`�  �m��`7  ����`7      E  , ,  �A��`7  �A��`�  �	��`�  �	��`7  �A��`7      E  , ,  ����`7  ����`�  ����`�  ����`7  ����`7      E  , ,  �y��`7  �y��`�  �A��`�  �A��`7  �y��`7      E  , ,  ����ha  ����i)  ����i)  ����ha  ����ha      E  , ,  �s��ha  �s��i)  �;��i)  �;��ha  �s��ha      E  , ,  ���ha  ���i)  ����i)  ����ha  ���ha      E  , ,  ����^�  ����_o  ����_o  ����^�  ����^�      E  , ,  �s��^�  �s��_o  �;��_o  �;��^�  �s��^�      E  , ,  ���^�  ���_o  ����_o  ����^�  ���^�      E  , ,  ����^�  ����_o  �s��_o  �s��^�  ����^�      E  , ,  �G��^�  �G��_o  ���_o  ���^�  �G��^�      E  , ,  �	��^�  �	��_o  ����_o  ����^�  �	��^�      E  , ,  ����^�  ����_o  �m��_o  �m��^�  ����^�      E  , ,  �A��^�  �A��_o  �	��_o  �	��^�  �A��^�      E  , ,  ����^�  ����_o  ����_o  ����^�  ����^�      E  , ,  �y��^�  �y��_o  �A��_o  �A��^�  �y��^�      E  , ,  ����ha  ����i)  �s��i)  �s��ha  ����ha      E  , ,  �G��ha  �G��i)  ���i)  ���ha  �G��ha      E  , ,  �	��ha  �	��i)  ����i)  ����ha  �	��ha      E  , ,  ����]  ����]�  ����]�  ����]  ����]      E  , ,  �s��]  �s��]�  �;��]�  �;��]  �s��]      E  , ,  ���]  ���]�  ����]�  ����]  ���]      E  , ,  ����]  ����]�  �s��]�  �s��]  ����]      E  , ,  �G��]  �G��]�  ���]�  ���]  �G��]      E  , ,  �	��]  �	��]�  ����]�  ����]  �	��]      E  , ,  ����]  ����]�  �m��]�  �m��]  ����]      E  , ,  �A��]  �A��]�  �	��]�  �	��]  �A��]      E  , ,  ����]  ����]�  ����]�  ����]  ����]      E  , ,  �y��]  �y��]�  �A��]�  �A��]  �y��]      E  , ,  ����ha  ����i)  �m��i)  �m��ha  ����ha      E  , ,  ����a�  ����b�  ����b�  ����a�  ����a�      E  , ,  �s��a�  �s��b�  �;��b�  �;��a�  �s��a�      E  , ,  ����[�  ����\O  ����\O  ����[�  ����[�      E  , ,  �s��[�  �s��\O  �;��\O  �;��[�  �s��[�      E  , ,  ���[�  ���\O  ����\O  ����[�  ���[�      E  , ,  ����[�  ����\O  �s��\O  �s��[�  ����[�      E  , ,  �G��[�  �G��\O  ���\O  ���[�  �G��[�      E  , ,  �	��[�  �	��\O  ����\O  ����[�  �	��[�      E  , ,  ����[�  ����\O  �m��\O  �m��[�  ����[�      E  , ,  �A��[�  �A��\O  �	��\O  �	��[�  �A��[�      E  , ,  ����[�  ����\O  ����\O  ����[�  ����[�      E  , ,  �y��[�  �y��\O  �A��\O  �A��[�  �y��[�      E  , ,  ���a�  ���b�  ����b�  ����a�  ���a�      E  , ,  ����a�  ����b�  �s��b�  �s��a�  ����a�      E  , ,  �G��a�  �G��b�  ���b�  ���a�  �G��a�      E  , ,  �	��a�  �	��b�  ����b�  ����a�  �	��a�      E  , ,  ����Y�  ����Z�  ����Z�  ����Y�  ����Y�      E  , ,  �s��Y�  �s��Z�  �;��Z�  �;��Y�  �s��Y�      E  , ,  ���Y�  ���Z�  ����Z�  ����Y�  ���Y�      E  , ,  ����Y�  ����Z�  �s��Z�  �s��Y�  ����Y�      E  , ,  �G��Y�  �G��Z�  ���Z�  ���Y�  �G��Y�      E  , ,  �	��Y�  �	��Z�  ����Z�  ����Y�  �	��Y�      E  , ,  ����Y�  ����Z�  �m��Z�  �m��Y�  ����Y�      E  , ,  �A��Y�  �A��Z�  �	��Z�  �	��Y�  �A��Y�      E  , ,  ����Y�  ����Z�  ����Z�  ����Y�  ����Y�      E  , ,  �y��Y�  �y��Z�  �A��Z�  �A��Y�  �y��Y�      E  , ,  ����a�  ����b�  �m��b�  �m��a�  ����a�      E  , ,  �A��a�  �A��b�  �	��b�  �	��a�  �A��a�      E  , ,  ����a�  ����b�  ����b�  ����a�  ����a�      E  , ,  �y��a�  �y��b�  �A��b�  �A��a�  �y��a�      E  , ,  ����Xg  ����Y/  ����Y/  ����Xg  ����Xg      E  , ,  �s��Xg  �s��Y/  �;��Y/  �;��Xg  �s��Xg      E  , ,  ���Xg  ���Y/  ����Y/  ����Xg  ���Xg      E  , ,  ����Xg  ����Y/  �s��Y/  �s��Xg  ����Xg      E  , ,  �G��Xg  �G��Y/  ���Y/  ���Xg  �G��Xg      E  , ,  �	��Xg  �	��Y/  ����Y/  ����Xg  �	��Xg      E  , ,  ����Xg  ����Y/  �m��Y/  �m��Xg  ����Xg      E  , ,  �A��Xg  �A��Y/  �	��Y/  �	��Xg  �A��Xg      E  , ,  ����Xg  ����Y/  ����Y/  ����Xg  ����Xg      E  , ,  �y��Xg  �y��Y/  �A��Y/  �A��Xg  �y��Xg      E  , ,  �A��ha  �A��i)  �	��i)  �	��ha  �A��ha      E  , ,  ����ha  ����i)  ����i)  ����ha  ����ha      E  , ,  �y��ha  �y��i)  �A��i)  �A��ha  �y��ha      E  , ,  ����`7  ����`�  ����`�  ����`7  ����`7      E  , ,  �s��`7  �s��`�  �;��`�  �;��`7  �s��`7      E  , ,  ���`7  ���`�  ����`�  ����`7  ���`7      E  , ,  ����`7  ����`�  �s��`�  �s��`7  ����`7      E  , ,  �G��`7  �G��`�  ���`�  ���`7  �G��`7      E  , ,  ����i�  ����ji  ����ji  ����i�  ����i�      E  , ,  ����i�  ����ji  �k��ji  �k��i�  ����i�      E  , ,  ����i�  ����ji  �O��ji  �O��i�  ����i�      E  , ,  �k��i�  �k��ji  �3��ji  �3��i�  �k��i�      E  , ,  O��i�  O��ji ��ji ��i�  O��i�      E  , , 3��i� 3��ji ���ji ���i� 3��i�      E  , , ��i� ��ji ���ji ���i� ��i�      E  , , ���i� ���ji 	���ji 	���i� ���i�      E  , , ���i� ���ji ���ji ���i� ���i�      E  , , ���i� ���ji ���ji ���i� ���i�      E  , , ���i� ���ji o��ji o��i� ���i�      E  , ,  ����o�  ����p�  ����p�  ����o�  ����o�      E  , ,  ����o�  ����p�  �k��p�  �k��o�  ����o�      E  , ,  ����o�  ����p�  �O��p�  �O��o�  ����o�      E  , ,  �k��o�  �k��p�  �3��p�  �3��o�  �k��o�      E  , ,  O��o�  O��p� ��p� ��o�  O��o�      E  , , 3��o� 3��p� ���p� ���o� 3��o�      E  , , ��o� ��p� ���p� ���o� ��o�      E  , , ���o� ���p� 	���p� 	���o� ���o�      E  , , ���o� ���p� ���p� ���o� ���o�      E  , , ���o� ���p� ���p� ���o� ���o�      E  , , ���o� ���p� o��p� o��o� ���o�      E  , ,  ����k1  ����k�  ����k�  ����k1  ����k1      E  , ,  ����k1  ����k�  �k��k�  �k��k1  ����k1      E  , ,  ����k1  ����k�  �O��k�  �O��k1  ����k1      E  , ,  �k��k1  �k��k�  �3��k�  �3��k1  �k��k1      E  , ,  O��k1  O��k� ��k� ��k1  O��k1      E  , , 3��k1 3��k� ���k� ���k1 3��k1      E  , , ��k1 ��k� ���k� ���k1 ��k1      E  , , ���k1 ���k� 	���k� 	���k1 ���k1      E  , , ���k1 ���k� ���k� ���k1 ���k1      E  , , ���k1 ���k� ���k� ���k1 ���k1      E  , , ���k1 ���k� o��k� o��k1 ���k1      E  , ,  ����qq  ����r9  ����r9  ����qq  ����qq      E  , ,  ����qq  ����r9  �k��r9  �k��qq  ����qq      E  , ,  ����qq  ����r9  �O��r9  �O��qq  ����qq      E  , ,  �k��qq  �k��r9  �3��r9  �3��qq  �k��qq      E  , ,  O��qq  O��r9 ��r9 ��qq  O��qq      E  , , 3��qq 3��r9 ���r9 ���qq 3��qq      E  , , ��qq ��r9 ���r9 ���qq ��qq      E  , , ���qq ���r9 	���r9 	���qq ���qq      E  , , ���qq ���r9 ���r9 ���qq ���qq      E  , , ���qq ���r9 ���r9 ���qq ���qq      E  , , ���qq ���r9 o��r9 o��qq ���qq      E  , ,  ����l�  ����m�  ����m�  ����l�  ����l�      E  , ,  ����l�  ����m�  �k��m�  �k��l�  ����l�      E  , ,  ����l�  ����m�  �O��m�  �O��l�  ����l�      E  , ,  �k��l�  �k��m�  �3��m�  �3��l�  �k��l�      E  , ,  O��l�  O��m� ��m� ��l�  O��l�      E  , , 3��l� 3��m� ���m� ���l� 3��l�      E  , , ��l� ��m� ���m� ���l� ��l�      E  , , ���l� ���m� 	���m� 	���l� ���l�      E  , , ���l� ���m� ���m� ���l� ���l�      E  , , ���l� ���m� ���m� ���l� ���l�      E  , , ���l� ���m� o��m� o��l� ���l�      E  , ,  ����nQ  ����o  ����o  ����nQ  ����nQ      E  , ,  ����nQ  ����o  �k��o  �k��nQ  ����nQ      E  , ,  ����nQ  ����o  �O��o  �O��nQ  ����nQ      E  , ,  �k��nQ  �k��o  �3��o  �3��nQ  �k��nQ      E  , ,  O��nQ  O��o ��o ��nQ  O��nQ      E  , , 3��nQ 3��o ���o ���nQ 3��nQ      E  , , ��nQ ��o ���o ���nQ ��nQ      E  , , ���nQ ���o 	���o 	���nQ ���nQ      E  , , ���nQ ���o ���o ���nQ ���nQ      E  , , ���nQ ���o ���o ���nQ ���nQ      E  , , ���nQ ���o o��o o��nQ ���nQ      E  , ,  �����  �����  ������  ������  �����      E  , ,  ���k�  ���lI  ����lI  ����k�  ���k�      E  , ,  ����k�  ����lI  �y��lI  �y��k�  ����k�      E  , ,  �k���l  �k���4  �3���4  �3���l  �k���l      E  , ,  ���i�  ���j�  ����j�  ����i�  ���i�      E  , ,  ����i�  ����j�  �y��j�  �y��i�  ����i�      E  , ,  �M��i�  �M��j�  ���j�  ���i�  �M��i�      E  , ,  �M��k�  �M��lI  ���lI  ���k�  �M��k�      E  , ,  ţ����  ţ����  �k����  �k����  ţ����      E  , ,  �?����  �?����  �����  �����  �?����      E  , ,  ������  ������  ϣ����  ϣ����  ������      E  , ,  ţ���l  ţ���4  �k���4  �k���l  ţ���l      E  , ,  �?���l  �?���4  ����4  ����l  �?���l      E  , ,  �����l  �����4  ϣ���4  ϣ���l  �����l      E  , ,  ���p1  ���p�  ����p�  ����p1  ���p1      E  , ,  ����p1  ����p�  �y��p�  �y��p1  ����p1      E  , ,  �M��p1  �M��p�  ���p�  ���p1  �M��p1      E  , ,  �3���l  �3���4  �����4  �����l  �3���l      E  , ,  ���n�  ���oi  ����oi  ����n�  ���n�      E  , ,  ����n�  ����oi  �y��oi  �y��n�  ����n�      E  , ,  �M��n�  �M��oi  ���oi  ���n�  �M��n�      E  , ,  �����l  �����4  �����4  �����l  �����l      E  , ,  ����q�  ����r�  �y��r�  �y��q�  ����q�      E  , ,  �M��q�  �M��r�  ���r�  ���q�  �M��q�      E  , ,  ���q�  ���r�  ����r�  ����q�  ���q�      E  , ,  ���m  ���m�  ����m�  ����m  ���m      E  , ,  ����m  ����m�  �y��m�  �y��m  ����m      E  , ,  �M��m  �M��m�  ���m�  ���m  �M��m      E  , ,  ����l  ����4  �����4  �����l  ����l      E  , ,  �3����  �3����  ������  ������  �3����      E  , ,  ������  ������  ������  ������  ������      E  , ,  �k����  �k����  �3����  �3����  �k����      E  , ,  ���Y�  ���Z�  ����Z�  ����Y�  ���Y�      E  , ,  ����Y�  ����Z�  �y��Z�  �y��Y�  ����Y�      E  , ,  �M��Y�  �M��Z�  ���Z�  ���Y�  �M��Y�      E  , ,  �M��[�  �M��\O  ���\O  ���[�  �M��[�      E  , ,  ����a�  ����b�  �y��b�  �y��a�  ����a�      E  , ,  ���^�  ���_o  ����_o  ����^�  ���^�      E  , ,  ����^�  ����_o  �y��_o  �y��^�  ����^�      E  , ,  �M��^�  �M��_o  ���_o  ���^�  �M��^�      E  , ,  �M��a�  �M��b�  ���b�  ���a�  �M��a�      E  , ,  ���a�  ���b�  ����b�  ����a�  ���a�      E  , ,  ���`7  ���`�  ����`�  ����`7  ���`7      E  , ,  ����`7  ����`�  �y��`�  �y��`7  ����`7      E  , ,  ���]  ���]�  ����]�  ����]  ���]      E  , ,  ����]  ����]�  �y��]�  �y��]  ����]      E  , ,  �M��]  �M��]�  ���]�  ���]  �M��]      E  , ,  �M��`7  �M��`�  ���`�  ���`7  �M��`7      E  , ,  ���[�  ���\O  ����\O  ����[�  ���[�      E  , ,  ���Xg  ���Y/  ����Y/  ����Xg  ���Xg      E  , ,  ����Xg  ����Y/  �y��Y/  �y��Xg  ����Xg      E  , ,  �M��Xg  �M��Y/  ���Y/  ���Xg  �M��Xg      E  , ,  ����[�  ����\O  �y��\O  �y��[�  ����[�      E  , ,  ���ha  ���i)  ����i)  ����ha  ���ha      E  , ,  ����ha  ����i)  �y��i)  �y��ha  ����ha      E  , ,  �M��ha  �M��i)  ���i)  ���ha  �M��ha      E  , ,  ����[  ����[�  ����[�  ����[  ����[      E  , ,  ����[  ����[�  �k��[�  �k��[  ����[      E  , ,  ����[  ����[�  �O��[�  �O��[  ����[      E  , ,  �k��[  �k��[�  �3��[�  �3��[  �k��[      E  , ,  O��[  O��[� ��[� ��[  O��[      E  , , 3��[ 3��[� ���[� ���[ 3��[      E  , , ��[ ��[� ���[� ���[ ��[      E  , , ���[ ���[� 	���[� 	���[ ���[      E  , , ���[ ���[� ���[� ���[ ���[      E  , , ���[ ���[� ���[� ���[ ���[      E  , , ���[ ���[� o��[� o��[ ���[      E  , , ���h ���h� 	���h� 	���h ���h      E  , , ���ca ���d) o��d) o��ca ���ca      E  , , ���h ���h� ���h� ���h ���h      E  , , ���h ���h� ���h� ���h ���h      E  , , ���h ���h� o��h� o��h ���h      E  , ,  O��h  O��h� ��h� ��h  O��h      E  , ,  �k��f�  �k��gI  �3��gI  �3��f�  �k��f�      E  , ,  O��f�  O��gI ��gI ��f�  O��f�      E  , , 3��f� 3��gI ���gI ���f� 3��f�      E  , , ��f� ��gI ���gI ���f� ��f�      E  , , ���f� ���gI 	���gI 	���f� ���f�      E  , , ���f� ���gI ���gI ���f� ���f�      E  , , ���f� ���gI ���gI ���f� ���f�      E  , , ���f� ���gI o��gI o��f� ���f�      E  , , 3��h 3��h� ���h� ���h 3��h      E  , ,  �k��d�  �k��e�  �3��e�  �3��d�  �k��d�      E  , ,  O��d�  O��e� ��e� ��d�  O��d�      E  , , 3��d� 3��e� ���e� ���d� 3��d�      E  , , ��d� ��e� ���e� ���d� ��d�      E  , , ���d� ���e� 	���e� 	���d� ���d�      E  , , ���d� ���e� ���e� ���d� ���d�      E  , , ���d� ���e� ���e� ���d� ���d�      E  , , ���d� ���e� o��e� o��d� ���d�      E  , , ��h ��h� ���h� ���h ��h      E  , ,  �k��ca  �k��d)  �3��d)  �3��ca  �k��ca      E  , ,  O��ca  O��d) ��d) ��ca  O��ca      E  , , 3��ca 3��d) ���d) ���ca 3��ca      E  , , ��ca ��d) ���d) ���ca ��ca      E  , , ���ca ���d) 	���d) 	���ca ���ca      E  , , ���ca ���d) ���d) ���ca ���ca      E  , , ���ca ���d) ���d) ���ca ���ca      E  , ,  �k��h  �k��h�  �3��h�  �3��h  �k��h      E  , ,  ����ca  ����d)  �O��d)  �O��ca  ����ca      E  , ,  ����d�  ����e�  ����e�  ����d�  ����d�      E  , ,  ����d�  ����e�  �k��e�  �k��d�  ����d�      E  , ,  ����d�  ����e�  �O��e�  �O��d�  ����d�      E  , ,  ����f�  ����gI  ����gI  ����f�  ����f�      E  , ,  ����f�  ����gI  �k��gI  �k��f�  ����f�      E  , ,  ����f�  ����gI  �O��gI  �O��f�  ����f�      E  , ,  ����ca  ����d)  ����d)  ����ca  ����ca      E  , ,  ����h  ����h�  ����h�  ����h  ����h      E  , ,  ����h  ����h�  �k��h�  �k��h  ����h      E  , ,  ����h  ����h�  �O��h�  �O��h  ����h      E  , ,  ����ca  ����d)  �k��d)  �k��ca  ����ca      E  , ,  ����V_  ����W'  �k��W'  �k��V_  ����V_      E  , ,  ����V_  ����W'  �O��W'  �O��V_  ����V_      E  , ,  ����Y  ����ZG  ����ZG  ����Y  ����Y      E  , ,  ����T�  ����U�  ����U�  ����T�  ����T�      E  , ,  ����T�  ����U�  �k��U�  �k��T�  ����T�      E  , ,  ����T�  ����U�  �O��U�  �O��T�  ����T�      E  , ,  ����Y  ����ZG  �k��ZG  �k��Y  ����Y      E  , ,  ����S?  ����T  ����T  ����S?  ����S?      E  , ,  ����S?  ����T  �k��T  �k��S?  ����S?      E  , ,  ����S?  ����T  �O��T  �O��S?  ����S?      E  , ,  ����W�  ����X�  ����X�  ����W�  ����W�      E  , ,  ����Q�  ����Rw  ����Rw  ����Q�  ����Q�      E  , ,  ����Q�  ����Rw  �k��Rw  �k��Q�  ����Q�      E  , ,  ����Q�  ����Rw  �O��Rw  �O��Q�  ����Q�      E  , ,  ����W�  ����X�  �k��X�  �k��W�  ����W�      E  , ,  ����P  ����P�  ����P�  ����P  ����P      E  , ,  ����P  ����P�  �k��P�  �k��P  ����P      E  , ,  ����P  ����P�  �O��P�  �O��P  ����P      E  , ,  ����W�  ����X�  �O��X�  �O��W�  ����W�      E  , ,  ����N�  ����OW  ����OW  ����N�  ����N�      E  , ,  ����N�  ����OW  �k��OW  �k��N�  ����N�      E  , ,  ����N�  ����OW  �O��OW  �O��N�  ����N�      E  , ,  ����Y  ����ZG  �O��ZG  �O��Y  ����Y      E  , ,  ����L�  ����M�  ����M�  ����L�  ����L�      E  , ,  ����L�  ����M�  �k��M�  �k��L�  ����L�      E  , ,  ����L�  ����M�  �O��M�  �O��L�  ����L�      E  , ,  ����V_  ����W'  ����W'  ����V_  ����V_      E  , ,  O��Y  O��ZG ��ZG ��Y  O��Y      E  , , 3��Y 3��ZG ���ZG ���Y 3��Y      E  , , ��Y ��ZG ���ZG ���Y ��Y      E  , ,  �k��T�  �k��U�  �3��U�  �3��T�  �k��T�      E  , ,  O��T�  O��U� ��U� ��T�  O��T�      E  , , 3��T� 3��U� ���U� ���T� 3��T�      E  , , ��T� ��U� ���U� ���T� ��T�      E  , , ���T� ���U� 	���U� 	���T� ���T�      E  , , ���T� ���U� ���U� ���T� ���T�      E  , , ���T� ���U� ���U� ���T� ���T�      E  , , ���T� ���U� o��U� o��T� ���T�      E  , ,  �k��W�  �k��X�  �3��X�  �3��W�  �k��W�      E  , ,  O��W�  O��X� ��X� ��W�  O��W�      E  , , 3��W� 3��X� ���X� ���W� 3��W�      E  , , ��W� ��X� ���X� ���W� ��W�      E  , ,  �k��S?  �k��T  �3��T  �3��S?  �k��S?      E  , ,  O��S?  O��T ��T ��S?  O��S?      E  , , 3��S? 3��T ���T ���S? 3��S?      E  , , ��S? ��T ���T ���S? ��S?      E  , , ���S? ���T 	���T 	���S? ���S?      E  , , ���S? ���T ���T ���S? ���S?      E  , , ���S? ���T ���T ���S? ���S?      E  , , ���S? ���T o��T o��S? ���S?      E  , , ���W� ���X� 	���X� 	���W� ���W�      E  , , ���W� ���X� ���X� ���W� ���W�      E  , , ���W� ���X� ���X� ���W� ���W�      E  , , ���W� ���X� o��X� o��W� ���W�      E  , ,  �k��Q�  �k��Rw  �3��Rw  �3��Q�  �k��Q�      E  , ,  O��Q�  O��Rw ��Rw ��Q�  O��Q�      E  , , 3��Q� 3��Rw ���Rw ���Q� 3��Q�      E  , , ��Q� ��Rw ���Rw ���Q� ��Q�      E  , , ���Q� ���Rw 	���Rw 	���Q� ���Q�      E  , , ���Q� ���Rw ���Rw ���Q� ���Q�      E  , , ���Q� ���Rw ���Rw ���Q� ���Q�      E  , , ���Q� ���Rw o��Rw o��Q� ���Q�      E  , , ���Y ���ZG 	���ZG 	���Y ���Y      E  , , ���Y ���ZG ���ZG ���Y ���Y      E  , , ���Y ���ZG ���ZG ���Y ���Y      E  , , ���Y ���ZG o��ZG o��Y ���Y      E  , ,  �k��P  �k��P�  �3��P�  �3��P  �k��P      E  , ,  O��P  O��P� ��P� ��P  O��P      E  , , 3��P 3��P� ���P� ���P 3��P      E  , , ��P ��P� ���P� ���P ��P      E  , , ���P ���P� 	���P� 	���P ���P      E  , , ���P ���P� ���P� ���P ���P      E  , , ���P ���P� ���P� ���P ���P      E  , , ���P ���P� o��P� o��P ���P      E  , ,  �k��V_  �k��W'  �3��W'  �3��V_  �k��V_      E  , ,  O��V_  O��W' ��W' ��V_  O��V_      E  , , 3��V_ 3��W' ���W' ���V_ 3��V_      E  , , ��V_ ��W' ���W' ���V_ ��V_      E  , ,  �k��N�  �k��OW  �3��OW  �3��N�  �k��N�      E  , ,  O��N�  O��OW ��OW ��N�  O��N�      E  , , 3��N� 3��OW ���OW ���N� 3��N�      E  , , ��N� ��OW ���OW ���N� ��N�      E  , , ���N� ���OW 	���OW 	���N� ���N�      E  , , ���N� ���OW ���OW ���N� ���N�      E  , , ���N� ���OW ���OW ���N� ���N�      E  , , ���N� ���OW o��OW o��N� ���N�      E  , , ���V_ ���W' 	���W' 	���V_ ���V_      E  , , ���V_ ���W' ���W' ���V_ ���V_      E  , , ���V_ ���W' ���W' ���V_ ���V_      E  , , ���V_ ���W' o��W' o��V_ ���V_      E  , ,  �k��L�  �k��M�  �3��M�  �3��L�  �k��L�      E  , ,  O��L�  O��M� ��M� ��L�  O��L�      E  , , 3��L� 3��M� ���M� ���L� 3��L�      E  , , ��L� ��M� ���M� ���L� ��L�      E  , , ���L� ���M� 	���M� 	���L� ���L�      E  , , ���L� ���M� ���M� ���L� ���L�      E  , , ���L� ���M� ���M� ���L� ���L�      E  , , ���L� ���M� o��M� o��L� ���L�      E  , ,  �k��Y  �k��ZG  �3��ZG  �3��Y  �k��Y      E  , , o��i� o��ji 7��ji 7��i� o��i�      E  , , S��i� S��ji ��ji ��i� S��i�      E  , , 7��i� 7��ji ���ji ���i� 7��i�      E  , ,  ��i�  ��ji  ���ji  ���i�  ��i�      E  , , "���i� "���ji #���ji #���i� "���i�      E  , , %���i� %���ji &���ji &���i� %���i�      E  , , (���i� (���ji )���ji )���i� (���i�      E  , , +���i� +���ji ,s��ji ,s��i� +���i�      E  , , .���i� .���ji /W��ji /W��i� .���i�      E  , , 1s��i� 1s��ji 2;��ji 2;��i� 1s��i�      E  , , 4W��i� 4W��ji 5��ji 5��i� 4W��i�      E  , , 7;��i� 7;��ji 8��ji 8��i� 7;��i�      E  , , :��i� :��ji :���ji :���i� :��i�      E  , , =��i� =��ji =���ji =���i� =��i�      E  , , ?���i� ?���ji @���ji @���i� ?���i�      E  , , B���i� B���ji C���ji C���i� B���i�      E  , , E���i� E���ji Fw��ji Fw��i� E���i�      E  , , H���i� H���ji I[��ji I[��i� H���i�      E  , , Kw��i� Kw��ji L?��ji L?��i� Kw��i�      E  , , N[��i� N[��ji O#��ji O#��i� N[��i�      E  , , Q?��i� Q?��ji R��ji R��i� Q?��i�      E  , , T#��i� T#��ji T���ji T���i� T#��i�      E  , , W��i� W��ji W���ji W���i� W��i�      E  , , Y���i� Y���ji Z���ji Z���i� Y���i�      E  , , \���i� \���ji ]���ji ]���i� \���i�      E  , , _���i� _���ji `{��ji `{��i� _���i�      E  , , b���i� b���ji c_��ji c_��i� b���i�      E  , , e{��i� e{��ji fC��ji fC��i� e{��i�      E  , , h_��i� h_��ji i'��ji i'��i� h_��i�      E  , , kC��i� kC��ji l��ji l��i� kC��i�      E  , , n'��i� n'��ji n���ji n���i� n'��i�      E  , , q��i� q��ji q���ji q���i� q��i�      E  , , s���i� s���ji t���ji t���i� s���i�      E  , , v���i� v���ji w���ji w���i� v���i�      E  , , h_��o� h_��p� i'��p� i'��o� h_��o�      E  , , kC��o� kC��p� l��p� l��o� kC��o�      E  , , n'��o� n'��p� n���p� n���o� n'��o�      E  , , q��o� q��p� q���p� q���o� q��o�      E  , , s���o� s���p� t���p� t���o� s���o�      E  , , v���o� v���p� w���p� w���o� v���o�      E  , , \���o� \���p� ]���p� ]���o� \���o�      E  , , _���o� _���p� `{��p� `{��o� _���o�      E  , , b���o� b���p� c_��p� c_��o� b���o�      E  , , e{��o� e{��p� fC��p� fC��o� e{��o�      E  , , kC��qq kC��r9 l��r9 l��qq kC��qq      E  , , n'��qq n'��r9 n���r9 n���qq n'��qq      E  , , q��qq q��r9 q���r9 q���qq q��qq      E  , , s���qq s���r9 t���r9 t���qq s���qq      E  , , v���qq v���r9 w���r9 w���qq v���qq      E  , , H���nQ H���o I[��o I[��nQ H���nQ      E  , , Kw��nQ Kw��o L?��o L?��nQ Kw��nQ      E  , , N[��nQ N[��o O#��o O#��nQ N[��nQ      E  , , Q?��nQ Q?��o R��o R��nQ Q?��nQ      E  , , T#��nQ T#��o T���o T���nQ T#��nQ      E  , , W��nQ W��o W���o W���nQ W��nQ      E  , , Y���nQ Y���o Z���o Z���nQ Y���nQ      E  , , \���nQ \���o ]���o ]���nQ \���nQ      E  , , _���nQ _���o `{��o `{��nQ _���nQ      E  , , b���nQ b���o c_��o c_��nQ b���nQ      E  , , e{��nQ e{��o fC��o fC��nQ e{��nQ      E  , , h_��nQ h_��o i'��o i'��nQ h_��nQ      E  , , kC��nQ kC��o l��o l��nQ kC��nQ      E  , , n'��nQ n'��o n���o n���nQ n'��nQ      E  , , q��nQ q��o q���o q���nQ q��nQ      E  , , s���nQ s���o t���o t���nQ s���nQ      E  , , v���nQ v���o w���o w���nQ v���nQ      E  , , H���qq H���r9 I[��r9 I[��qq H���qq      E  , , Kw��qq Kw��r9 L?��r9 L?��qq Kw��qq      E  , , N[��qq N[��r9 O#��r9 O#��qq N[��qq      E  , , Q?��qq Q?��r9 R��r9 R��qq Q?��qq      E  , , H���l� H���m� I[��m� I[��l� H���l�      E  , , Kw��l� Kw��m� L?��m� L?��l� Kw��l�      E  , , N[��l� N[��m� O#��m� O#��l� N[��l�      E  , , Q?��l� Q?��m� R��m� R��l� Q?��l�      E  , , T#��l� T#��m� T���m� T���l� T#��l�      E  , , W��l� W��m� W���m� W���l� W��l�      E  , , Y���l� Y���m� Z���m� Z���l� Y���l�      E  , , \���l� \���m� ]���m� ]���l� \���l�      E  , , _���l� _���m� `{��m� `{��l� _���l�      E  , , b���l� b���m� c_��m� c_��l� b���l�      E  , , e{��l� e{��m� fC��m� fC��l� e{��l�      E  , , h_��l� h_��m� i'��m� i'��l� h_��l�      E  , , kC��l� kC��m� l��m� l��l� kC��l�      E  , , n'��l� n'��m� n���m� n���l� n'��l�      E  , , q��l� q��m� q���m� q���l� q��l�      E  , , s���l� s���m� t���m� t���l� s���l�      E  , , v���l� v���m� w���m� w���l� v���l�      E  , , T#��qq T#��r9 T���r9 T���qq T#��qq      E  , , W��qq W��r9 W���r9 W���qq W��qq      E  , , Y���qq Y���r9 Z���r9 Z���qq Y���qq      E  , , \���qq \���r9 ]���r9 ]���qq \���qq      E  , , _���qq _���r9 `{��r9 `{��qq _���qq      E  , , b���qq b���r9 c_��r9 c_��qq b���qq      E  , , e{��qq e{��r9 fC��r9 fC��qq e{��qq      E  , , h_��qq h_��r9 i'��r9 i'��qq h_��qq      E  , , H���o� H���p� I[��p� I[��o� H���o�      E  , , Kw��o� Kw��p� L?��p� L?��o� Kw��o�      E  , , N[��o� N[��p� O#��p� O#��o� N[��o�      E  , , H���k1 H���k� I[��k� I[��k1 H���k1      E  , , Kw��k1 Kw��k� L?��k� L?��k1 Kw��k1      E  , , N[��k1 N[��k� O#��k� O#��k1 N[��k1      E  , , Q?��k1 Q?��k� R��k� R��k1 Q?��k1      E  , , T#��k1 T#��k� T���k� T���k1 T#��k1      E  , , W��k1 W��k� W���k� W���k1 W��k1      E  , , Y���k1 Y���k� Z���k� Z���k1 Y���k1      E  , , \���k1 \���k� ]���k� ]���k1 \���k1      E  , , _���k1 _���k� `{��k� `{��k1 _���k1      E  , , b���k1 b���k� c_��k� c_��k1 b���k1      E  , , e{��k1 e{��k� fC��k� fC��k1 e{��k1      E  , , h_��k1 h_��k� i'��k� i'��k1 h_��k1      E  , , kC��k1 kC��k� l��k� l��k1 kC��k1      E  , , n'��k1 n'��k� n���k� n���k1 n'��k1      E  , , q��k1 q��k� q���k� q���k1 q��k1      E  , , s���k1 s���k� t���k� t���k1 s���k1      E  , , v���k1 v���k� w���k� w���k1 v���k1      E  , , Q?��o� Q?��p� R��p� R��o� Q?��o�      E  , , T#��o� T#��p� T���p� T���o� T#��o�      E  , , W��o� W��p� W���p� W���o� W��o�      E  , , Y���o� Y���p� Z���p� Z���o� Y���o�      E  , , B���l� B���m� C���m� C���l� B���l�      E  , , E���l� E���m� Fw��m� Fw��l� E���l�      E  , , "���nQ "���o #���o #���nQ "���nQ      E  , , %���nQ %���o &���o &���nQ %���nQ      E  , , (���nQ (���o )���o )���nQ (���nQ      E  , , +���nQ +���o ,s��o ,s��nQ +���nQ      E  , , .���nQ .���o /W��o /W��nQ .���nQ      E  , , 1s��nQ 1s��o 2;��o 2;��nQ 1s��nQ      E  , , 4W��nQ 4W��o 5��o 5��nQ 4W��nQ      E  , , 7;��nQ 7;��o 8��o 8��nQ 7;��nQ      E  , , :��nQ :��o :���o :���nQ :��nQ      E  , , =��nQ =��o =���o =���nQ =��nQ      E  , , ?���nQ ?���o @���o @���nQ ?���nQ      E  , , B���nQ B���o C���o C���nQ B���nQ      E  , , E���nQ E���o Fw��o Fw��nQ E���nQ      E  , , o��qq o��r9 7��r9 7��qq o��qq      E  , , S��qq S��r9 ��r9 ��qq S��qq      E  , , 7��qq 7��r9 ���r9 ���qq 7��qq      E  , ,  ��qq  ��r9  ���r9  ���qq  ��qq      E  , , "���qq "���r9 #���r9 #���qq "���qq      E  , , %���qq %���r9 &���r9 &���qq %���qq      E  , , (���qq (���r9 )���r9 )���qq (���qq      E  , , +���qq +���r9 ,s��r9 ,s��qq +���qq      E  , , .���qq .���r9 /W��r9 /W��qq .���qq      E  , , 1s��qq 1s��r9 2;��r9 2;��qq 1s��qq      E  , , 4W��qq 4W��r9 5��r9 5��qq 4W��qq      E  , , 7;��qq 7;��r9 8��r9 8��qq 7;��qq      E  , , o��o� o��p� 7��p� 7��o� o��o�      E  , , S��o� S��p� ��p� ��o� S��o�      E  , , 7��o� 7��p� ���p� ���o� 7��o�      E  , ,  ��o�  ��p�  ���p�  ���o�  ��o�      E  , , "���o� "���p� #���p� #���o� "���o�      E  , , %���o� %���p� &���p� &���o� %���o�      E  , , (���o� (���p� )���p� )���o� (���o�      E  , , +���o� +���p� ,s��p� ,s��o� +���o�      E  , , .���o� .���p� /W��p� /W��o� .���o�      E  , , 1s��o� 1s��p� 2;��p� 2;��o� 1s��o�      E  , , 4W��o� 4W��p� 5��p� 5��o� 4W��o�      E  , , 7;��o� 7;��p� 8��p� 8��o� 7;��o�      E  , , :��o� :��p� :���p� :���o� :��o�      E  , , =��o� =��p� =���p� =���o� =��o�      E  , , ?���o� ?���p� @���p� @���o� ?���o�      E  , , B���o� B���p� C���p� C���o� B���o�      E  , , E���o� E���p� Fw��p� Fw��o� E���o�      E  , , :��qq :��r9 :���r9 :���qq :��qq      E  , , =��qq =��r9 =���r9 =���qq =��qq      E  , , ?���qq ?���r9 @���r9 @���qq ?���qq      E  , , o��k1 o��k� 7��k� 7��k1 o��k1      E  , , S��k1 S��k� ��k� ��k1 S��k1      E  , , 7��k1 7��k� ���k� ���k1 7��k1      E  , ,  ��k1  ��k�  ���k�  ���k1  ��k1      E  , , "���k1 "���k� #���k� #���k1 "���k1      E  , , %���k1 %���k� &���k� &���k1 %���k1      E  , , (���k1 (���k� )���k� )���k1 (���k1      E  , , +���k1 +���k� ,s��k� ,s��k1 +���k1      E  , , .���k1 .���k� /W��k� /W��k1 .���k1      E  , , 1s��k1 1s��k� 2;��k� 2;��k1 1s��k1      E  , , 4W��k1 4W��k� 5��k� 5��k1 4W��k1      E  , , 7;��k1 7;��k� 8��k� 8��k1 7;��k1      E  , , :��k1 :��k� :���k� :���k1 :��k1      E  , , =��k1 =��k� =���k� =���k1 =��k1      E  , , ?���k1 ?���k� @���k� @���k1 ?���k1      E  , , B���k1 B���k� C���k� C���k1 B���k1      E  , , E���k1 E���k� Fw��k� Fw��k1 E���k1      E  , , B���qq B���r9 C���r9 C���qq B���qq      E  , , E���qq E���r9 Fw��r9 Fw��qq E���qq      E  , , o��nQ o��o 7��o 7��nQ o��nQ      E  , , S��nQ S��o ��o ��nQ S��nQ      E  , , 7��nQ 7��o ���o ���nQ 7��nQ      E  , ,  ��nQ  ��o  ���o  ���nQ  ��nQ      E  , , o��l� o��m� 7��m� 7��l� o��l�      E  , , S��l� S��m� ��m� ��l� S��l�      E  , , 7��l� 7��m� ���m� ���l� 7��l�      E  , ,  ��l�  ��m�  ���m�  ���l�  ��l�      E  , , "���l� "���m� #���m� #���l� "���l�      E  , , %���l� %���m� &���m� &���l� %���l�      E  , , (���l� (���m� )���m� )���l� (���l�      E  , , +���l� +���m� ,s��m� ,s��l� +���l�      E  , , .���l� .���m� /W��m� /W��l� .���l�      E  , , 1s��l� 1s��m� 2;��m� 2;��l� 1s��l�      E  , , 4W��l� 4W��m� 5��m� 5��l� 4W��l�      E  , , 7;��l� 7;��m� 8��m� 8��l� 7;��l�      E  , , :��l� :��m� :���m� :���l� :��l�      E  , , =��l� =��m� =���m� =���l� =��l�      E  , , ?���l� ?���m� @���m� @���l� ?���l�      E  , , :��[ :��[� :���[� :���[ :��[      E  , , =��[ =��[� =���[� =���[ =��[      E  , , ?���[ ?���[� @���[� @���[ ?���[      E  , , B���[ B���[� C���[� C���[ B���[      E  , , E���[ E���[� Fw��[� Fw��[ E���[      E  , , o��[ o��[� 7��[� 7��[ o��[      E  , , S��[ S��[� ��[� ��[ S��[      E  , , 7��[ 7��[� ���[� ���[ 7��[      E  , ,  ��[  ��[�  ���[�  ���[  ��[      E  , , "���[ "���[� #���[� #���[ "���[      E  , , %���[ %���[� &���[� &���[ %���[      E  , , (���[ (���[� )���[� )���[ (���[      E  , , +���[ +���[� ,s��[� ,s��[ +���[      E  , , .���[ .���[� /W��[� /W��[ .���[      E  , , 1s��[ 1s��[� 2;��[� 2;��[ 1s��[      E  , , 4W��[ 4W��[� 5��[� 5��[ 4W��[      E  , , 7;��[ 7;��[� 8��[� 8��[ 7;��[      E  , , 7;��f� 7;��gI 8��gI 8��f� 7;��f�      E  , , :��f� :��gI :���gI :���f� :��f�      E  , , =��f� =��gI =���gI =���f� =��f�      E  , , ?���f� ?���gI @���gI @���f� ?���f�      E  , , B���f� B���gI C���gI C���f� B���f�      E  , , E���f� E���gI Fw��gI Fw��f� E���f�      E  , , .���d� .���e� /W��e� /W��d� .���d�      E  , , 1s��d� 1s��e� 2;��e� 2;��d� 1s��d�      E  , , 4W��d� 4W��e� 5��e� 5��d� 4W��d�      E  , , 7;��d� 7;��e� 8��e� 8��d� 7;��d�      E  , , :��d� :��e� :���e� :���d� :��d�      E  , , =��d� =��e� =���e� =���d� =��d�      E  , , ?���d� ?���e� @���e� @���d� ?���d�      E  , , B���d� B���e� C���e� C���d� B���d�      E  , , E���d� E���e� Fw��e� Fw��d� E���d�      E  , , .���h .���h� /W��h� /W��h .���h      E  , , 1s��h 1s��h� 2;��h� 2;��h 1s��h      E  , , 4W��h 4W��h� 5��h� 5��h 4W��h      E  , , 7;��h 7;��h� 8��h� 8��h 7;��h      E  , , :��h :��h� :���h� :���h :��h      E  , , =��h =��h� =���h� =���h =��h      E  , , ?���h ?���h� @���h� @���h ?���h      E  , , B���h B���h� C���h� C���h B���h      E  , , E���h E���h� Fw��h� Fw��h E���h      E  , , .���ca .���d) /W��d) /W��ca .���ca      E  , , 1s��ca 1s��d) 2;��d) 2;��ca 1s��ca      E  , , 4W��ca 4W��d) 5��d) 5��ca 4W��ca      E  , , 7;��ca 7;��d) 8��d) 8��ca 7;��ca      E  , , :��ca :��d) :���d) :���ca :��ca      E  , , =��ca =��d) =���d) =���ca =��ca      E  , , ?���ca ?���d) @���d) @���ca ?���ca      E  , , B���ca B���d) C���d) C���ca B���ca      E  , , E���ca E���d) Fw��d) Fw��ca E���ca      E  , , .���f� .���gI /W��gI /W��f� .���f�      E  , , 1s��f� 1s��gI 2;��gI 2;��f� 1s��f�      E  , , 4W��f� 4W��gI 5��gI 5��f� 4W��f�      E  , , "���f� "���gI #���gI #���f� "���f�      E  , , %���f� %���gI &���gI &���f� %���f�      E  , , (���f� (���gI )���gI )���f� (���f�      E  , , +���f� +���gI ,s��gI ,s��f� +���f�      E  , , o��h o��h� 7��h� 7��h o��h      E  , , S��h S��h� ��h� ��h S��h      E  , , 7��h 7��h� ���h� ���h 7��h      E  , ,  ��h  ��h�  ���h�  ���h  ��h      E  , , "���h "���h� #���h� #���h "���h      E  , , %���h %���h� &���h� &���h %���h      E  , , (���h (���h� )���h� )���h (���h      E  , , +���h +���h� ,s��h� ,s��h +���h      E  , , o��d� o��e� 7��e� 7��d� o��d�      E  , , o��f� o��gI 7��gI 7��f� o��f�      E  , , S��f� S��gI ��gI ��f� S��f�      E  , , 7��f� 7��gI ���gI ���f� 7��f�      E  , , o��ca o��d) 7��d) 7��ca o��ca      E  , , S��ca S��d) ��d) ��ca S��ca      E  , , 7��ca 7��d) ���d) ���ca 7��ca      E  , ,  ��ca  ��d)  ���d)  ���ca  ��ca      E  , , S��d� S��e� ��e� ��d� S��d�      E  , , 7��d� 7��e� ���e� ���d� 7��d�      E  , ,  ��d�  ��e�  ���e�  ���d�  ��d�      E  , , "���d� "���e� #���e� #���d� "���d�      E  , , %���d� %���e� &���e� &���d� %���d�      E  , , (���d� (���e� )���e� )���d� (���d�      E  , , +���d� +���e� ,s��e� ,s��d� +���d�      E  , , %���ca %���d) &���d) &���ca %���ca      E  , , (���ca (���d) )���d) )���ca (���ca      E  , , +���ca +���d) ,s��d) ,s��ca +���ca      E  , , "���ca "���d) #���d) #���ca "���ca      E  , ,  ��f�  ��gI  ���gI  ���f�  ��f�      E  , , (���T� (���U� )���U� )���T� (���T�      E  , , +���T� +���U� ,s��U� ,s��T� +���T�      E  , , o��W� o��X� 7��X� 7��W� o��W�      E  , , S��W� S��X� ��X� ��W� S��W�      E  , , 7��W� 7��X� ���X� ���W� 7��W�      E  , ,  ��W�  ��X�  ���X�  ���W�  ��W�      E  , , o��V_ o��W' 7��W' 7��V_ o��V_      E  , , S��V_ S��W' ��W' ��V_ S��V_      E  , , 7��V_ 7��W' ���W' ���V_ 7��V_      E  , ,  ��V_  ��W'  ���W'  ���V_  ��V_      E  , , "���V_ "���W' #���W' #���V_ "���V_      E  , , %���V_ %���W' &���W' &���V_ %���V_      E  , , (���V_ (���W' )���W' )���V_ (���V_      E  , , +���V_ +���W' ,s��W' ,s��V_ +���V_      E  , , o��S? o��T 7��T 7��S? o��S?      E  , , S��S? S��T ��T ��S? S��S?      E  , , 7��S? 7��T ���T ���S? 7��S?      E  , ,  ��S?  ��T  ���T  ���S?  ��S?      E  , , "���S? "���T #���T #���S? "���S?      E  , , %���S? %���T &���T &���S? %���S?      E  , , (���S? (���T )���T )���S? (���S?      E  , , +���S? +���T ,s��T ,s��S? +���S?      E  , , "���W� "���X� #���X� #���W� "���W�      E  , , %���W� %���X� &���X� &���W� %���W�      E  , , (���W� (���X� )���X� )���W� (���W�      E  , , +���W� +���X� ,s��X� ,s��W� +���W�      E  , , "���Y "���ZG #���ZG #���Y "���Y      E  , , %���Y %���ZG &���ZG &���Y %���Y      E  , , (���Y (���ZG )���ZG )���Y (���Y      E  , , +���Y +���ZG ,s��ZG ,s��Y +���Y      E  , , o��Y o��ZG 7��ZG 7��Y o��Y      E  , , S��Y S��ZG ��ZG ��Y S��Y      E  , , 7��Y 7��ZG ���ZG ���Y 7��Y      E  , ,  ��Y  ��ZG  ���ZG  ���Y  ��Y      E  , , o��Q� o��Rw 7��Rw 7��Q� o��Q�      E  , , S��Q� S��Rw ��Rw ��Q� S��Q�      E  , , 7��Q� 7��Rw ���Rw ���Q� 7��Q�      E  , ,  ��Q�  ��Rw  ���Rw  ���Q�  ��Q�      E  , , "���Q� "���Rw #���Rw #���Q� "���Q�      E  , , %���Q� %���Rw &���Rw &���Q� %���Q�      E  , , (���Q� (���Rw )���Rw )���Q� (���Q�      E  , , +���Q� +���Rw ,s��Rw ,s��Q� +���Q�      E  , , o��T� o��U� 7��U� 7��T� o��T�      E  , , S��T� S��U� ��U� ��T� S��T�      E  , , o��P o��P� 7��P� 7��P o��P      E  , , S��P S��P� ��P� ��P S��P      E  , , 7��P 7��P� ���P� ���P 7��P      E  , ,  ��P  ��P�  ���P�  ���P  ��P      E  , , "���P "���P� #���P� #���P "���P      E  , , %���P %���P� &���P� &���P %���P      E  , , (���P (���P� )���P� )���P (���P      E  , , +���P +���P� ,s��P� ,s��P +���P      E  , , o��N� o��OW 7��OW 7��N� o��N�      E  , , S��N� S��OW ��OW ��N� S��N�      E  , , 7��N� 7��OW ���OW ���N� 7��N�      E  , ,  ��N�  ��OW  ���OW  ���N�  ��N�      E  , , "���N� "���OW #���OW #���N� "���N�      E  , , %���N� %���OW &���OW &���N� %���N�      E  , , (���N� (���OW )���OW )���N� (���N�      E  , , +���N� +���OW ,s��OW ,s��N� +���N�      E  , , 7��T� 7��U� ���U� ���T� 7��T�      E  , ,  ��T�  ��U�  ���U�  ���T�  ��T�      E  , , "���T� "���U� #���U� #���T� "���T�      E  , , %���T� %���U� &���U� &���T� %���T�      E  , , o��L� o��M� 7��M� 7��L� o��L�      E  , , S��L� S��M� ��M� ��L� S��L�      E  , , 7��L� 7��M� ���M� ���L� 7��L�      E  , ,  ��L�  ��M�  ���M�  ���L�  ��L�      E  , , "���L� "���M� #���M� #���L� "���L�      E  , , %���L� %���M� &���M� &���L� %���L�      E  , , (���L� (���M� )���M� )���L� (���L�      E  , , +���L� +���M� ,s��M� ,s��L� +���L�      E  , , .���V_ .���W' /W��W' /W��V_ .���V_      E  , , 1s��V_ 1s��W' 2;��W' 2;��V_ 1s��V_      E  , , .���T� .���U� /W��U� /W��T� .���T�      E  , , 1s��T� 1s��U� 2;��U� 2;��T� 1s��T�      E  , , 4W��T� 4W��U� 5��U� 5��T� 4W��T�      E  , , 7;��T� 7;��U� 8��U� 8��T� 7;��T�      E  , , :��T� :��U� :���U� :���T� :��T�      E  , , =��T� =��U� =���U� =���T� =��T�      E  , , ?���T� ?���U� @���U� @���T� ?���T�      E  , , B���T� B���U� C���U� C���T� B���T�      E  , , E���T� E���U� Fw��U� Fw��T� E���T�      E  , , 4W��V_ 4W��W' 5��W' 5��V_ 4W��V_      E  , , 7;��V_ 7;��W' 8��W' 8��V_ 7;��V_      E  , , :��V_ :��W' :���W' :���V_ :��V_      E  , , =��V_ =��W' =���W' =���V_ =��V_      E  , , .���Q� .���Rw /W��Rw /W��Q� .���Q�      E  , , 1s��Q� 1s��Rw 2;��Rw 2;��Q� 1s��Q�      E  , , 4W��Q� 4W��Rw 5��Rw 5��Q� 4W��Q�      E  , , 7;��Q� 7;��Rw 8��Rw 8��Q� 7;��Q�      E  , , :��Q� :��Rw :���Rw :���Q� :��Q�      E  , , =��Q� =��Rw =���Rw =���Q� =��Q�      E  , , ?���Q� ?���Rw @���Rw @���Q� ?���Q�      E  , , B���Q� B���Rw C���Rw C���Q� B���Q�      E  , , E���Q� E���Rw Fw��Rw Fw��Q� E���Q�      E  , , ?���V_ ?���W' @���W' @���V_ ?���V_      E  , , B���V_ B���W' C���W' C���V_ B���V_      E  , , E���V_ E���W' Fw��W' Fw��V_ E���V_      E  , , :��Y :��ZG :���ZG :���Y :��Y      E  , , =��Y =��ZG =���ZG =���Y =��Y      E  , , ?���Y ?���ZG @���ZG @���Y ?���Y      E  , , B���Y B���ZG C���ZG C���Y B���Y      E  , , E���Y E���ZG Fw��ZG Fw��Y E���Y      E  , , .���Y .���ZG /W��ZG /W��Y .���Y      E  , , 1s��Y 1s��ZG 2;��ZG 2;��Y 1s��Y      E  , , .���P .���P� /W��P� /W��P .���P      E  , , 1s��P 1s��P� 2;��P� 2;��P 1s��P      E  , , 4W��P 4W��P� 5��P� 5��P 4W��P      E  , , 7;��P 7;��P� 8��P� 8��P 7;��P      E  , , :��P :��P� :���P� :���P :��P      E  , , =��P =��P� =���P� =���P =��P      E  , , ?���P ?���P� @���P� @���P ?���P      E  , , B���P B���P� C���P� C���P B���P      E  , , E���P E���P� Fw��P� Fw��P E���P      E  , , .���W� .���X� /W��X� /W��W� .���W�      E  , , 1s��W� 1s��X� 2;��X� 2;��W� 1s��W�      E  , , 4W��W� 4W��X� 5��X� 5��W� 4W��W�      E  , , 7;��W� 7;��X� 8��X� 8��W� 7;��W�      E  , , :��W� :��X� :���X� :���W� :��W�      E  , , =��W� =��X� =���X� =���W� =��W�      E  , , .���S? .���T /W��T /W��S? .���S?      E  , , 1s��S? 1s��T 2;��T 2;��S? 1s��S?      E  , , .���N� .���OW /W��OW /W��N� .���N�      E  , , 1s��N� 1s��OW 2;��OW 2;��N� 1s��N�      E  , , 4W��N� 4W��OW 5��OW 5��N� 4W��N�      E  , , 7;��N� 7;��OW 8��OW 8��N� 7;��N�      E  , , :��N� :��OW :���OW :���N� :��N�      E  , , =��N� =��OW =���OW =���N� =��N�      E  , , ?���N� ?���OW @���OW @���N� ?���N�      E  , , B���N� B���OW C���OW C���N� B���N�      E  , , E���N� E���OW Fw��OW Fw��N� E���N�      E  , , 4W��S? 4W��T 5��T 5��S? 4W��S?      E  , , 7;��S? 7;��T 8��T 8��S? 7;��S?      E  , , :��S? :��T :���T :���S? :��S?      E  , , =��S? =��T =���T =���S? =��S?      E  , , ?���S? ?���T @���T @���S? ?���S?      E  , , B���S? B���T C���T C���S? B���S?      E  , , E���S? E���T Fw��T Fw��S? E���S?      E  , , ?���W� ?���X� @���X� @���W� ?���W�      E  , , B���W� B���X� C���X� C���W� B���W�      E  , , E���W� E���X� Fw��X� Fw��W� E���W�      E  , , 4W��Y 4W��ZG 5��ZG 5��Y 4W��Y      E  , , 7;��Y 7;��ZG 8��ZG 8��Y 7;��Y      E  , , .���L� .���M� /W��M� /W��L� .���L�      E  , , 1s��L� 1s��M� 2;��M� 2;��L� 1s��L�      E  , , 4W��L� 4W��M� 5��M� 5��L� 4W��L�      E  , , 7;��L� 7;��M� 8��M� 8��L� 7;��L�      E  , , :��L� :��M� :���M� :���L� :��L�      E  , , =��L� =��M� =���M� =���L� =��L�      E  , , ?���L� ?���M� @���M� @���L� ?���L�      E  , , B���L� B���M� C���M� C���L� B���L�      E  , , E���L� E���M� Fw��M� Fw��L� E���L�      E  , , H���[ H���[� I[��[� I[��[ H���[      E  , , Kw��[ Kw��[� L?��[� L?��[ Kw��[      E  , , N[��[ N[��[� O#��[� O#��[ N[��[      E  , , Q?��[ Q?��[� R��[� R��[ Q?��[      E  , , T#��[ T#��[� T���[� T���[ T#��[      E  , , W��[ W��[� W���[� W���[ W��[      E  , , Y���[ Y���[� Z���[� Z���[ Y���[      E  , , \���[ \���[� ]���[� ]���[ \���[      E  , , _���[ _���[� `{��[� `{��[ _���[      E  , , b���[ b���[� c_��[� c_��[ b���[      E  , , e{��[ e{��[� fC��[� fC��[ e{��[      E  , , h_��[ h_��[� i'��[� i'��[ h_��[      E  , , kC��[ kC��[� l��[� l��[ kC��[      E  , , n'��[ n'��[� n���[� n���[ n'��[      E  , , q��[ q��[� q���[� q���[ q��[      E  , , s���[ s���[� t���[� t���[ s���[      E  , , v���[ v���[� w���[� w���[ v���[      E  , , e{��h e{��h� fC��h� fC��h e{��h      E  , , h_��h h_��h� i'��h� i'��h h_��h      E  , , kC��h kC��h� l��h� l��h kC��h      E  , , n'��h n'��h� n���h� n���h n'��h      E  , , q��h q��h� q���h� q���h q��h      E  , , s���h s���h� t���h� t���h s���h      E  , , v���h v���h� w���h� w���h v���h      E  , , _���ca _���d) `{��d) `{��ca _���ca      E  , , b���ca b���d) c_��d) c_��ca b���ca      E  , , e{��ca e{��d) fC��d) fC��ca e{��ca      E  , , h_��ca h_��d) i'��d) i'��ca h_��ca      E  , , kC��ca kC��d) l��d) l��ca kC��ca      E  , , n'��ca n'��d) n���d) n���ca n'��ca      E  , , q��ca q��d) q���d) q���ca q��ca      E  , , s���ca s���d) t���d) t���ca s���ca      E  , , v���ca v���d) w���d) w���ca v���ca      E  , , h_��d� h_��e� i'��e� i'��d� h_��d�      E  , , kC��d� kC��e� l��e� l��d� kC��d�      E  , , n'��d� n'��e� n���e� n���d� n'��d�      E  , , q��d� q��e� q���e� q���d� q��d�      E  , , s���d� s���e� t���e� t���d� s���d�      E  , , v���d� v���e� w���e� w���d� v���d�      E  , , _���f� _���gI `{��gI `{��f� _���f�      E  , , b���f� b���gI c_��gI c_��f� b���f�      E  , , e{��f� e{��gI fC��gI fC��f� e{��f�      E  , , h_��f� h_��gI i'��gI i'��f� h_��f�      E  , , kC��f� kC��gI l��gI l��f� kC��f�      E  , , n'��f� n'��gI n���gI n���f� n'��f�      E  , , q��f� q��gI q���gI q���f� q��f�      E  , , s���f� s���gI t���gI t���f� s���f�      E  , , v���f� v���gI w���gI w���f� v���f�      E  , , _���h _���h� `{��h� `{��h _���h      E  , , b���h b���h� c_��h� c_��h b���h      E  , , _���d� _���e� `{��e� `{��d� _���d�      E  , , b���d� b���e� c_��e� c_��d� b���d�      E  , , e{��d� e{��e� fC��e� fC��d� e{��d�      E  , , T#��f� T#��gI T���gI T���f� T#��f�      E  , , W��f� W��gI W���gI W���f� W��f�      E  , , Y���f� Y���gI Z���gI Z���f� Y���f�      E  , , Kw��f� Kw��gI L?��gI L?��f� Kw��f�      E  , , N[��f� N[��gI O#��gI O#��f� N[��f�      E  , , H���ca H���d) I[��d) I[��ca H���ca      E  , , Kw��ca Kw��d) L?��d) L?��ca Kw��ca      E  , , N[��ca N[��d) O#��d) O#��ca N[��ca      E  , , Q?��ca Q?��d) R��d) R��ca Q?��ca      E  , , T#��ca T#��d) T���d) T���ca T#��ca      E  , , W��ca W��d) W���d) W���ca W��ca      E  , , Y���ca Y���d) Z���d) Z���ca Y���ca      E  , , \���ca \���d) ]���d) ]���ca \���ca      E  , , Kw��h Kw��h� L?��h� L?��h Kw��h      E  , , N[��h N[��h� O#��h� O#��h N[��h      E  , , Q?��h Q?��h� R��h� R��h Q?��h      E  , , T#��h T#��h� T���h� T���h T#��h      E  , , W��h W��h� W���h� W���h W��h      E  , , Y���h Y���h� Z���h� Z���h Y���h      E  , , \���h \���h� ]���h� ]���h \���h      E  , , \���f� \���gI ]���gI ]���f� \���f�      E  , , H���d� H���e� I[��e� I[��d� H���d�      E  , , Kw��d� Kw��e� L?��e� L?��d� Kw��d�      E  , , N[��d� N[��e� O#��e� O#��d� N[��d�      E  , , Q?��d� Q?��e� R��e� R��d� Q?��d�      E  , , T#��d� T#��e� T���e� T���d� T#��d�      E  , , W��d� W��e� W���e� W���d� W��d�      E  , , Y���d� Y���e� Z���e� Z���d� Y���d�      E  , , \���d� \���e� ]���e� ]���d� \���d�      E  , , H���h H���h� I[��h� I[��h H���h      E  , , H���f� H���gI I[��gI I[��f� H���f�      E  , , Q?��f� Q?��gI R��gI R��f� Q?��f�      E  , , W��Q� W��Rw W���Rw W���Q� W��Q�      E  , , Y���Q� Y���Rw Z���Rw Z���Q� Y���Q�      E  , , \���Q� \���Rw ]���Rw ]���Q� \���Q�      E  , , W��Y W��ZG W���ZG W���Y W��Y      E  , , H���S? H���T I[��T I[��S? H���S?      E  , , Kw��S? Kw��T L?��T L?��S? Kw��S?      E  , , N[��S? N[��T O#��T O#��S? N[��S?      E  , , Q?��S? Q?��T R��T R��S? Q?��S?      E  , , T#��S? T#��T T���T T���S? T#��S?      E  , , W��S? W��T W���T W���S? W��S?      E  , , Y���S? Y���T Z���T Z���S? Y���S?      E  , , \���S? \���T ]���T ]���S? \���S?      E  , , Y���Y Y���ZG Z���ZG Z���Y Y���Y      E  , , \���Y \���ZG ]���ZG ]���Y \���Y      E  , , H���Y H���ZG I[��ZG I[��Y H���Y      E  , , Kw��Y Kw��ZG L?��ZG L?��Y Kw��Y      E  , , H���T� H���U� I[��U� I[��T� H���T�      E  , , Kw��T� Kw��U� L?��U� L?��T� Kw��T�      E  , , N[��T� N[��U� O#��U� O#��T� N[��T�      E  , , H���P H���P� I[��P� I[��P H���P      E  , , Kw��P Kw��P� L?��P� L?��P Kw��P      E  , , N[��P N[��P� O#��P� O#��P N[��P      E  , , Q?��P Q?��P� R��P� R��P Q?��P      E  , , T#��P T#��P� T���P� T���P T#��P      E  , , W��P W��P� W���P� W���P W��P      E  , , Y���P Y���P� Z���P� Z���P Y���P      E  , , \���P \���P� ]���P� ]���P \���P      E  , , Q?��T� Q?��U� R��U� R��T� Q?��T�      E  , , T#��T� T#��U� T���U� T���T� T#��T�      E  , , W��T� W��U� W���U� W���T� W��T�      E  , , Y���T� Y���U� Z���U� Z���T� Y���T�      E  , , \���T� \���U� ]���U� ]���T� \���T�      E  , , N[��Y N[��ZG O#��ZG O#��Y N[��Y      E  , , Q?��Y Q?��ZG R��ZG R��Y Q?��Y      E  , , T#��Y T#��ZG T���ZG T���Y T#��Y      E  , , H���W� H���X� I[��X� I[��W� H���W�      E  , , Kw��W� Kw��X� L?��X� L?��W� Kw��W�      E  , , N[��W� N[��X� O#��X� O#��W� N[��W�      E  , , Q?��W� Q?��X� R��X� R��W� Q?��W�      E  , , T#��W� T#��X� T���X� T���W� T#��W�      E  , , H���V_ H���W' I[��W' I[��V_ H���V_      E  , , Kw��V_ Kw��W' L?��W' L?��V_ Kw��V_      E  , , N[��V_ N[��W' O#��W' O#��V_ N[��V_      E  , , Q?��V_ Q?��W' R��W' R��V_ Q?��V_      E  , , H���N� H���OW I[��OW I[��N� H���N�      E  , , Kw��N� Kw��OW L?��OW L?��N� Kw��N�      E  , , N[��N� N[��OW O#��OW O#��N� N[��N�      E  , , Q?��N� Q?��OW R��OW R��N� Q?��N�      E  , , T#��N� T#��OW T���OW T���N� T#��N�      E  , , W��N� W��OW W���OW W���N� W��N�      E  , , Y���N� Y���OW Z���OW Z���N� Y���N�      E  , , \���N� \���OW ]���OW ]���N� \���N�      E  , , T#��V_ T#��W' T���W' T���V_ T#��V_      E  , , W��V_ W��W' W���W' W���V_ W��V_      E  , , Y���V_ Y���W' Z���W' Z���V_ Y���V_      E  , , \���V_ \���W' ]���W' ]���V_ \���V_      E  , , W��W� W��X� W���X� W���W� W��W�      E  , , Y���W� Y���X� Z���X� Z���W� Y���W�      E  , , \���W� \���X� ]���X� ]���W� \���W�      E  , , H���Q� H���Rw I[��Rw I[��Q� H���Q�      E  , , Kw��Q� Kw��Rw L?��Rw L?��Q� Kw��Q�      E  , , N[��Q� N[��Rw O#��Rw O#��Q� N[��Q�      E  , , Q?��Q� Q?��Rw R��Rw R��Q� Q?��Q�      E  , , T#��Q� T#��Rw T���Rw T���Q� T#��Q�      E  , , H���L� H���M� I[��M� I[��L� H���L�      E  , , Kw��L� Kw��M� L?��M� L?��L� Kw��L�      E  , , N[��L� N[��M� O#��M� O#��L� N[��L�      E  , , Q?��L� Q?��M� R��M� R��L� Q?��L�      E  , , T#��L� T#��M� T���M� T���L� T#��L�      E  , , W��L� W��M� W���M� W���L� W��L�      E  , , Y���L� Y���M� Z���M� Z���L� Y���L�      E  , , \���L� \���M� ]���M� ]���L� \���L�      E  , , _���P _���P� `{��P� `{��P _���P      E  , , b���P b���P� c_��P� c_��P b���P      E  , , e{��P e{��P� fC��P� fC��P e{��P      E  , , h_��P h_��P� i'��P� i'��P h_��P      E  , , kC��P kC��P� l��P� l��P kC��P      E  , , n'��P n'��P� n���P� n���P n'��P      E  , , q��P q��P� q���P� q���P q��P      E  , , s���P s���P� t���P� t���P s���P      E  , , v���P v���P� w���P� w���P v���P      E  , , n'��W� n'��X� n���X� n���W� n'��W�      E  , , n'��S? n'��T n���T n���S? n'��S?      E  , , q��S? q��T q���T q���S? q��S?      E  , , s���S? s���T t���T t���S? s���S?      E  , , v���S? v���T w���T w���S? v���S?      E  , , b���T� b���U� c_��U� c_��T� b���T�      E  , , e{��T� e{��U� fC��U� fC��T� e{��T�      E  , , h_��T� h_��U� i'��U� i'��T� h_��T�      E  , , kC��T� kC��U� l��U� l��T� kC��T�      E  , , _���Q� _���Rw `{��Rw `{��Q� _���Q�      E  , , b���Q� b���Rw c_��Rw c_��Q� b���Q�      E  , , e{��Q� e{��Rw fC��Rw fC��Q� e{��Q�      E  , , h_��Q� h_��Rw i'��Rw i'��Q� h_��Q�      E  , , kC��Q� kC��Rw l��Rw l��Q� kC��Q�      E  , , n'��Q� n'��Rw n���Rw n���Q� n'��Q�      E  , , q��Q� q��Rw q���Rw q���Q� q��Q�      E  , , s���Q� s���Rw t���Rw t���Q� s���Q�      E  , , v���Q� v���Rw w���Rw w���Q� v���Q�      E  , , q��W� q��X� q���X� q���W� q��W�      E  , , s���W� s���X� t���X� t���W� s���W�      E  , , v���W� v���X� w���X� w���W� v���W�      E  , , n'��T� n'��U� n���U� n���T� n'��T�      E  , , _���Y _���ZG `{��ZG `{��Y _���Y      E  , , b���Y b���ZG c_��ZG c_��Y b���Y      E  , , e{��Y e{��ZG fC��ZG fC��Y e{��Y      E  , , _���N� _���OW `{��OW `{��N� _���N�      E  , , b���N� b���OW c_��OW c_��N� b���N�      E  , , e{��N� e{��OW fC��OW fC��N� e{��N�      E  , , h_��N� h_��OW i'��OW i'��N� h_��N�      E  , , kC��N� kC��OW l��OW l��N� kC��N�      E  , , n'��N� n'��OW n���OW n���N� n'��N�      E  , , q��N� q��OW q���OW q���N� q��N�      E  , , s���N� s���OW t���OW t���N� s���N�      E  , , v���N� v���OW w���OW w���N� v���N�      E  , , h_��Y h_��ZG i'��ZG i'��Y h_��Y      E  , , kC��Y kC��ZG l��ZG l��Y kC��Y      E  , , n'��Y n'��ZG n���ZG n���Y n'��Y      E  , , q��Y q��ZG q���ZG q���Y q��Y      E  , , _���V_ _���W' `{��W' `{��V_ _���V_      E  , , b���V_ b���W' c_��W' c_��V_ b���V_      E  , , e{��V_ e{��W' fC��W' fC��V_ e{��V_      E  , , h_��V_ h_��W' i'��W' i'��V_ h_��V_      E  , , kC��V_ kC��W' l��W' l��V_ kC��V_      E  , , n'��V_ n'��W' n���W' n���V_ n'��V_      E  , , q��V_ q��W' q���W' q���V_ q��V_      E  , , s���V_ s���W' t���W' t���V_ s���V_      E  , , v���V_ v���W' w���W' w���V_ v���V_      E  , , s���Y s���ZG t���ZG t���Y s���Y      E  , , v���Y v���ZG w���ZG w���Y v���Y      E  , , q��T� q��U� q���U� q���T� q��T�      E  , , s���T� s���U� t���U� t���T� s���T�      E  , , v���T� v���U� w���U� w���T� v���T�      E  , , _���T� _���U� `{��U� `{��T� _���T�      E  , , _���S? _���T `{��T `{��S? _���S?      E  , , b���S? b���T c_��T c_��S? b���S?      E  , , e{��S? e{��T fC��T fC��S? e{��S?      E  , , h_��S? h_��T i'��T i'��S? h_��S?      E  , , kC��S? kC��T l��T l��S? kC��S?      E  , , _���W� _���X� `{��X� `{��W� _���W�      E  , , b���W� b���X� c_��X� c_��W� b���W�      E  , , e{��W� e{��X� fC��X� fC��W� e{��W�      E  , , h_��W� h_��X� i'��X� i'��W� h_��W�      E  , , kC��W� kC��X� l��X� l��W� kC��W�      E  , , _���L� _���M� `{��M� `{��L� _���L�      E  , , b���L� b���M� c_��M� c_��L� b���L�      E  , , e{��L� e{��M� fC��M� fC��L� e{��L�      E  , , h_��L� h_��M� i'��M� i'��L� h_��L�      E  , , kC��L� kC��M� l��M� l��L� kC��L�      E  , , n'��L� n'��M� n���M� n���L� n'��L�      E  , , q��L� q��M� q���M� q���L� q��L�      E  , , s���L� s���M� t���M� t���L� s���L�      E  , , v���L� v���M� w���M� w���L� v���L�      E  , , ����i� ����ji ����ji ����i� ����i�      E  , , ����i� ����ji ŧ��ji ŧ��i� ����i�      E  , , ����i� ����ji ȋ��ji ȋ��i� ����i�      E  , , ʧ��i� ʧ��ji �o��ji �o��i� ʧ��i�      E  , , ͋��i� ͋��ji �S��ji �S��i� ͋��i�      E  , , y���i� y���ji z��ji z��i� y���i�      E  , , |���i� |���ji }c��ji }c��i� |���i�      E  , , ��i� ��ji �G��ji �G��i� ��i�      E  , , �c��i� �c��ji �+��ji �+��i� �c��i�      E  , , �G��i� �G��ji ���ji ���i� �G��i�      E  , , �+��i� �+��ji ����ji ����i� �+��i�      E  , , ���i� ���ji ����ji ����i� ���i�      E  , , ����i� ����ji ����ji ����i� ����i�      E  , , ����i� ����ji ����ji ����i� ����i�      E  , , ����i� ����ji ����ji ����i� ����i�      E  , , ����i� ����ji �g��ji �g��i� ����i�      E  , , ����i� ����ji �K��ji �K��i� ����i�      E  , , �g��i� �g��ji �/��ji �/��i� �g��i�      E  , , �K��i� �K��ji ���ji ���i� �K��i�      E  , , �/��i� �/��ji ����ji ����i� �/��i�      E  , , ���i� ���ji ����ji ����i� ���i�      E  , , ����i� ����ji ����ji ����i� ����i�      E  , , ����i� ����ji ����ji ����i� ����i�      E  , , ����i� ����ji ����ji ����i� ����i�      E  , , ����i� ����ji �k��ji �k��i� ����i�      E  , , ����i� ����ji �O��ji �O��i� ����i�      E  , , �k��i� �k��ji �3��ji �3��i� �k��i�      E  , , �O��i� �O��ji ���ji ���i� �O��i�      E  , , �3��i� �3��ji ����ji ����i� �3��i�      E  , , ���i� ���ji ����ji ����i� ���i�      E  , , ʧ��o� ʧ��p� �o��p� �o��o� ʧ��o�      E  , , ͋��o� ͋��p� �S��p� �S��o� ͋��o�      E  , , ����nQ ����o ����o ����nQ ����nQ      E  , , ����nQ ����o ����o ����nQ ����nQ      E  , , ����nQ ����o �k��o �k��nQ ����nQ      E  , , ����nQ ����o �O��o �O��nQ ����nQ      E  , , �k��nQ �k��o �3��o �3��nQ �k��nQ      E  , , �O��nQ �O��o ���o ���nQ �O��nQ      E  , , �3��nQ �3��o ����o ����nQ �3��nQ      E  , , ���nQ ���o ����o ����nQ ���nQ      E  , , ����nQ ����o ����o ����nQ ����nQ      E  , , ����nQ ����o ŧ��o ŧ��nQ ����nQ      E  , , ����nQ ����o ȋ��o ȋ��nQ ����nQ      E  , , ʧ��nQ ʧ��o �o��o �o��nQ ʧ��nQ      E  , , ͋��nQ ͋��o �S��o �S��nQ ͋��nQ      E  , , �3��qq �3��r9 ����r9 ����qq �3��qq      E  , , ���qq ���r9 ����r9 ����qq ���qq      E  , , ����qq ����r9 ����r9 ����qq ����qq      E  , , ����qq ����r9 ŧ��r9 ŧ��qq ����qq      E  , , ����qq ����r9 ȋ��r9 ȋ��qq ����qq      E  , , ʧ��qq ʧ��r9 �o��r9 �o��qq ʧ��qq      E  , , ͋��qq ͋��r9 �S��r9 �S��qq ͋��qq      E  , , ����qq ����r9 �k��r9 �k��qq ����qq      E  , , ����qq ����r9 �O��r9 �O��qq ����qq      E  , , �k��qq �k��r9 �3��r9 �3��qq �k��qq      E  , , �O��qq �O��r9 ���r9 ���qq �O��qq      E  , , �3��l� �3��m� ����m� ����l� �3��l�      E  , , ���l� ���m� ����m� ����l� ���l�      E  , , ����l� ����m� ����m� ����l� ����l�      E  , , ����l� ����m� ŧ��m� ŧ��l� ����l�      E  , , ����l� ����m� ȋ��m� ȋ��l� ����l�      E  , , ʧ��l� ʧ��m� �o��m� �o��l� ʧ��l�      E  , , ͋��l� ͋��m� �S��m� �S��l� ͋��l�      E  , , ����qq ����r9 ����r9 ����qq ����qq      E  , , ����qq ����r9 ����r9 ����qq ����qq      E  , , ����l� ����m� ����m� ����l� ����l�      E  , , ����l� ����m� �k��m� �k��l� ����l�      E  , , ����l� ����m� �O��m� �O��l� ����l�      E  , , �k��l� �k��m� �3��m� �3��l� �k��l�      E  , , �O��l� �O��m� ���m� ���l� �O��l�      E  , , ����o� ����p� ����p� ����o� ����o�      E  , , ����o� ����p� ����p� ����o� ����o�      E  , , ����o� ����p� �k��p� �k��o� ����o�      E  , , ����o� ����p� �O��p� �O��o� ����o�      E  , , �k��o� �k��p� �3��p� �3��o� �k��o�      E  , , �O��o� �O��p� ���p� ���o� �O��o�      E  , , �3��o� �3��p� ����p� ����o� �3��o�      E  , , ���o� ���p� ����p� ����o� ���o�      E  , , ����o� ����p� ����p� ����o� ����o�      E  , , ����o� ����p� ŧ��p� ŧ��o� ����o�      E  , , ����o� ����p� ȋ��p� ȋ��o� ����o�      E  , , ����k1 ����k� ����k� ����k1 ����k1      E  , , ����k1 ����k� ����k� ����k1 ����k1      E  , , ����k1 ����k� �k��k� �k��k1 ����k1      E  , , ����k1 ����k� �O��k� �O��k1 ����k1      E  , , �k��k1 �k��k� �3��k� �3��k1 �k��k1      E  , , �O��k1 �O��k� ���k� ���k1 �O��k1      E  , , �3��k1 �3��k� ����k� ����k1 �3��k1      E  , , ���k1 ���k� ����k� ����k1 ���k1      E  , , ����k1 ����k� ����k� ����k1 ����k1      E  , , ����k1 ����k� ŧ��k� ŧ��k1 ����k1      E  , , ����k1 ����k� ȋ��k� ȋ��k1 ����k1      E  , , ʧ��k1 ʧ��k� �o��k� �o��k1 ʧ��k1      E  , , ͋��k1 ͋��k� �S��k� �S��k1 ͋��k1      E  , , ����l� ����m� ����m� ����l� ����l�      E  , , ���nQ ���o ����o ����nQ ���nQ      E  , , ����nQ ����o ����o ����nQ ����nQ      E  , , ����nQ ����o ����o ����nQ ����nQ      E  , , ����o� ����p� �K��p� �K��o� ����o�      E  , , �g��o� �g��p� �/��p� �/��o� �g��o�      E  , , �K��o� �K��p� ���p� ���o� �K��o�      E  , , y���o� y���p� z��p� z��o� y���o�      E  , , |���o� |���p� }c��p� }c��o� |���o�      E  , , ��o� ��p� �G��p� �G��o� ��o�      E  , , �c��o� �c��p� �+��p� �+��o� �c��o�      E  , , �G��o� �G��p� ���p� ���o� �G��o�      E  , , �+��o� �+��p� ����p� ����o� �+��o�      E  , , ����nQ ����o ����o ����nQ ����nQ      E  , , ����nQ ����o �g��o �g��nQ ����nQ      E  , , ����nQ ����o �K��o �K��nQ ����nQ      E  , , �g��nQ �g��o �/��o �/��nQ �g��nQ      E  , , �K��nQ �K��o ���o ���nQ �K��nQ      E  , , �/��nQ �/��o ����o ����nQ �/��nQ      E  , , ���nQ ���o ����o ����nQ ���nQ      E  , , ����nQ ����o ����o ����nQ ����nQ      E  , , �/��qq �/��r9 ����r9 ����qq �/��qq      E  , , ���qq ���r9 ����r9 ����qq ���qq      E  , , ����qq ����r9 ����r9 ����qq ����qq      E  , , ����qq ����r9 ����r9 ����qq ����qq      E  , , ����qq ����r9 ����r9 ����qq ����qq      E  , , ����qq ����r9 ����r9 ����qq ����qq      E  , , ����qq ����r9 �g��r9 �g��qq ����qq      E  , , ����qq ����r9 �K��r9 �K��qq ����qq      E  , , �g��qq �g��r9 �/��r9 �/��qq �g��qq      E  , , �K��qq �K��r9 ���r9 ���qq �K��qq      E  , , �/��o� �/��p� ����p� ����o� �/��o�      E  , , ���o� ���p� ����p� ����o� ���o�      E  , , y���k1 y���k� z��k� z��k1 y���k1      E  , , |���k1 |���k� }c��k� }c��k1 |���k1      E  , , ��k1 ��k� �G��k� �G��k1 ��k1      E  , , �c��k1 �c��k� �+��k� �+��k1 �c��k1      E  , , �G��k1 �G��k� ���k� ���k1 �G��k1      E  , , �+��k1 �+��k� ����k� ����k1 �+��k1      E  , , ���k1 ���k� ����k� ����k1 ���k1      E  , , ����k1 ����k� ����k� ����k1 ����k1      E  , , ����k1 ����k� ����k� ����k1 ����k1      E  , , ����k1 ����k� ����k� ����k1 ����k1      E  , , ����o� ����p� ����p� ����o� ����o�      E  , , ���o� ���p� ����p� ����o� ���o�      E  , , ����o� ����p� ����p� ����o� ����o�      E  , , y���nQ y���o z��o z��nQ y���nQ      E  , , |���nQ |���o }c��o }c��nQ |���nQ      E  , , y���l� y���m� z��m� z��l� y���l�      E  , , |���l� |���m� }c��m� }c��l� |���l�      E  , , ��l� ��m� �G��m� �G��l� ��l�      E  , , �c��l� �c��m� �+��m� �+��l� �c��l�      E  , , �G��l� �G��m� ���m� ���l� �G��l�      E  , , �+��l� �+��m� ����m� ����l� �+��l�      E  , , ���l� ���m� ����m� ����l� ���l�      E  , , ����l� ����m� ����m� ����l� ����l�      E  , , ����l� ����m� ����m� ����l� ����l�      E  , , ����l� ����m� ����m� ����l� ����l�      E  , , ����k1 ����k� �g��k� �g��k1 ����k1      E  , , ����k1 ����k� �K��k� �K��k1 ����k1      E  , , �g��k1 �g��k� �/��k� �/��k1 �g��k1      E  , , �K��k1 �K��k� ���k� ���k1 �K��k1      E  , , �/��k1 �/��k� ����k� ����k1 �/��k1      E  , , ���k1 ���k� ����k� ����k1 ���k1      E  , , ����k1 ����k� ����k� ����k1 ����k1      E  , , ��nQ ��o �G��o �G��nQ ��nQ      E  , , �c��nQ �c��o �+��o �+��nQ �c��nQ      E  , , �G��nQ �G��o ���o ���nQ �G��nQ      E  , , ����o� ����p� ����p� ����o� ����o�      E  , , ����o� ����p� ����p� ����o� ����o�      E  , , ����l� ����m� �g��m� �g��l� ����l�      E  , , ����l� ����m� �K��m� �K��l� ����l�      E  , , �g��l� �g��m� �/��m� �/��l� �g��l�      E  , , �K��l� �K��m� ���m� ���l� �K��l�      E  , , ����o� ����p� �g��p� �g��o� ����o�      E  , , y���qq y���r9 z��r9 z��qq y���qq      E  , , |���qq |���r9 }c��r9 }c��qq |���qq      E  , , ��qq ��r9 �G��r9 �G��qq ��qq      E  , , �c��qq �c��r9 �+��r9 �+��qq �c��qq      E  , , �G��qq �G��r9 ���r9 ���qq �G��qq      E  , , �+��qq �+��r9 ����r9 ����qq �+��qq      E  , , ���qq ���r9 ����r9 ����qq ���qq      E  , , �/��l� �/��m� ����m� ����l� �/��l�      E  , , ���l� ���m� ����m� ����l� ���l�      E  , , ����l� ����m� ����m� ����l� ����l�      E  , , �+��nQ �+��o ����o ����nQ �+��nQ      E  , , ����V_ ����W' ����W' ����V_ ����V_      E  , , ����S? ����T ����T ����S? ����S?      E  , , ����W� ����X� ����X� ����W� ����W�      E  , , ����ca ����d) ����d) ����ca ����ca      E  , , y���[ y���[� z��[� z��[ y���[      E  , , |���[ |���[� }c��[� }c��[ |���[      E  , , ��[ ��[� �G��[� �G��[ ��[      E  , , �c��[ �c��[� �+��[� �+��[ �c��[      E  , , �G��[ �G��[� ���[� ���[ �G��[      E  , , �+��[ �+��[� ����[� ����[ �+��[      E  , , ���[ ���[� ����[� ����[ ���[      E  , , ����[ ����[� ����[� ����[ ����[      E  , , ����[ ����[� ����[� ����[ ����[      E  , , ����[ ����[� ����[� ����[ ����[      E  , , ����[ ����[� �g��[� �g��[ ����[      E  , , ����[ ����[� �K��[� �K��[ ����[      E  , , �g��[ �g��[� �/��[� �/��[ �g��[      E  , , �K��[ �K��[� ���[� ���[ �K��[      E  , , �/��[ �/��[� ����[� ����[ �/��[      E  , , ���[ ���[� ����[� ����[ ���[      E  , , ����[ ����[� ����[� ����[ ����[      E  , , ����Q� ����Rw ����Rw ����Q� ����Q�      E  , , ����P ����P� ����P� ����P ����P      E  , , ����T� ����U� ����U� ����T� ����T�      E  , , ����d� ����e� ����e� ����d� ����d�      E  , , ����N� ����OW ����OW ����N� ����N�      E  , , ����h ����h� ����h� ����h ����h      E  , , ����Y ����ZG ����ZG ����Y ����Y      E  , , ����f� ����gI ����gI ����f� ����f�      E  , , ����L� ����M� ����M� ����L� ����L�      E  , , �g��ca �g��d) �/��d) �/��ca �g��ca      E  , , �K��ca �K��d) ���d) ���ca �K��ca      E  , , �/��ca �/��d) ����d) ����ca �/��ca      E  , , ���ca ���d) ����d) ����ca ���ca      E  , , ����ca ����d) ����d) ����ca ����ca      E  , , ���h ���h� ����h� ����h ���h      E  , , ����h ����h� ����h� ����h ����h      E  , , ����h ����h� �K��h� �K��h ����h      E  , , �g��h �g��h� �/��h� �/��h �g��h      E  , , �K��h �K��h� ���h� ���h �K��h      E  , , �/��h �/��h� ����h� ����h �/��h      E  , , ����f� ����gI ����gI ����f� ����f�      E  , , �g��f� �g��gI �/��gI �/��f� �g��f�      E  , , �K��f� �K��gI ���gI ���f� �K��f�      E  , , ����d� ����e� ����e� ����d� ����d�      E  , , ����d� ����e� �g��e� �g��d� ����d�      E  , , ����d� ����e� �K��e� �K��d� ����d�      E  , , �g��d� �g��e� �/��e� �/��d� �g��d�      E  , , �K��d� �K��e� ���e� ���d� �K��d�      E  , , �/��d� �/��e� ����e� ����d� �/��d�      E  , , ���d� ���e� ����e� ����d� ���d�      E  , , ����d� ����e� ����e� ����d� ����d�      E  , , �/��f� �/��gI ����gI ����f� �/��f�      E  , , ���f� ���gI ����gI ����f� ���f�      E  , , ����h ����h� ����h� ����h ����h      E  , , ����h ����h� �g��h� �g��h ����h      E  , , ����ca ����d) ����d) ����ca ����ca      E  , , ����ca ����d) �g��d) �g��ca ����ca      E  , , ����f� ����gI ����gI ����f� ����f�      E  , , ����f� ����gI �g��gI �g��f� ����f�      E  , , ����f� ����gI �K��gI �K��f� ����f�      E  , , ����ca ����d) �K��d) �K��ca ����ca      E  , , �c��d� �c��e� �+��e� �+��d� �c��d�      E  , , �G��d� �G��e� ���e� ���d� �G��d�      E  , , �+��d� �+��e� ����e� ����d� �+��d�      E  , , ���d� ���e� ����e� ����d� ���d�      E  , , ����d� ����e� ����e� ����d� ����d�      E  , , �c��ca �c��d) �+��d) �+��ca �c��ca      E  , , �G��ca �G��d) ���d) ���ca �G��ca      E  , , �+��ca �+��d) ����d) ����ca �+��ca      E  , , y���ca y���d) z��d) z��ca y���ca      E  , , |���ca |���d) }c��d) }c��ca |���ca      E  , , ��ca ��d) �G��d) �G��ca ��ca      E  , , y���h y���h� z��h� z��h y���h      E  , , |���h |���h� }c��h� }c��h |���h      E  , , ��h ��h� �G��h� �G��h ��h      E  , , �c��h �c��h� �+��h� �+��h �c��h      E  , , y���f� y���gI z��gI z��f� y���f�      E  , , |���f� |���gI }c��gI }c��f� |���f�      E  , , ��f� ��gI �G��gI �G��f� ��f�      E  , , �c��f� �c��gI �+��gI �+��f� �c��f�      E  , , �G��f� �G��gI ���gI ���f� �G��f�      E  , , �+��f� �+��gI ����gI ����f� �+��f�      E  , , ���f� ���gI ����gI ����f� ���f�      E  , , ����f� ����gI ����gI ����f� ����f�      E  , , �G��h �G��h� ���h� ���h �G��h      E  , , �+��h �+��h� ����h� ����h �+��h      E  , , ���h ���h� ����h� ����h ���h      E  , , ����h ����h� ����h� ����h ����h      E  , , y���d� y���e� z��e� z��d� y���d�      E  , , ���ca ���d) ����d) ����ca ���ca      E  , , ����ca ����d) ����d) ����ca ����ca      E  , , |���d� |���e� }c��e� }c��d� |���d�      E  , , ��d� ��e� �G��e� �G��d� ��d�      E  , , �c��P �c��P� �+��P� �+��P �c��P      E  , , �G��P �G��P� ���P� ���P �G��P      E  , , �+��P �+��P� ����P� ����P �+��P      E  , , ���P ���P� ����P� ����P ���P      E  , , ����P ����P� ����P� ����P ����P      E  , , ��S? ��T �G��T �G��S? ��S?      E  , , �+��T� �+��U� ����U� ����T� �+��T�      E  , , ���T� ���U� ����U� ����T� ���T�      E  , , ����T� ����U� ����U� ����T� ����T�      E  , , �c��S? �c��T �+��T �+��S? �c��S?      E  , , |���V_ |���W' }c��W' }c��V_ |���V_      E  , , ��V_ ��W' �G��W' �G��V_ ��V_      E  , , �c��V_ �c��W' �+��W' �+��V_ �c��V_      E  , , �G��V_ �G��W' ���W' ���V_ �G��V_      E  , , �G��S? �G��T ���T ���S? �G��S?      E  , , �+��S? �+��T ����T ����S? �+��S?      E  , , ���S? ���T ����T ����S? ���S?      E  , , ����S? ����T ����T ����S? ����S?      E  , , ���V_ ���W' ����W' ����V_ ���V_      E  , , ���W� ���X� ����X� ����W� ���W�      E  , , ����W� ����X� ����X� ����W� ����W�      E  , , ����V_ ����W' ����W' ����V_ ����V_      E  , , �+��V_ �+��W' ����W' ����V_ �+��V_      E  , , y���Q� y���Rw z��Rw z��Q� y���Q�      E  , , y���W� y���X� z��X� z��W� y���W�      E  , , |���W� |���X� }c��X� }c��W� |���W�      E  , , |���Q� |���Rw }c��Rw }c��Q� |���Q�      E  , , ��Q� ��Rw �G��Rw �G��Q� ��Q�      E  , , �c��Q� �c��Rw �+��Rw �+��Q� �c��Q�      E  , , �G��Q� �G��Rw ���Rw ���Q� �G��Q�      E  , , y���N� y���OW z��OW z��N� y���N�      E  , , |���N� |���OW }c��OW }c��N� |���N�      E  , , ��N� ��OW �G��OW �G��N� ��N�      E  , , �c��N� �c��OW �+��OW �+��N� �c��N�      E  , , �G��N� �G��OW ���OW ���N� �G��N�      E  , , �+��N� �+��OW ����OW ����N� �+��N�      E  , , ���N� ���OW ����OW ����N� ���N�      E  , , ����N� ����OW ����OW ����N� ����N�      E  , , �+��Q� �+��Rw ����Rw ����Q� �+��Q�      E  , , ���Q� ���Rw ����Rw ����Q� ���Q�      E  , , ����Q� ����Rw ����Rw ����Q� ����Q�      E  , , y���S? y���T z��T z��S? y���S?      E  , , |���S? |���T }c��T }c��S? |���S?      E  , , ��W� ��X� �G��X� �G��W� ��W�      E  , , �c��W� �c��X� �+��X� �+��W� �c��W�      E  , , �G��W� �G��X� ���X� ���W� �G��W�      E  , , �+��W� �+��X� ����X� ����W� �+��W�      E  , , y���V_ y���W' z��W' z��V_ y���V_      E  , , y���T� y���U� z��U� z��T� y���T�      E  , , |���T� |���U� }c��U� }c��T� |���T�      E  , , y���Y y���ZG z��ZG z��Y y���Y      E  , , |���Y |���ZG }c��ZG }c��Y |���Y      E  , , ��Y ��ZG �G��ZG �G��Y ��Y      E  , , �c��Y �c��ZG �+��ZG �+��Y �c��Y      E  , , �G��Y �G��ZG ���ZG ���Y �G��Y      E  , , �+��Y �+��ZG ����ZG ����Y �+��Y      E  , , ���Y ���ZG ����ZG ����Y ���Y      E  , , ����Y ����ZG ����ZG ����Y ����Y      E  , , ��T� ��U� �G��U� �G��T� ��T�      E  , , �c��T� �c��U� �+��U� �+��T� �c��T�      E  , , �G��T� �G��U� ���U� ���T� �G��T�      E  , , y���P y���P� z��P� z��P y���P      E  , , |���P |���P� }c��P� }c��P |���P      E  , , y���L� y���M� z��M� z��L� y���L�      E  , , |���L� |���M� }c��M� }c��L� |���L�      E  , , ��L� ��M� �G��M� �G��L� ��L�      E  , , �c��L� �c��M� �+��M� �+��L� �c��L�      E  , , �G��L� �G��M� ���M� ���L� �G��L�      E  , , �+��L� �+��M� ����M� ����L� �+��L�      E  , , ���L� ���M� ����M� ����L� ���L�      E  , , ����L� ����M� ����M� ����L� ����L�      E  , , ��P ��P� �G��P� �G��P ��P      E  , , �/��Q� �/��Rw ����Rw ����Q� �/��Q�      E  , , ���Q� ���Rw ����Rw ����Q� ���Q�      E  , , ����Q� ����Rw ����Rw ����Q� ����Q�      E  , , ����V_ ����W' ����W' ����V_ ����V_      E  , , ����V_ ����W' ����W' ����V_ ����V_      E  , , ����V_ ����W' �g��W' �g��V_ ����V_      E  , , ����V_ ����W' �K��W' �K��V_ ����V_      E  , , ����W� ����X� ����X� ����W� ����W�      E  , , ����W� ����X� �g��X� �g��W� ����W�      E  , , ����W� ����X� �K��X� �K��W� ����W�      E  , , �g��W� �g��X� �/��X� �/��W� �g��W�      E  , , �K��W� �K��X� ���X� ���W� �K��W�      E  , , �/��W� �/��X� ����X� ����W� �/��W�      E  , , ���W� ���X� ����X� ����W� ���W�      E  , , ����P ����P� ����P� ����P ����P      E  , , ����N� ����OW ����OW ����N� ����N�      E  , , ����N� ����OW �g��OW �g��N� ����N�      E  , , ����N� ����OW �K��OW �K��N� ����N�      E  , , �g��N� �g��OW �/��OW �/��N� �g��N�      E  , , �K��N� �K��OW ���OW ���N� �K��N�      E  , , �/��N� �/��OW ����OW ����N� �/��N�      E  , , ���N� ���OW ����OW ����N� ���N�      E  , , ����N� ����OW ����OW ����N� ����N�      E  , , ����P ����P� �g��P� �g��P ����P      E  , , ����P ����P� �K��P� �K��P ����P      E  , , �g��P �g��P� �/��P� �/��P �g��P      E  , , �K��P �K��P� ���P� ���P �K��P      E  , , �/��P �/��P� ����P� ����P �/��P      E  , , ���P ���P� ����P� ����P ���P      E  , , ����P ����P� ����P� ����P ����P      E  , , ����W� ����X� ����X� ����W� ����W�      E  , , ����S? ����T ����T ����S? ����S?      E  , , ����S? ����T �g��T �g��S? ����S?      E  , , ����S? ����T �K��T �K��S? ����S?      E  , , ����T� ����U� ����U� ����T� ����T�      E  , , ����T� ����U� �g��U� �g��T� ����T�      E  , , ����T� ����U� �K��U� �K��T� ����T�      E  , , �g��T� �g��U� �/��U� �/��T� �g��T�      E  , , �K��T� �K��U� ���U� ���T� �K��T�      E  , , �/��T� �/��U� ����U� ����T� �/��T�      E  , , ���T� ���U� ����U� ����T� ���T�      E  , , ����T� ����U� ����U� ����T� ����T�      E  , , �g��S? �g��T �/��T �/��S? �g��S?      E  , , ����Y ����ZG ����ZG ����Y ����Y      E  , , ����Y ����ZG �g��ZG �g��Y ����Y      E  , , ����Y ����ZG �K��ZG �K��Y ����Y      E  , , �g��Y �g��ZG �/��ZG �/��Y �g��Y      E  , , �K��Y �K��ZG ���ZG ���Y �K��Y      E  , , �/��Y �/��ZG ����ZG ����Y �/��Y      E  , , ���Y ���ZG ����ZG ����Y ���Y      E  , , ����Y ����ZG ����ZG ����Y ����Y      E  , , �K��S? �K��T ���T ���S? �K��S?      E  , , �/��S? �/��T ����T ����S? �/��S?      E  , , ���S? ���T ����T ����S? ���S?      E  , , ����S? ����T ����T ����S? ����S?      E  , , �g��V_ �g��W' �/��W' �/��V_ �g��V_      E  , , �K��V_ �K��W' ���W' ���V_ �K��V_      E  , , �/��V_ �/��W' ����W' ����V_ �/��V_      E  , , ���V_ ���W' ����W' ����V_ ���V_      E  , , ����Q� ����Rw ����Rw ����Q� ����Q�      E  , , ����Q� ����Rw �g��Rw �g��Q� ����Q�      E  , , ����Q� ����Rw �K��Rw �K��Q� ����Q�      E  , , �g��Q� �g��Rw �/��Rw �/��Q� �g��Q�      E  , , �K��Q� �K��Rw ���Rw ���Q� �K��Q�      E  , , ����L� ����M� ����M� ����L� ����L�      E  , , ����L� ����M� �g��M� �g��L� ����L�      E  , , ����L� ����M� �K��M� �K��L� ����L�      E  , , �g��L� �g��M� �/��M� �/��L� �g��L�      E  , , �K��L� �K��M� ���M� ���L� �K��L�      E  , , �/��L� �/��M� ����M� ����L� �/��L�      E  , , ���L� ���M� ����M� ����L� ���L�      E  , , ����L� ����M� ����M� ����L� ����L�      E  , , ����[ ����[� ����[� ����[ ����[      E  , , ����[ ����[� ����[� ����[ ����[      E  , , ����[ ����[� �k��[� �k��[ ����[      E  , , ����[ ����[� �O��[� �O��[ ����[      E  , , �k��[ �k��[� �3��[� �3��[ �k��[      E  , , �O��[ �O��[� ���[� ���[ �O��[      E  , , �3��[ �3��[� ����[� ����[ �3��[      E  , , ���[ ���[� ����[� ����[ ���[      E  , , ����[ ����[� ����[� ����[ ����[      E  , , ����[ ����[� ŧ��[� ŧ��[ ����[      E  , , ����[ ����[� ȋ��[� ȋ��[ ����[      E  , , ʧ��[ ʧ��[� �o��[� �o��[ ʧ��[      E  , , ͋��[ ͋��[� �S��[� �S��[ ͋��[      E  , , �T��Z� �T��[� ���[� ���Z� �T��Z�      E  , , ����ca ����d) ŧ��d) ŧ��ca ����ca      E  , , ����]� ����^p ۖ��^p ۖ��]� ����]�      E  , , �T��\Y �T��]! ���]! ���\Y �T��\Y      E  , , ����ca ����d) ȋ��d) ȋ��ca ����ca      E  , , ʧ��ca ʧ��d) �o��d) �o��ca ʧ��ca      E  , , ͋��ca ͋��d) �S��d) �S��ca ͋��ca      E  , , ͋��h ͋��h� �S��h� �S��h ͋��h      E  , , ����bX ����c  ۖ��c  ۖ��bX ����bX      E  , , ����h� ����i` ۖ��i` ۖ��h� ����h�      E  , , ����c� ����d� ۖ��d� ۖ��c� ����c�      E  , , �T��b� �T��ca ���ca ���b� �T��b�      E  , , ʧ��h ʧ��h� �o��h� �o��h ʧ��h      E  , , ����`� ����a� ۖ��a� ۖ��`� ����`�      E  , , �T��_y �T��`A ���`A ���_y �T��_y      E  , , ����\ ����\� ۖ��\� ۖ��\ ����\      E  , , �T��d) �T��d� ���d� ���d) �T��d)      E  , , �T��gI �T��h ���h ���gI �T��gI      E  , , ����_8 ����`  ۖ��`  ۖ��_8 ����_8      E  , , ����f� ����gI ŧ��gI ŧ��f� ����f�      E  , , ����f� ����gI ȋ��gI ȋ��f� ����f�      E  , , ʧ��f� ʧ��gI �o��gI �o��f� ʧ��f�      E  , , ͋��f� ͋��gI �S��gI �S��f� ͋��f�      E  , , ����g ����g� ۖ��g� ۖ��g ����g      E  , , �T��e� �T��f� ���f� ���e� �T��e�      E  , , �T��]� �T��^� ���^� ���]� �T��]�      E  , , ����h ����h� ŧ��h� ŧ��h ����h      E  , , ����h ����h� ȋ��h� ȋ��h ����h      E  , , �T��a	 �T��a� ���a� ���a	 �T��a	      E  , , ����d� ����e� ŧ��e� ŧ��d� ����d�      E  , , ����d� ����e� ȋ��e� ȋ��d� ����d�      E  , , ʧ��d� ʧ��e� �o��e� �o��d� ʧ��d�      E  , , ͋��d� ͋��e� �S��e� �S��d� ͋��d�      E  , , ����ex ����f@ ۖ��f@ ۖ��ex ����ex      E  , , �T��h� �T��i� ���i� ���h� �T��h�      E  , , ����h ����h� �k��h� �k��h ����h      E  , , �k��ca �k��d) �3��d) �3��ca �k��ca      E  , , �O��ca �O��d) ���d) ���ca �O��ca      E  , , �3��ca �3��d) ����d) ����ca �3��ca      E  , , ���ca ���d) ����d) ����ca ���ca      E  , , ����d� ����e� ����e� ����d� ����d�      E  , , ����d� ����e� ����e� ����d� ����d�      E  , , ����f� ����gI ����gI ����f� ����f�      E  , , ����f� ����gI ����gI ����f� ����f�      E  , , ����d� ����e� �k��e� �k��d� ����d�      E  , , ����f� ����gI �k��gI �k��f� ����f�      E  , , ����d� ����e� �O��e� �O��d� ����d�      E  , , ����f� ����gI �O��gI �O��f� ����f�      E  , , �k��f� �k��gI �3��gI �3��f� �k��f�      E  , , �k��d� �k��e� �3��e� �3��d� �k��d�      E  , , �O��d� �O��e� ���e� ���d� �O��d�      E  , , �O��f� �O��gI ���gI ���f� �O��f�      E  , , �3��f� �3��gI ����gI ����f� �3��f�      E  , , ���f� ���gI ����gI ����f� ���f�      E  , , ����f� ����gI ����gI ����f� ����f�      E  , , �3��d� �3��e� ����e� ����d� �3��d�      E  , , ���d� ���e� ����e� ����d� ���d�      E  , , ����d� ����e� ����e� ����d� ����d�      E  , , ����h ����h� �O��h� �O��h ����h      E  , , �k��h �k��h� �3��h� �3��h �k��h      E  , , �O��h �O��h� ���h� ���h �O��h      E  , , �3��h �3��h� ����h� ����h �3��h      E  , , ���h ���h� ����h� ����h ���h      E  , , ����ca ����d) ����d) ����ca ����ca      E  , , ����h ����h� ����h� ����h ����h      E  , , ����h ����h� ����h� ����h ����h      E  , , ����h ����h� ����h� ����h ����h      E  , , ����ca ����d) ����d) ����ca ����ca      E  , , ����ca ����d) ����d) ����ca ����ca      E  , , ����ca ����d) �k��d) �k��ca ����ca      E  , , ����ca ����d) �O��d) �O��ca ����ca      E  , , ����T� ����U� ����U� ����T� ����T�      E  , , ����T� ����U� ����U� ����T� ����T�      E  , , ����T� ����U� �k��U� �k��T� ����T�      E  , , ����T� ����U� �O��U� �O��T� ����T�      E  , , �k��T� �k��U� �3��U� �3��T� �k��T�      E  , , ����W� ����X� ����X� ����W� ����W�      E  , , ����W� ����X� ����X� ����W� ����W�      E  , , ����W� ����X� �k��X� �k��W� ����W�      E  , , ����W� ����X� �O��X� �O��W� ����W�      E  , , ����N� ����OW ����OW ����N� ����N�      E  , , ����N� ����OW ����OW ����N� ����N�      E  , , ����N� ����OW �k��OW �k��N� ����N�      E  , , ����N� ����OW �O��OW �O��N� ����N�      E  , , �k��N� �k��OW �3��OW �3��N� �k��N�      E  , , �O��N� �O��OW ���OW ���N� �O��N�      E  , , �3��N� �3��OW ����OW ����N� �3��N�      E  , , ���N� ���OW ����OW ����N� ���N�      E  , , ����N� ����OW ����OW ����N� ����N�      E  , , �O��T� �O��U� ���U� ���T� �O��T�      E  , , �3��T� �3��U� ����U� ����T� �3��T�      E  , , �k��W� �k��X� �3��X� �3��W� �k��W�      E  , , �O��W� �O��X� ���X� ���W� �O��W�      E  , , ���T� ���U� ����U� ����T� ���T�      E  , , ����T� ����U� ����U� ����T� ����T�      E  , , �O��S? �O��T ���T ���S? �O��S?      E  , , �3��S? �3��T ����T ����S? �3��S?      E  , , ���S? ���T ����T ����S? ���S?      E  , , ����S? ����T ����T ����S? ����S?      E  , , ����S? ����T ����T ����S? ����S?      E  , , ����Q� ����Rw ����Rw ����Q� ����Q�      E  , , ����Q� ����Rw ����Rw ����Q� ����Q�      E  , , ����Q� ����Rw �k��Rw �k��Q� ����Q�      E  , , ����Q� ����Rw �O��Rw �O��Q� ����Q�      E  , , �k��Q� �k��Rw �3��Rw �3��Q� �k��Q�      E  , , �O��Q� �O��Rw ���Rw ���Q� �O��Q�      E  , , �3��Q� �3��Rw ����Rw ����Q� �3��Q�      E  , , ���Q� ���Rw ����Rw ����Q� ���Q�      E  , , ����Q� ����Rw ����Rw ����Q� ����Q�      E  , , ����S? ����T ����T ����S? ����S?      E  , , ����S? ����T �k��T �k��S? ����S?      E  , , ����S? ����T �O��T �O��S? ����S?      E  , , ����P ����P� ����P� ����P ����P      E  , , ����P ����P� ����P� ����P ����P      E  , , ����Y ����ZG ����ZG ����Y ����Y      E  , , ����Y ����ZG ����ZG ����Y ����Y      E  , , ����Y ����ZG �k��ZG �k��Y ����Y      E  , , ����Y ����ZG �O��ZG �O��Y ����Y      E  , , �k��Y �k��ZG �3��ZG �3��Y �k��Y      E  , , �O��Y �O��ZG ���ZG ���Y �O��Y      E  , , �3��Y �3��ZG ����ZG ����Y �3��Y      E  , , ���Y ���ZG ����ZG ����Y ���Y      E  , , ����Y ����ZG ����ZG ����Y ����Y      E  , , ����P ����P� �k��P� �k��P ����P      E  , , ����P ����P� �O��P� �O��P ����P      E  , , �k��P �k��P� �3��P� �3��P �k��P      E  , , �O��P �O��P� ���P� ���P �O��P      E  , , �3��P �3��P� ����P� ����P �3��P      E  , , ���P ���P� ����P� ����P ���P      E  , , ����P ����P� ����P� ����P ����P      E  , , �k��S? �k��T �3��T �3��S? �k��S?      E  , , ����V_ ����W' ����W' ����V_ ����V_      E  , , ����V_ ����W' ����W' ����V_ ����V_      E  , , ����V_ ����W' �k��W' �k��V_ ����V_      E  , , ����V_ ����W' �O��W' �O��V_ ����V_      E  , , �k��V_ �k��W' �3��W' �3��V_ �k��V_      E  , , �O��V_ �O��W' ���W' ���V_ �O��V_      E  , , �3��V_ �3��W' ����W' ����V_ �3��V_      E  , , ���V_ ���W' ����W' ����V_ ���V_      E  , , �3��W� �3��X� ����X� ����W� �3��W�      E  , , ���W� ���X� ����X� ����W� ���W�      E  , , ����W� ����X� ����X� ����W� ����W�      E  , , ����V_ ����W' ����W' ����V_ ����V_      E  , , ����L� ����M� ����M� ����L� ����L�      E  , , ����L� ����M� ����M� ����L� ����L�      E  , , ����L� ����M� �k��M� �k��L� ����L�      E  , , ����L� ����M� �O��M� �O��L� ����L�      E  , , �k��L� �k��M� �3��M� �3��L� �k��L�      E  , , �O��L� �O��M� ���M� ���L� �O��L�      E  , , �3��L� �3��M� ����M� ����L� �3��L�      E  , , ���L� ���M� ����M� ����L� ���L�      E  , , ����L� ����M� ����M� ����L� ����L�      E  , , ����Y ����ZG ȋ��ZG ȋ��Y ����Y      E  , , ʧ��Y ʧ��ZG �o��ZG �o��Y ʧ��Y      E  , , ͋��Y ͋��ZG �S��ZG �S��Y ͋��Y      E  , , ͋��W� ͋��X� �S��X� �S��W� ͋��W�      E  , , ����T� ����U� ŧ��U� ŧ��T� ����T�      E  , , ����T� ����U� ȋ��U� ȋ��T� ����T�      E  , , ʧ��T� ʧ��U� �o��U� �o��T� ʧ��T�      E  , , ͋��T� ͋��U� �S��U� �S��T� ͋��T�      E  , , ����S? ����T ŧ��T ŧ��S? ����S?      E  , , ����P ����P� ŧ��P� ŧ��P ����P      E  , , ����P ����P� ȋ��P� ȋ��P ����P      E  , , ����V_ ����W' ŧ��W' ŧ��V_ ����V_      E  , , ����V_ ����W' ȋ��W' ȋ��V_ ����V_      E  , , ����Q� ����Rw ŧ��Rw ŧ��Q� ����Q�      E  , , ����Q� ����Rw ȋ��Rw ȋ��Q� ����Q�      E  , , ʧ��Q� ʧ��Rw �o��Rw �o��Q� ʧ��Q�      E  , , ͋��Q� ͋��Rw �S��Rw �S��Q� ͋��Q�      E  , , ����N� ����OW ŧ��OW ŧ��N� ����N�      E  , , ����N� ����OW ȋ��OW ȋ��N� ����N�      E  , , ʧ��N� ʧ��OW �o��OW �o��N� ʧ��N�      E  , , ͋��N� ͋��OW �S��OW �S��N� ͋��N�      E  , , ʧ��V_ ʧ��W' �o��W' �o��V_ ʧ��V_      E  , , ����W� ����X� ŧ��X� ŧ��W� ����W�      E  , , ͋��V_ ͋��W' �S��W' �S��V_ ͋��V_      E  , , ʧ��P ʧ��P� �o��P� �o��P ʧ��P      E  , , ͋��P ͋��P� �S��P� �S��P ͋��P      E  , , ����S? ����T ȋ��T ȋ��S? ����S?      E  , , ʧ��S? ʧ��T �o��T �o��S? ʧ��S?      E  , , ͋��S? ͋��T �S��T �S��S? ͋��S?      E  , , ����W� ����X� ȋ��X� ȋ��W� ����W�      E  , , ʧ��W� ʧ��X� �o��X� �o��W� ʧ��W�      E  , , ����Z� ����[P ۖ��[P ۖ��Z� ����Z�      E  , , ����Y ����ZG ŧ��ZG ŧ��Y ����Y      E  , , ����L� ����M� ŧ��M� ŧ��L� ����L�      E  , , ����L� ����M� ȋ��M� ȋ��L� ����L�      E  , , ʧ��L� ʧ��M� �o��M� �o��L� ʧ��L�      E  , , ͋��L� ͋��M� �S��M� �S��L� ͋��L�      E   ,  ;8����  ;8����  T����  T����  ;8����      E   ,  ;8����  ;8����  T����  T����  ;8����      E   ,  (i  $�  (i  (  Y�  (  Y�  $�  (i  $�      E     G���� vin       E     G����3 vcm       E     A#  &m iref      G   , ����� ����@ ����@ ����� �����      G    
����� vout     �     "�     " user_project_wrapper 
  opamp_v1    C�       +D� ��      �   ,             5�  ,�@ 5�  ,�@               	   E   !        +k5 �� +k5 �� +i� ��   	   E   !        +k9 �� +k9 	[   	   E   !        *�� �� *�� 2r   	   E   !        +:  �� +:  �      E   , EJ���@ EJ  	` Gz  	` Gz���@ EJ���@      E   , !v 5�� !v 5�� #� 5�� #� 5�� !v 5��      E   , ]� 5�� ]� 5�� _� 5�� _� 5�� ]� 5��      E   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      E   , � 5�� � 5�� �2 5�� �2 5�� � 5��      E   , B 5�� B 5�� r 5�� r 5�� B 5��      E   , RN 5�� RN 5�� T~ 5�� T~ 5�� RN 5��      E   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      E   ,  �� 5��  �� 5��  �� 5��  �� 5��  �� 5��      E   , "� 5�� "� 5�� "
 5�� "
 5�� "� 5��      E   , #E 5�� #E 5�� #GJ 5�� #GJ 5�� #E 5��      E   , $�Z 5�� $�Z 5�� $�� 5�� $�� 5�� $�Z 5��      E   , %�f 5�� %�f 5�� %�� 5�� %�� 5�� %�f 5��      E   , &�� 5�� &�� 5�� &�� 5�� &�� 5�� &�� 5��      E   , (7� 5�� (7� 5�� (: 5�� (: 5�� (7� 5��      E   , )u� 5�� )u� 5�� )x" 5�� )x" 5�� )u� 5��      E   , *�2 5�� *�2 5�� *�b 5�� *�b 5�� *�2 5��      E   , +�r 5�� +�r 5�� +� 5�� +� 5�� +�r 5��      E   , �6 5�� �6 5�� �f 5�� �f 5�� �6 5��      E   , �. 5�� �. 5�� �^ 5�� �^ 5�� �. 5��      E   , n 5�� n 5�� � 5�� � 5�� n 5��      E   , Tz 5�� Tz 5�� V� 5�� V� 5�� Tz 5��      E   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      E   , �� 5�� �� 5�� �* 5�� �* 5�� �� 5��      E   ,  5��  5�� 6 5�� 6 5��  5��      E   , 	GF 5�� 	GF 5�� 	Iv 5�� 	Iv 5�� 	GF 5��      E   , 
�� 5�� 
�� 5�� 
�� 5�� 
�� 5�� 
�� 5��      E   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      E   , �� 5�� �� 5��   5��   5�� �� 5��      E   , : 5�� : 5�� <B 5�� <B 5�� : 5��      E   , x 5�� x 5�� zN 5�� zN 5�� x 5��      E   , �^ 5�� �^ 5�� �� 5�� �� 5�� �^ 5��      E   , � 5�� � 5�� �� 5�� �� 5�� � 5��      E   , .� 5�� .� 5�� 0� 5�� 0� 5�� .� 5��      E   , j� 5�� j� 5�� m 5�� m 5�� j� 5��      E   , �* 5�� �* 5�� �Z 5�� �Z 5�� �* 5��      E   ,  �� 5��  �� 5��  � 5��  � 5��  �� 5��      E   ,   &���@   &  	`  "V  	`  "V���@   &���@      E   ,  7����@  7�  	`  9�  	`  9����@  7����@      E   ,  N����@  N�  	`  Q  	`  Q���@  N����@      E   ,  f:���@  f:  	`  hj  	`  hj���@  f:���@      E   ,  }����@  }�  	`  �  	`  ����@  }����@      E   ,  �����@  ��  	`  �"  	`  �"���@  �����@      E   ,  �N���@  �N  	`  �~  	`  �~���@  �N���@      E   ,  ê���@  ê  	`  ��  	`  �����@  ê���@      E   ,  ����@  �  	`  �6  	`  �6���@  ����@      E   ,  �b���@  �b  	`  ��  	`  �����@  �b���@      E   , 	����@ 	�  	` �  	` ����@ 	����@      E   , !���@ !  	` #J  	` #J���@ !���@      E   , 8v���@ 8v  	` :�  	` :����@ 8v���@      E   , O����@ O�  	` R  	` R���@ O����@      E   , eb���@ eb  	` g�  	` g����@ eb���@      E   , |����@ |�  	` ~�  	` ~����@ |����@      E   , ����@ �  	` �J  	` �J���@ ����@      E   , �v���@ �v  	` ��  	` �����@ �v���@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �.���@ �.  	` �^  	` �^���@ �.���@      E   , ����@ �  	` �  	` ����@ ����@      E   , ����@ �  	`   	` ���@ ����@      E   ,  B���@  B  	` "r  	` "r���@  B���@      E   , 7����@ 7�  	` 9�  	` 9����@ 7����@      E   , N����@ N�  	` Q*  	` Q*���@ N����@      E   , fV���@ fV  	` h�  	` h����@ fV���@      E   , }����@ }�  	` �  	` ����@ }����@      E   , ����@ �  	` �>  	` �>���@ ����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �*  	` �*���@ �����@      E   , �V���@ �V  	` ۆ  	` ۆ���@ �V���@      E   , ����@ �  	` ��  	` �����@ ����@      E   , ���@   	` 
>  	` 
>���@ ���@      E   , j���@ j  	` !�  	` !����@ j���@      E   , 6����@ 6�  	` 8�  	` 8����@ 6����@      E   , N"���@ N"  	` PR  	` PR���@ N"���@      E   , e~���@ e~  	` g�  	` g����@ e~���@      E   , |����@ |�  	` 
  	` 
���@ |����@      E   , �6���@ �6  	` �f  	` �f���@ �6���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �J���@ �J  	` �z  	` �z���@ �J���@      E   , �����@ ��  	` �
  	` �
���@ �����@      E   , 6���@ 6  	` 	f  	` 	f���@ 6���@      E   , ����@ �  	`  �  	`  ����@ ����@      E   , 5����@ 5�  	` 8  	` 8���@ 5����@      E   , MJ���@ MJ  	` Oz  	` Oz���@ MJ���@      E   , d����@ d�  	` f�  	` f����@ d����@      E   , |���@ |  	` ~2  	` ~2���@ |���@      E   , �^���@ �^  	` ��  	` �����@ �^���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �F  	` �F���@ ����@      E   , �r���@ �r  	` ۢ  	` ۢ���@ �r���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , *���@ *  	` 
Z  	` 
Z���@ *���@      E   , ����@ �  	` !�  	` !����@ ����@      E   , 5���@ 5  	` 7F  	` 7F���@ 5���@      E   , Lr���@ Lr  	` N�  	` N����@ Lr���@      E   , c����@ c�  	` e�  	` e����@ c����@      E   , {*���@ {*  	` }Z  	` }Z���@ {*���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   ,  
����@  
�  	`  �  	`  ����@  
����@      E   , �>���@ �>  	` �n  	` �n���@ �>���@      E   , ؚ���@ ؚ  	` ��  	` �����@ ؚ���@      E   , �����@ ��  	` �&  	` �&���@ �����@      E   , R���@ R  	` 	�  	` 	����@ R���@      E   , ����@ �  	`  �  	`  ����@ ����@      E   , 6
���@ 6
  	` 8:  	` 8:���@ 6
���@      E   , Mf���@ Mf  	` O�  	` O����@ Mf���@      E   , d����@ d�  	` f�  	` f����@ d����@      E   , zR���@ zR  	` |�  	` |����@ zR���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �
���@ �
  	` �:  	` �:���@ �
���@      E   , �f���@ �f  	`   	` ���@ �f���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �N  	` �N���@ ����@      E   , z���@ z  	` �  	` ����@ z���@      E   , ����@ �  	`    	`  ���@ ����@      E   , 52���@ 52  	` 7b  	` 7b���@ 52���@      E   , L����@ L�  	` N�  	` N����@ L����@      E   , c����@ c�  	` f  	` f���@ c����@      E   , {F���@ {F  	` }v  	` }v���@ {F���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �.  	` �.���@ �����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �F���@ �F  	` �v  	` �v���@ �F���@      E   , ����@ �  	` �  	` ����@ ����@      E   , ����@ �  	` .  	` .���@ ����@      E   , 4Z���@ 4Z  	` 6�  	` 6����@ 4Z���@      E   , K����@ K�  	` M�  	` M����@ K����@      E   , c���@ c  	` eB  	` eB���@ c���@      E   , zn���@ zn  	` |�  	` |����@ zn���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �&���@ �&  	` �V  	` �V���@ �&���@      E   , �����@ ��  	` ²  	` ²���@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �:���@ �:  	` �j  	` �j���@ �:���@      E   , 	����@ 	�  	` 	�  	` 	����@ 	����@      E   , 	&���@ 	&  	` 	V  	` 	V���@ 	&���@      E   , 	3����@ 	3�  	` 	5�  	` 	5����@ 	3����@      E   , 	J����@ 	J�  	` 	M  	` 	M���@ 	J����@      E   , 	b:���@ 	b:  	` 	dj  	` 	dj���@ 	b:���@      E   , 	y����@ 	y�  	` 	{�  	` 	{����@ 	y����@      E   , 	�����@ 	��  	` 	�"  	` 	�"���@ 	�����@      E   , 	�N���@ 	�N  	` 	�~  	` 	�~���@ 	�N���@      E   , 	�����@ 	��  	` 	��  	` 	�����@ 	�����@      E   , 	����@ 	�  	` 	�6  	` 	�6���@ 	����@      E   , 	�b���@ 	�b  	` 	�  	` 	����@ 	�b���@      E   , 
����@ 
�  	` 
�  	` 
����@ 
����@      E   , 
���@ 
  	` 
J  	` 
J���@ 
���@      E   , 
4v���@ 
4v  	` 
6�  	` 
6����@ 
4v���@      E   , 
J���@ 
J  	` 
L6  	` 
L6���@ 
J���@      E   , 
ab���@ 
ab  	` 
c�  	` 
c����@ 
ab���@      E   , 
x����@ 
x�  	` 
z�  	` 
z����@ 
x����@      E   , 
����@ 
�  	` 
�J  	` 
�J���@ 
����@      E   , 
�v���@ 
�v  	` 
��  	` 
�����@ 
�v���@      E   , 
�����@ 
��  	` 
�  	` 
����@ 
�����@      E   , 
�.���@ 
�.  	` 
�^  	` 
�^���@ 
�.���@      E   , 
����@ 
�  	` 
�  	` 
����@ 
����@      E   , ����@ �  	`   	` ���@ ����@      E   , B���@ B  	` r  	` r���@ B���@      E   , �����@ ��  	` �  	` ����@ �����@      E   , J����@ J�  	` M*  	` M*���@ J����@      E   , bV���@ bV  	` d�  	` d����@ bV���@      E   , y����@ y�  	` {�  	` {����@ y����@      E   , �B���@ �B  	` �r  	` �r���@ �B���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �*  	` �*���@ �����@      E   , �V���@ �V  	` ׆  	` ׆���@ �V���@      E   , ����@ �  	` ��  	` �����@ ����@      E   , ���@   	` >  	` >���@ ���@      E   , j���@ j  	` �  	` ����@ j���@      E   , 2����@ 2�  	` 4�  	` 4����@ 2����@      E   , J"���@ J"  	` LR  	` LR���@ J"���@      E   , a~���@ a~  	` c�  	` c����@ a~���@      E   , x����@ x�  	` {
  	` {
���@ x����@      E   , �6���@ �6  	` �f  	` �f���@ �6���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �~���@ �~  	` ֮  	` ֮���@ �~���@      E   , �����@ ��  	` �
  	` �
���@ �����@      E   , 6���@ 6  	` f  	` f���@ 6���@      E   , ����@ �  	` �  	` ����@ ����@      E   , 1����@ 1�  	` 4  	` 4���@ 1����@      E   , IJ���@ IJ  	` Kz  	` Kz���@ IJ���@      E   , `����@ `�  	` b�  	` b����@ `����@      E   , x���@ x  	` z2  	` z2���@ x���@      E   , �^���@ �^  	` ��  	` �����@ �^���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �F  	` �F���@ ����@      E   , �r���@ �r  	` ע  	` ע���@ �r���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , *���@ *  	` Z  	` Z���@ *���@      E   , ����@ �  	` �  	` ����@ ����@      E   , 1���@ 1  	` 3F  	` 3F���@ 1���@      E   , Hr���@ Hr  	` J�  	` J����@ Hr���@      E   , _����@ _�  	` a�  	` a����@ _����@      E   , w*���@ w*  	` yZ  	` yZ���@ w*���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �>���@ �>  	` �n  	` �n���@ �>���@      E   , Ԛ���@ Ԛ  	` ��  	` �����@ Ԛ���@      E   , �����@ ��  	` �&  	` �&���@ �����@      E   , R���@ R  	` �  	` ����@ R���@      E   , ����@ �  	` �  	` ����@ ����@      E   , 2
���@ 2
  	` 4:  	` 4:���@ 2
���@      E   , If���@ If  	` K�  	` K����@ If���@      E   , ^����@ ^�  	` a&  	` a&���@ ^����@      E   , vR���@ vR  	` x�  	` x����@ vR���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �
���@ �
  	` �:  	` �:���@ �
���@      E   , �f���@ �f  	` ��  	` �����@ �f���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �N  	` �N���@ ����@      E   , z���@ z  	` �  	` ����@ z���@      E   , ����@ �  	`   	` ���@ ����@      E   , 12���@ 12  	` 3b  	` 3b���@ 12���@      E   , H����@ H�  	` J�  	` J����@ H����@      E   , _����@ _�  	` b  	` b���@ _����@      E   , wF���@ wF  	` yv  	` yv���@ wF���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �2���@ �2  	` �b  	` �b���@ �2���@      E   , 3����@ 3�  	` 5�  	` 5����@ 3����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �F���@ �F  	` �v  	` �v���@ �F���@      E   , ����@ �  	` �  	` ����@ ����@      E   , ����@ �  	` .  	` .���@ ����@      E   , 0Z���@ 0Z  	` 2�  	` 2����@ 0Z���@      E   , G����@ G�  	` I�  	` I����@ G����@      E   , _���@ _  	` aB  	` aB���@ _���@      E   , vn���@ vn  	` x�  	` x����@ vn���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �&���@ �&  	` �V  	` �V���@ �&���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �n���@ �n  	` �  	` ����@ �n���@      E   ,  ����@  �  	` �  	` ����@  ����@      E   , &���@ &  	` V  	` V���@ &���@      E   , /����@ /�  	` 1�  	` 1����@ /����@      E   , F����@ F�  	` I  	` I���@ F����@      E   , ^:���@ ^:  	` `j  	` `j���@ ^:���@      E   , u����@ u�  	` w�  	` w����@ u����@      E   , �����@ ��  	` �"  	` �"���@ �����@      E   , �N���@ �N  	` �~  	` �~���@ �N���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �6  	` �6���@ ����@      E   , �b���@ �b  	` �  	` ����@ �b���@      E   , ����@ �  	` �  	` ����@ ����@      E   , ���@   	` J  	` J���@ ���@      E   , .����@ .�  	` 0�  	` 0����@ .����@      E   , F���@ F  	` H6  	` H6���@ F���@      E   , ]b���@ ]b  	` _�  	` _����@ ]b���@      E   , t����@ t�  	` v�  	` v����@ t����@      E   , ����@ �  	` �J  	` �J���@ ����@      E   , �v���@ �v  	` ��  	` �����@ �v���@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �.���@ �.  	` �^  	` �^���@ �.���@      E   , ����@ �  	` �  	` ����@ ����@      E   ,  ����@  �  	`   	` ���@  ����@      E   , B���@ B  	` r  	` r���@ B���@      E   , /����@ /�  	` 1�  	` 1����@ /����@      E   , F����@ F�  	` I*  	` I*���@ F����@      E   , ^V���@ ^V  	` `�  	` `����@ ^V���@      E   , s����@ s�  	` v  	` v���@ s����@      E   , �B���@ �B  	` �r  	` �r���@ �B���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �*  	` �*���@ �����@      E   , �V���@ �V  	` ӆ  	` ӆ���@ �V���@      E   , ����@ �  	` ��  	` �����@ ����@      E   ,  ���@    	` >  	` >���@  ���@      E   , j���@ j  	` �  	` ����@ j���@      E   , .����@ .�  	` 0�  	` 0����@ .����@      E   , F"���@ F"  	` HR  	` HR���@ F"���@      E   , ]~���@ ]~  	` _�  	` _����@ ]~���@      E   , t����@ t�  	` w
  	` w
���@ t����@      E   , �6���@ �6  	` �f  	` �f���@ �6���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �"���@ �"  	` �R  	` �R���@ �"���@      E   , �~���@ �~  	` Ү  	` Ү���@ �~���@      E   , �����@ ��  	` �
  	` �
���@ �����@      E   , �6���@ �6  	` f  	` f���@ �6���@      E   , ����@ �  	` �  	` ����@ ����@      E   , -����@ -�  	` 0  	` 0���@ -����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , \����@ \�  	` ^�  	` ^����@ \����@      E   , t���@ t  	` v2  	` v2���@ t���@      E   , �^���@ �^  	` ��  	` �����@ �^���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �F  	` �F���@ ����@      E   , �r���@ �r  	` Ӣ  	` Ӣ���@ �r���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �^���@ �^  	`  �  	`  ����@ �^���@      E   , ����@ �  	` �  	` ����@ ����@      E   , -���@ -  	` /F  	` /F���@ -���@      E   , Dr���@ Dr  	` F�  	` F����@ Dr���@      E   , [����@ [�  	` ]�  	` ]����@ [����@      E   , s*���@ s*  	` uZ  	` uZ���@ s*���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �>���@ �>  	` �n  	` �n���@ �>���@      E   , К���@ К  	` ��  	` �����@ К���@      E   , �����@ ��  	` �&  	` �&���@ �����@      E   , �R���@ �R  	` �  	` ����@ �R���@      E   , ����@ �  	` �  	` ����@ ����@      E   , .
���@ .
  	` 0:  	` 0:���@ .
���@      E   , C����@ C�  	` E�  	` E����@ C����@      E   , Z����@ Z�  	` ]&  	` ]&���@ Z����@      E   , rR���@ rR  	` t�  	` t����@ rR���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �
���@ �
  	` �:  	` �:���@ �
���@      E   , �f���@ �f  	` ��  	` �����@ �f���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �N  	` �N���@ ����@      E   , �z���@ �z  	`  �  	`  ����@ �z���@      E   , ����@ �  	`   	` ���@ ����@      E   , -2���@ -2  	` /b  	` /b���@ -2���@      E   , D����@ D�  	` F�  	` F����@ D����@      E   , [����@ [�  	` ^  	` ^���@ [����@      E   , sF���@ sF  	` uv  	` uv���@ sF���@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �2���@ �2  	` �b  	` �b���@ �2���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �F���@ �F  	` �v  	` �v���@ �F���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` .  	` .���@ ����@      E   , ,Z���@ ,Z  	` .�  	` .����@ ,Z���@      E   , C����@ C�  	` E�  	` E����@ C����@      E   , [���@ [  	` ]B  	` ]B���@ [���@      E   , rn���@ rn  	` t�  	` t����@ rn���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �&���@ �&  	` �V  	` �V���@ �&���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �B  	` �B���@ ����@      E   , �n���@ �n  	` �  	` ����@ �n���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , &���@ &  	` V  	` V���@ &���@      E   , +����@ +�  	` -�  	` -����@ +����@      E   , B����@ B�  	` E  	` E���@ B����@      E   , Z:���@ Z:  	` \j  	` \j���@ Z:���@      E   , q����@ q�  	` s�  	` s����@ q����@      E   , �����@ ��  	` �"  	` �"���@ �����@      E   , �N���@ �N  	` �~  	` �~���@ �N���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �6  	` �6���@ ����@      E   , �b���@ �b  	` �  	` ����@ �b���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , N���@ N  	` ~  	` ~���@ N���@      E   , *����@ *�  	` ,�  	` ,����@ *����@      E   , B���@ B  	` D6  	` D6���@ B���@      E   , Yb���@ Yb  	` [�  	` [����@ Yb���@      E   , p����@ p�  	` r�  	` r����@ p����@      E   , ����@ �  	` �J  	` �J���@ ����@      E   , �v���@ �v  	` ��  	` �����@ �v���@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �.���@ �.  	` �^  	` �^���@ �.���@      E   , ����@ �  	` �  	` ����@ ����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , B���@ B  	` r  	` r���@ B���@      E   , +����@ +�  	` -�  	` -����@ +����@      E   , B����@ B�  	` E*  	` E*���@ B����@      E   , X����@ X�  	` Z�  	` Z����@ X����@      E   , o����@ o�  	` r  	` r���@ o����@      E   , �B���@ �B  	` �r  	` �r���@ �B���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �*  	` �*���@ �����@      E   , �V���@ �V  	` φ  	` φ���@ �V���@      E   , ����@ �  	` ��  	` �����@ ����@      E   , ����@ �  	` �>  	` �>���@ ����@      E   , j���@ j  	` �  	` ����@ j���@      E   , *����@ *�  	` ,�  	` ,����@ *����@      E   , B"���@ B"  	` DR  	` DR���@ B"���@      E   , Y~���@ Y~  	` [�  	` [����@ Y~���@      E   , p����@ p�  	` s
  	` s
���@ p����@      E   , �6���@ �6  	` �f  	` �f���@ �6���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �"���@ �"  	` �R  	` �R���@ �"���@      E   , �~���@ �~  	` ή  	` ή���@ �~���@      E   , �����@ ��  	` �
  	` �
���@ �����@      E   , �6���@ �6  	` �f  	` �f���@ �6���@      E   , ����@ �  	` �  	` ����@ ����@      E   , )����@ )�  	` ,  	` ,���@ )����@      E   , AJ���@ AJ  	` Cz  	` Cz���@ AJ���@      E   , X����@ X�  	` Z�  	` Z����@ X����@      E   , p���@ p  	` r2  	` r2���@ p���@      E   , �^���@ �^  	` ��  	` �����@ �^���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �F  	` �F���@ ����@      E   , �r���@ �r  	` Ϣ  	` Ϣ���@ �r���@      E   , ����@ �  	` �2  	` �2���@ ����@      E   , �^���@ �^  	` ��  	` �����@ �^���@      E   ,  ����@  �  	`  �  	`  ����@  ����@      E   ,  )���@  )  	`  +F  	`  +F���@  )���@      E   ,  @r���@  @r  	`  B�  	`  B����@  @r���@      E   ,  W����@  W�  	`  Y�  	`  Y����@  W����@      E   ,  o*���@  o*  	`  qZ  	`  qZ���@  o*���@      E   ,  �����@  ��  	`  ��  	`  �����@  �����@      E   ,  �����@  ��  	`  �  	`  ����@  �����@      E   ,  �>���@  �>  	`  �n  	`  �n���@  �>���@      E   ,  ̚���@  ̚  	`  ��  	`  �����@  ̚���@      E   ,  �����@  ��  	`  �&  	`  �&���@  �����@      E   ,  �R���@  �R  	`  ��  	`  �����@  �R���@      E   , !����@ !�  	` !�  	` !����@ !����@      E   , !(>���@ !(>  	` !*n  	` !*n���@ !(>���@      E   , !?����@ !?�  	` !A�  	` !A����@ !?����@      E   , !V����@ !V�  	` !Y&  	` !Y&���@ !V����@      E   , !nR���@ !nR  	` !p�  	` !p����@ !nR���@      E   , !�����@ !��  	` !��  	` !�����@ !�����@      E   , !�
���@ !�
  	` !�:  	` !�:���@ !�
���@      E   , !�f���@ !�f  	` !��  	` !�����@ !�f���@      E   , !�����@ !��  	` !��  	` !�����@ !�����@      E   , !����@ !�  	` !�N  	` !�N���@ !����@      E   , !�z���@ !�z  	` !��  	` !�����@ !�z���@      E   , "����@ "�  	` "  	` "���@ "����@      E   , ")2���@ ")2  	` "+b  	` "+b���@ ")2���@      E   , "@����@ "@�  	` "B�  	` "B����@ "@����@      E   , "W����@ "W�  	` "Z  	` "Z���@ "W����@      E   , "mz���@ "mz  	` "o�  	` "o����@ "mz���@      E   , "�����@ "��  	` "�  	` "����@ "�����@      E   , "�2���@ "�2  	` "�b  	` "�b���@ "�2���@      E   , "�����@ "��  	` "��  	` "�����@ "�����@      E   , "�����@ "��  	` "�  	` "����@ "�����@      E   , "�F���@ "�F  	` "�v  	` "�v���@ "�F���@      E   , "�����@ "��  	` "��  	` "�����@ "�����@      E   , #����@ #�  	` #.  	` #.���@ #����@      E   , #(Z���@ #(Z  	` #*�  	` #*����@ #(Z���@      E   , #?����@ #?�  	` #A�  	` #A����@ #?����@      E   , #W���@ #W  	` #YB  	` #YB���@ #W���@      E   , #nn���@ #nn  	` #p�  	` #p����@ #nn���@      E   , #�����@ #��  	` #��  	` #�����@ #�����@      E   , #�&���@ #�&  	` #�V  	` #�V���@ #�&���@      E   , #�����@ #��  	` #��  	` #�����@ #�����@      E   , #����@ #�  	` #�B  	` #�B���@ #����@      E   , #�n���@ #�n  	` #�  	` #����@ #�n���@      E   , #�����@ #��  	` #��  	` #�����@ #�����@      E   , $&���@ $&  	` $V  	` $V���@ $&���@      E   , $'����@ $'�  	` $)�  	` $)����@ $'����@      E   , $>����@ $>�  	` $A  	` $A���@ $>����@      E   , $V:���@ $V:  	` $Xj  	` $Xj���@ $V:���@      E   , $m����@ $m�  	` $o�  	` $o����@ $m����@      E   , $�����@ $��  	` $�"  	` $�"���@ $�����@      E   , $�N���@ $�N  	` $�~  	` $�~���@ $�N���@      E   , $�����@ $��  	` $��  	` $�����@ $�����@      E   , $����@ $�  	` $�6  	` $�6���@ $����@      E   , $�b���@ $�b  	` $�  	` $����@ $�b���@      E   , $�����@ $��  	` $�"  	` $�"���@ $�����@      E   , %N���@ %N  	` %~  	` %~���@ %N���@      E   , %&����@ %&�  	` %(�  	` %(����@ %&����@      E   , %>���@ %>  	` %@6  	` %@6���@ %>���@      E   , %Ub���@ %Ub  	` %W�  	` %W����@ %Ub���@      E   , %l����@ %l�  	` %n�  	` %n����@ %l����@      E   , %����@ %�  	` %�J  	` %�J���@ %����@      E   , %�v���@ %�v  	` %��  	` %�����@ %�v���@      E   , %�����@ %��  	` %�  	` %����@ %�����@      E   , %�.���@ %�.  	` %�^  	` %�^���@ %�.���@      E   , %����@ %�  	` %�  	` %����@ %����@      E   , %�����@ %��  	` %�  	` %����@ %�����@      E   , &B���@ &B  	` &r  	` &r���@ &B���@      E   , &'����@ &'�  	` &)�  	` &)����@ &'����@      E   , &=.���@ &=.  	` &?^  	` &?^���@ &=.���@      E   , &T����@ &T�  	` &V�  	` &V����@ &T����@      E   , &k����@ &k�  	` &n  	` &n���@ &k����@      E   , &�B���@ &�B  	` &�r  	` &�r���@ &�B���@      E   , &�����@ &��  	` &��  	` &�����@ &�����@      E   , &�����@ &��  	` &�*  	` &�*���@ &�����@      E   , &�V���@ &�V  	` &ˆ  	` &ˆ���@ &�V���@      E   , &����@ &�  	` &��  	` &�����@ &����@      E   , &����@ &�  	` &�>  	` &�>���@ &����@      E   , 'j���@ 'j  	` '�  	` '����@ 'j���@      E   , '&����@ '&�  	` '(�  	` '(����@ '&����@      E   , '>"���@ '>"  	` '@R  	` '@R���@ '>"���@      E   , 'U~���@ 'U~  	` 'W�  	` 'W����@ 'U~���@      E   , 'l����@ 'l�  	` 'o
  	` 'o
���@ 'l����@      E   , '�j���@ '�j  	` '��  	` '�����@ '�j���@      E   , '�����@ '��  	` '��  	` '�����@ '�����@      E   , '�"���@ '�"  	` '�R  	` '�R���@ '�"���@      E   , '�~���@ '�~  	` 'ʮ  	` 'ʮ���@ '�~���@      E   , '�����@ '��  	` '�
  	` '�
���@ '�����@      E   , '�6���@ '�6  	` '�f  	` '�f���@ '�6���@      E   , (����@ (�  	` (�  	` (����@ (����@      E   , (%����@ (%�  	` ((  	` ((���@ (%����@      E   , (=J���@ (=J  	` (?z  	` (?z���@ (=J���@      E   , (T����@ (T�  	` (V�  	` (V����@ (T����@      E   , (l���@ (l  	` (n2  	` (n2���@ (l���@      E   , (�^���@ (�^  	` (��  	` (�����@ (�^���@      E   , (�����@ (��  	` (��  	` (�����@ (�����@      E   , (����@ (�  	` (�F  	` (�F���@ (����@      E   , (Ǧ���@ (Ǧ  	` (��  	` (�����@ (Ǧ���@      E   , (����@ (�  	` (�2  	` (�2���@ (����@      E   , (�^���@ (�^  	` (��  	` (�����@ (�^���@      E   , )����@ )�  	` )�  	` )����@ )����@      E   , )%���@ )%  	` )'F  	` )'F���@ )%���@      E   , )<r���@ )<r  	` )>�  	` )>����@ )<r���@      E   , )S����@ )S�  	` )U�  	` )U����@ )S����@      E   , )k*���@ )k*  	` )mZ  	` )mZ���@ )k*���@      E   , )�����@ )��  	` )��  	` )�����@ )�����@      E   , )�����@ )��  	` )�  	` )����@ )�����@      E   , )�>���@ )�>  	` )�n  	` )�n���@ )�>���@      E   , )Ț���@ )Ț  	` )��  	` )�����@ )Ț���@      E   , )�����@ )��  	` )�&  	` )�&���@ )�����@      E   , )�R���@ )�R  	` )��  	` )�����@ )�R���@      E   , *����@ *�  	` *  	` *���@ *����@      E   , *$>���@ *$>  	` *&n  	` *&n���@ *$>���@      E   , *;����@ *;�  	` *=�  	` *=����@ *;����@      E   , *R����@ *R�  	` *U&  	` *U&���@ *R����@      E   , *jR���@ *jR  	` *l�  	` *l����@ *jR���@      E   , *�����@ *��  	` *��  	` *�����@ *�����@      E   , *�
���@ *�
  	` *�:  	` *�:���@ *�
���@      E   , *�f���@ *�f  	` *��  	` *�����@ *�f���@      E   , *�����@ *��  	` *��  	` *�����@ *�����@      E   , *����@ *�  	` *�N  	` *�N���@ *����@      E   , *�z���@ *�z  	` *��  	` *�����@ *�z���@      E   , +����@ +�  	` +  	` +���@ +����@      E   , +%2���@ +%2  	` +'b  	` +'b���@ +%2���@      E   , +<����@ +<�  	` +>�  	` +>����@ +<����@      E   , +R���@ +R  	` +TN  	` +TN���@ +R���@      E   , +iz���@ +iz  	` +k�  	` +k����@ +iz���@      E   , +�����@ +��  	` +�  	` +����@ +�����@      E   , +�2���@ +�2  	` +�b  	` +�b���@ +�2���@      E   , +�����@ +��  	` +��  	` +�����@ +�����@      E   , +�����@ +��  	` +�  	` +����@ +�����@      E   , +�F���@ +�F  	` +�v  	` +�v���@ +�F���@      E   , +�����@ +��  	` +��  	` +�����@ +�����@      E   , ,����@ ,�  	` ,.  	` ,.���@ ,����@      E   , ,$Z���@ ,$Z  	` ,&�  	` ,&����@ ,$Z���@      E   , ,;����@ ,;�  	` ,=�  	` ,=����@ ,;����@      E   , ,S���@ ,S  	` ,UB  	` ,UB���@ ,S���@      E   , ,jn���@ ,jn  	` ,l�  	` ,l����@ ,jn���@      E   , ,�����@ ,��  	` ,��  	` ,�����@ ,�����@   	   F   !        ,�  s� +�  s�   	   F   !        ,� � +i� �   	   F   !        ,�� �� +8r ��   	   F   !        ,�� 0� *�< 0�      F   ,���@ ִ���@ �d  	` �d  	` ִ���@ ִ      F   , ,�� 4Zl ,�� 4_ ,�  4_ ,�  4Zl ,�� 4Zl      F   , ,�� 3u� ,�� 3z� ,�  3z� ,�  3u� ,�� 3u�      F   , ,�� 2�� ,�� 2�� ,�  2�� ,�  2�� ,�� 2��      F   , ,�� 1�t ,�� 1�$ ,�  1�$ ,�  1�t ,�� 1�t      F   , ,�� 0� ,�� 0ʴ ,�  0ʴ ,�  0� ,�� 0�      F   , ,�� /� ,�� /�D ,�  /�D ,�  /� ,�� /�      F   , ,�� .�| ,�� .�, ,�  .�, ,�  .�| ,�� .�|      F   , ,�� . ,�� .� ,�  .� ,�  . ,�� .      F   , ,�� -1� ,�� -6L ,�  -6L ,�  -1� ,�� -1�      F   , ,�� ,M, ,�� ,Q� ,�  ,Q� ,�  ,M, ,�� ,M,      F   , ,�� +f ,�� +j� ,�  +j� ,�  +f ,�� +f      F   , ,�� *�� ,�� *�T ,�  *�T ,�  *�� ,�� *��      F   , ,�� )�4 ,�� )�� ,�  )�� ,�  )�4 ,�� )�4      F   , ,�� (�� ,�� (�t ,�  (�t ,�  (�� ,�� (��      F   , ,�� 'Ѭ ,�� '�\ ,�  '�\ ,�  'Ѭ ,�� 'Ѭ      F   , ,�� &�< ,�� &�� ,�  &�� ,�  &�< ,�� &�<      F   , ,�� &� ,�� &| ,�  &| ,�  &� ,�� &�      F   , ,�� %!� ,�� %&d ,�  %&d ,�  %!� ,�� %!�      F   , ,�� $=D ,�� $A� ,�  $A� ,�  $=D ,�� $=D      F   , ,�� #X� ,�� #]� ,�  #]� ,�  #X� ,�� #X�      F   , ,�� "td ,�� "y ,�  "y ,�  "td ,�� "td      F   , ,�� !�L ,�� !�� ,�  !�� ,�  !�L ,�� !�L      F   , ,��  �� ,��  �� ,�   �� ,�   �� ,��  ��      F   , ,�� �l ,�� � ,�  � ,�  �l ,�� �l      F   , ,�� �� ,�� � ,�  � ,�  �� ,�� ��      F   , ,�� �� ,�� �� ,�  �� ,�  �� ,�� ��      F   , ,�� t ,�� $ ,�  $ ,�  t ,�� t      F   , ,�� 0 ,�� 4� ,�  4� ,�  0 ,�� 0      F   , ,�� K� ,�� PD ,�  PD ,�  K� ,�� K�      F   , ,�� 5>� ,�� 5C� ,�  5C� ,�  5>� ,�� 5>�      F   ,���@ 2�����@ 2��  	` 2��  	` 2�����@ 2��      F   ,���@ %˴���@ %�d  	` %�d  	` %˴���@ %˴      F   ,���@ ,_����@ ,dt  	` ,dt  	` ,_����@ ,_�      F   ,���@ $�$���@ $��  	` $��  	` $�$���@ $�$      F   ,���@ 0�����@ 0�d  	` 0�d  	` 0�����@ 0��      F   ,���@ #�<���@ #��  	` #��  	` #�<���@ #�<      F   ,���@ 4
����@ 4l  	` 4l  	` 4
����@ 4
�      F   ,���@ "�����@ "�\  	` "�\  	` "�����@ "��      F   ,���@ +F4���@ +J�  	` +J�  	` +F4���@ +F4      F   ,���@ /�����@ /�|  	` /�|  	` /�����@ /��      F   ,���@ !h���@ !l�  	` !l�  	` !h���@ !h      F   ,���@ */L���@ *3�  	` *3�  	` */L���@ */L      F   ,���@  Q4���@  U�  	`  U�  	`  Q4���@  Q4      F   ,���@ 1�D���@ 1��  	` 1��  	` 1�D���@ 1�D      F   ,���@ 7����@ <T  	` <T  	` 7����@ 7�      F   ,���@ )����@ )l  	` )l  	` )����@ )�      F   ,���@  ����@ %l  	` %l  	`  ����@  �      F   ,���@ .�<���@ .��  	` .��  	` .�<���@ .�<      F   ,���@ '�,���@ ( �  	` ( �  	` '�,���@ '�,      F   ,���@ ,���@ �  	` �  	` ,���@ ,      F   ,���@ 5$L���@ 5(�  	` 5(�  	` 5$L���@ 5$L      F   ,���@ ����@ �L  	` �L  	` ����@ �      F   ,���@ -v����@ -{\  	` -{\  	` -v����@ -v�      F   ,���@ &�D���@ &��  	` &��  	` &�D���@ &�D      F   ,���@ �$���@ ��  	` ��  	` �$���@ �$      F   ,���@ �����@ �D  	` �D  	` �����@ ��      F   ,���@ �����@ �\  	` �\  	` �����@ ��      F   ,���@ s���@ w�  	` w�  	` s���@ s      F   ,���@ \4���@ `�  	` `�  	` \4���@ \4      F   ,���@ B����@ GT  	` GT  	` B����@ B�      F   ,���@ )���@ -�  	` -�  	` )���@ )      F   ,���@ ,���@ �  	` �  	` ,���@ ,      F   ,���@ �����@ �L  	` �L  	` �����@ ��      F   ,���@ ����@ �  	` �  	` ����@ �      F   ,���@ �$���@ ��  	` ��  	` �$���@ �$      F   ,���@ �����@ �D  	` �D  	` �����@ ��      F   ,���@ ����@ ��  	` ��  	` ����@ �      F   ,���@ ~���@ ��  	` ��  	` ~���@ ~      F   ,���@ 
d����@ 
i<  	` 
i<  	` 
d����@ 
d�      F   ,���@ 	M����@ 	RT  	` 	RT  	` 	M����@ 	M�      F   ,���@ 4���@ 8�  	` 8�  	` 4���@ 4      F   ,���@ ����@ 4  	` 4  	` ����@ �      F   ,���@ ����@ L  	` L  	` ����@ �      F   ,���@ ����@ �  	` �  	` ����@ �      F   ,���@ �|���@ �,  	` �,  	` �|���@ �|      F   ,���@ �����@ �D  	` �D  	` �����@ ��      F   ,���@ ����@ ��  	` ��  	` ����@ �      F   ,���@  ����@  ��  	`  ��  	`  ����@  �      F   , ,�� �� ,�� Ǆ ,�  Ǆ ,�  �� ,�� ��      F   , ,�� �d ,�� � ,�  � ,�  �d ,�� �d      F   , ,�� 4 ,�� � ,�  � ,�  4 ,�� 4      F   , ,�� �L ,�� �� ,�  �� ,�  �L ,�� �L      F   , ,�� �� ,�� �4 ,�  �4 ,�  �� ,�� ��      F   , ,�� � ,�� � ,�  � ,�  � ,�� �      F   , ,��   ,�� $� ,�  $� ,�    ,��        F   , ,�� .l ,�� 3 ,�  3 ,�  .l ,�� .l      F   , ,�� ;� ,�� @\ ,�  @\ ,�  ;� ,�� ;�      F   , ,�� 
GT ,�� 
L ,�  
L ,�  
GT ,�� 
GT      F   , ,�� 	b� ,�� 	g� ,�  	g� ,�  	b� ,�� 	b�      F   , ,�� � ,�� �� ,�  �� ,�  � ,�� �      F   , ,�� ~t ,�� �$ ,�  �$ ,�  ~t ,�� ~t      F   , ,�� W< ,�� [� ,�  [� ,�  W< ,�� W<      F   , ,�� � ,�� �� ,�  �� ,�  � ,�� �      F   , ,�� � ,�� �� ,�  �� ,�  � ,�� �      F   , ,�� �� ,�� �� ,�  �� ,�  �� ,�� ��      F   , ,�� r� ,�� w| ,�  w| ,�  r� ,�� r�      F   , ,�� �| ,�� �, ,�  �, ,�  �| ,�� �|      F   , ,�� d| ,�� i, ,�  i, ,�  d| ,�� d|      F   , ,�� � ,�� � ,�  � ,�  � ,�� �      F   , ,�� � ,�� 
L ,�  
L ,�  � ,�� �      F   , ,�� �� ,�� �d ,�  �d ,�  �� ,�� ��      F   , ,�� � ,�� #4 ,�  #4 ,�  � ,�� �      F   , ,�� � ,�� �T ,�  �T ,�  � ,�� �      F   , ,�� : ,�� >� ,�  >� ,�  : ,�� :      F   , ,�� �D ,�� �� ,�  �� ,�  �D ,�� �D      F   , ,�� U� ,�� ZT ,�  ZT ,�  U� ,�� U�      F   , ,�� �� ,�� �L ,�  �L ,�  �� ,�� ��      F   , ,��  q4 ,��  u� ,�   u� ,�   q4 ,��  q4   	   G   !        +�  � +�  s� +P  s�   	   G   !       $ *��  � *�� � *�� � *�� o      G   ,��[<��p,��[< 6D���f� 6D���f���p,��[<��p,      G   ,��m4���$��m4 62���x� 62���x����$��m4���$      G   ,��,�����, 6 ����� 6 ����������,���      G   ,���$������$ 6����� 6�����������$���      G   ,��������� 5������ 5���������������      G   ,��������� 5����� 5��������������      G   ,���������� 5������ 5�����������������      G   ,���������� 5����� 5����������������      G   , ,����� ,� 5�� ,�� 5�� ,������ ,�����      G   , ,� ���� ,�  5�� ,Ÿ 5�� ,Ÿ���� ,� ����      G   , ,����� ,�� 5� ,װ 5� ,װ��� ,�����      G   , ,����� ,�� 5�� ,� 5�� ,���� ,�����      G   , ,����� ,�� 6� ,�� 6� ,����� ,�����      G   , -���� -� 6 � -� 6 � -���� -����      G   , -����$ -� 62� -� 62� -����$ -����$      G   , -%���p, -%� 6D� -1� 6D� -1���p, -%���p,      G   , $ 5�� $ 5�� � 5�� � 5�� $ 5��      G   , Tt 5�� Tt 6 � `, 6 � `, 5�� Tt 5��      G   , �� 5�� �� 6D� �| 6D� �| 5�� �� 5��      G   , 'd 5�� 'd 5�� 3 5�� 3 5�� 'd 5��      G   , m� 5�� m� 5�� yl 5�� yl 5�� m� 5��      G   , � 5�� � 6 � �� 6 � �� 5�� � 5��      G   , �T 5�� �T 6D�  6D�  5�� �T 5��      G   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      G   , �D 5�� �D 5�� �� 5�� �� 5�� �D 5��      G   , � 5�� � 6 � L 6 � L 5�� � 5��      G   , Y� 5�� Y� 6D� e� 6D� e� 5�� Y� 5��      G   , � 5�� � 5�� �< 5�� �< 5�� � 5��      G   , ,� 5�� ,� 5�� 8� 5�� 8� 5�� ,� 5��      G   , s$ 5�� s$ 6 � ~� 6 � ~� 5�� s$ 5��      G   , �t 5�� �t 6D� �, 6D� �, 5�� �t 5��      G   , F 5�� F 5�� Q� 5�� Q� 5�� F 5��      G   , �d 5�� �d 5�� � 5�� � 5�� �d 5��      G   , Ҵ 5�� Ҵ 6 � �l 6 � �l 5�� Ҵ 5��      G   ,  5��  6D� $� 6D� $� 5��  5��      G   , �� 5�� �� 5�� �\ 5�� �\ 5�� �� 5��      G   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      G   ,  2D 5��  2D 6 �  =� 6 �  =� 5��  2D 5��      G   ,  x� 5��  x� 6D�  �L 6D�  �L 5��  x� 5��      G   , !4 5�� !4 5�� !� 5�� !� 5�� !4 5��      G   , !K� 5�� !K� 5�� !W< 5�� !W< 5�� !K� 5��      G   , !�� 5�� !�� 6 � !�� 6 � !�� 5�� !�� 5��      G   , !�$ 5�� !�$ 6D� !�� 6D� !�� 5�� !�$ 5��      G   , "d� 5�� "d� 5�� "p| 5�� "p| 5�� "d� 5��      G   , "� 5�� "� 5�� "�� 5�� "�� 5�� "� 5��      G   , "�d 5�� "�d 6 � "� 6 � "� 5�� "�d 5��      G   , #7� 5�� #7� 6D� #Cl 6D� #Cl 5�� #7� 5��      G   , #�T 5�� #�T 5�� #� 5�� #� 5�� #�T 5��      G   , $
� 5�� $
� 5�� $\ 5�� $\ 5�� $
� 5��      G   , $P� 5�� $P� 6 � $\� 6 � $\� 5�� $P� 5��      G   , $�D 5�� $�D 6D� $�� 6D� $�� 5�� $�D 5��      G   , %#� 5�� %#� 5�� %/� 5�� %/� 5�� %#� 5��      G   , %j4 5�� %j4 5�� %u� 5�� %u� 5�� %j4 5��      G   , %�� 5�� %�� 6 � %�< 6 � %�< 5�� %�� 5��      G   , %�� 5�� %�� 6D� &� 6D� &� 5�� %�� 5��      G   , &�t 5�� &�t 5�� &�, 5�� &�, 5�� &�t 5��      G   , &�� 5�� &�� 5�� &�| 5�� &�| 5�� &�� 5��      G   , ' 5�� ' 6 � '� 6 � '� 5�� ' 5��      G   , 'Vd 5�� 'Vd 6D� 'b 6D� 'b 5�� 'Vd 5��      G   , '� 5�� '� 5�� '� 5�� '� 5�� '� 5��      G   , ()T 5�� ()T 5�� (5 5�� (5 5�� ()T 5��      G   , (o� 5�� (o� 6 � ({\ 6 � ({\ 5�� (o� 5��      G   , (�� 5�� (�� 6D� (�� 6D� (�� 5�� (�� 5��      G   , )B� 5�� )B� 5�� )NL 5�� )NL 5�� )B� 5��      G   , )�� 5�� )�� 5�� )�� 5�� )�� 5�� )�� 5��      G   , )�4 5�� )�4 6 � )�� 6 � )�� 5�� )�4 5��      G   , *� 5�� *� 6D� *!< 6D� *!< 5�� *� 5��      G   , *�$ 5�� *�$ 5�� *�� 5�� *�� 5�� *�$ 5��      G   , *�t 5�� *�t 5�� *�, 5�� *�, 5�� *�t 5��      G   , +.� 5�� +.� 6 � +:| 6 � +:| 5�� +.� 5��      G   , +u 5�� +u 6D� +�� 6D� +�� 5�� +u 5��      G   , ,� 5�� ,� 5�� ,l 5�� ,l 5�� ,� 5��      G   , ,H 5�� ,H 5�� ,S� 5�� ,S� 5�� ,H 5��      G   , O 5�� O 5�� Z� 5�� Z� 5�� O 5��      G   , �T 5�� �T 6 � � 6 � � 5�� �T 5��      G   , ۤ 5�� ۤ 6D� �\ 6D� �\ 5�� ۤ 5��      G   , hD 5�� hD 5�� s� 5�� s� 5�� hD 5��      G   , �� 5�� �� 5�� �L 5�� �L 5�� �� 5��      G   , �� 5�� �� 6 �  � 6 �  � 5�� �� 5��      G   , ;4 5�� ;4 6D� F� 6D� F� 5�� ;4 5��      G   , �� 5�� �� 5�� ӌ 5�� ӌ 5�� �� 5��      G   , �� 5�� �� 5�� ڌ 5�� ڌ 5�� �� 5��      G   , $ 5�� $ 5��  � 5��  � 5�� $ 5��      G   , [t 5�� [t 6 � g, 6 � g, 5�� [t 5��      G   , �� 5�� �� 6D� �| 6D� �| 5�� �� 5��      G   , .d 5�� .d 5�� : 5�� : 5�� .d 5��      G   , t� 5�� t� 5�� �l 5�� �l 5�� t� 5��      G   , � 5�� � 6 � Ƽ 6 � Ƽ 5�� � 5��      G   , T 5�� T 6D�  6D�  5�� T 5��      G   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      G   , �D 5�� �D 5�� �� 5�� �� 5�� �D 5��      G   , � 5�� � 6 � &L 6 � &L 5�� � 5��      G   , `� 5�� `� 6D� l� 6D� l� 5�� `� 5��      G   , � 5�� � 5�� �< 5�� �< 5�� � 5��      G   , 3� 5�� 3� 5�� ?� 5�� ?� 5�� 3� 5��      G   , z$ 5�� z$ 6 � �� 6 � �� 5�� z$ 5��      G   , �t 5�� �t 6D� �, 6D� �, 5�� �t 5��      G   , M 5�� M 5�� X� 5�� X� 5�� M 5��      G   , �d 5�� �d 5�� � 5�� � 5�� �d 5��      G   , ٴ 5�� ٴ 6 � �l 6 � �l 5�� ٴ 5��      G   , 	  5�� 	  6D� 	+� 6D� 	+� 5�� 	  5��      G   , 	�� 5�� 	�� 5�� 	�\ 5�� 	�\ 5�� 	�� 5��      G   , 	�� 5�� 	�� 5�� 	�� 5�� 	�� 5�� 	�� 5��      G   , 
9D 5�� 
9D 6 � 
D� 6 � 
D� 5�� 
9D 5��      G   , 
� 5�� 
� 6D� 
�L 6D� 
�L 5�� 
� 5��      G   , 4 5�� 4 5�� � 5�� � 5�� 4 5��      G   , R� 5�� R� 5�� ^< 5�� ^< 5�� R� 5��      G   , �� 5�� �� 6 � �� 6 � �� 5�� �� 5��      G   , �$ 5�� �$ 6D� �� 6D� �� 5�� �$ 5��      G   , k� 5�� k� 5�� w| 5�� w| 5�� k� 5��      G   , � 5�� � 5�� �� 5�� �� 5�� � 5��      G   , �d 5�� �d 6 �  6 �  5�� �d 5��      G   , >� 5�� >� 6D� Jl 6D� Jl 5�� >� 5��      G   , �T 5�� �T 5�� � 5�� � 5�� �T 5��      G   , � 5�� � 5�� \ 5�� \ 5�� � 5��      G   , W� 5�� W� 6 � c� 6 � c� 5�� W� 5��      G   , �D 5�� �D 6D� �� 6D� �� 5�� �D 5��      G   , *� 5�� *� 5�� 6� 5�� 6� 5�� *� 5��      G   , q4 5�� q4 5�� |� 5�� |� 5�� q4 5��      G   , �� 5�� �� 6 � �< 6 � �< 5�� �� 5��      G   , �� 5�� �� 6D� 	� 6D� 	� 5�� �� 5��      G   , �t 5�� �t 5�� �, 5�� �, 5�� �t 5��      G   , �� 5�� �� 5�� �| 5�� �| 5�� �� 5��      G   ,  5��  6 � "� 6 � "� 5��  5��      G   , ]d 5�� ]d 6D� i 6D� i 5�� ]d 5��      G   , � 5�� � 5�� �� 5�� �� 5�� � 5��      G   , 0T 5�� 0T 5�� < 5�� < 5�� 0T 5��      G   , v� 5�� v� 6 � �\ 6 � �\ 5�� v� 5��      G   , �� 5�� �� 6D� Ȭ 6D� Ȭ 5�� �� 5��      G   , I� 5�� I� 5�� UL 5�� UL 5�� I� 5��      G   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      G   , �4 5�� �4 6 � �� 6 � �� 5�� �4 5��      G   , � 5�� � 6D� (< 6D� (< 5�� � 5��      G   , �$ 5�� �$ 5�� �� 5�� �� 5�� �$ 5��      G   , �t 5�� �t 5�� �, 5�� �, 5�� �t 5��      G   , 5� 5�� 5� 6 � A| 6 � A| 5�� 5� 5��      G   , | 5�� | 6D� �� 6D� �� 5�� | 5��      G   , � 5�� � 5�� l 5�� l 5�� � 5��      G   ,  � 5��  � 5��  l 5��  l 5��  � 5��      G   ,  V 5��  V 5��  a� 5��  a� 5��  V 5��      G   ,  �T 5��  �T 6 �  � 6 �  � 5��  �T 5��      G   ,  � 5��  � 6D�  �\ 6D�  �\ 5��  � 5��      G   , oD 5�� oD 5�� z� 5�� z� 5�� oD 5��      G   , �� 5�� �� 5�� �L 5�� �L 5�� �� 5��      G   , �� 5�� �� 6 � � 6 � � 5�� �� 5��      G   , B4 5�� B4 6D� M� 6D� M� 5�� B4 5��      G   , ������ ��  	` ڌ  	` ڌ���� ������      G   , $��� $  	`  �  	`  ���� $���      G   , [t��� [t  	` g,  	` g,��� [t���      G   , ����p, ��  	` �|  	` �|��p, ����p,      G   , .d���� .d  	` :  	` :���� .d����      G   , t���� t�  	` �l  	` �l��� t����      G   , ���� �  	` Ƽ  	` Ƽ��� ����      G   , T��p, T  	`   	` ��p, T��p,      G   , ������ ��  	` ��  	` ������ ������      G   , �D��� �D  	` ��  	` ����� �D���      G   , ���� �  	` &L  	` &L��� ����      G   , `���p, `�  	` l�  	` l���p, `���p,      G   , ����� �  	` �<  	` �<���� �����      G   , 3���� 3�  	` ?�  	` ?���� 3����      G   , z$��� z$  	` ��  	` ����� z$���      G   , �t��p, �t  	` �,  	` �,��p, �t��p,      G   , M���� M  	` X�  	` X����� M����      G   , �d��� �d  	` �  	` ���� �d���      G   , ٴ��� ٴ  	` �l  	` �l��� ٴ���      G   , 	 ��p, 	   	` 	+�  	` 	+���p, 	 ��p,      G   , 	������ 	��  	` 	�\  	` 	�\���� 	������      G   , 	����� 	��  	` 	��  	` 	����� 	�����      G   , 
9D��� 
9D  	` 
D�  	` 
D���� 
9D���      G   , 
���p, 
�  	` 
�L  	` 
�L��p, 
���p,      G   , 4���� 4  	` �  	` ����� 4����      G   , R���� R�  	` ^<  	` ^<��� R����      G   , ����� ��  	` ��  	` ����� �����      G   , �$��p, �$  	` ��  	` ����p, �$��p,      G   , k����� k�  	` w|  	` w|���� k�����      G   , ���� �  	` ��  	` ����� ����      G   , �d��� �d  	`   	` ��� �d���      G   , >���p, >�  	` Jl  	` Jl��p, >���p,      G   , �T���� �T  	` �  	` ����� �T����      G   , ���� �  	` \  	` \��� ����      G   , W���� W�  	` c�  	` c���� W����      G   , �D��p, �D  	` ��  	` ����p, �D��p,      G   , *����� *�  	` 6�  	` 6����� *�����      G   , q4��� q4  	` |�  	` |���� q4���      G   , ����� ��  	` �<  	` �<��� �����      G   , ����p, ��  	` 	�  	` 	���p, ����p,      G   , �t���� �t  	` �,  	` �,���� �t����      G   , ����� ��  	` �|  	` �|��� �����      G   , ���   	` "�  	` "���� ���      G   , ]d��p, ]d  	` i  	` i��p, ]d��p,      G   , ����� �  	` ��  	` ������ �����      G   , 0T��� 0T  	` <  	` <��� 0T���      G   , v���� v�  	` �\  	` �\��� v����      G   , ����p, ��  	` Ȭ  	` Ȭ��p, ����p,      G   , I����� I�  	` UL  	` UL���� I�����      G   , ����� ��  	` ��  	` ����� �����      G   , �4��� �4  	` ��  	` ����� �4���      G   , ���p, �  	` (<  	` (<��p, ���p,      G   , �$���� �$  	` ��  	` ������ �$����      G   , �t��� �t  	` �,  	` �,��� �t���      G   , 5���� 5�  	` A|  	` A|��� 5����      G   , |��p, |  	` ��  	` ����p, |��p,      G   , ����� �  	` l  	` l���� �����      G   ,  �����  �  	`  l  	`  l����  �����      G   ,  V���  V  	`  a�  	`  a����  V���      G   ,  �T���  �T  	`  �  	`  ����  �T���      G   ,  ���p,  �  	`  �\  	`  �\��p,  ���p,      G   , oD���� oD  	` z�  	` z����� oD����      G   , ����� ��  	` �L  	` �L��� �����      G   , ����� ��  	` �  	` ���� �����      G   , B4��p, B4  	` M�  	` M���p, B4��p,      G   , $��� $  	` �  	` ���� $���      G   , Tt��� Tt  	` `,  	` `,��� Tt���      G   , ����p, ��  	` �|  	` �|��p, ����p,      G   , 'd���� 'd  	` 3  	` 3���� 'd����      G   , m���� m�  	` yl  	` yl��� m����      G   , ���� �  	` ��  	` ����� ����      G   , �T��p, �T  	`   	` ��p, �T��p,      G   , ������ ��  	` ��  	` ������ ������      G   , �D��� �D  	` ��  	` ����� �D���      G   , ���� �  	` L  	` L��� ����      G   , Y���p, Y�  	` e�  	` e���p, Y���p,      G   , ����� �  	` �<  	` �<���� �����      G   , ,���� ,�  	` 8�  	` 8���� ,����      G   , s$��� s$  	` ~�  	` ~���� s$���      G   , �t��p, �t  	` �,  	` �,��p, �t��p,      G   , F���� F  	` Q�  	` Q����� F����      G   , �d��� �d  	` �  	` ���� �d���      G   , Ҵ��� Ҵ  	` �l  	` �l��� Ҵ���      G   , ��p,   	` $�  	` $���p, ��p,      G   , ������ ��  	` �\  	` �\���� ������      G   , ����� ��  	` ��  	` ����� �����      G   ,  2D���  2D  	`  =�  	`  =����  2D���      G   ,  x���p,  x�  	`  �L  	`  �L��p,  x���p,      G   , !4���� !4  	` !�  	` !����� !4����      G   , !K���� !K�  	` !W<  	` !W<��� !K����      G   , !����� !��  	` !��  	` !����� !�����      G   , !�$��p, !�$  	` !��  	` !����p, !�$��p,      G   , "d����� "d�  	` "p|  	` "p|���� "d�����      G   , "���� "�  	` "��  	` "����� "����      G   , "�d��� "�d  	` "�  	` "���� "�d���      G   , #7���p, #7�  	` #Cl  	` #Cl��p, #7���p,      G   , #�T���� #�T  	` #�  	` #����� #�T����      G   , $
���� $
�  	` $\  	` $\��� $
����      G   , $P���� $P�  	` $\�  	` $\���� $P����      G   , $�D��p, $�D  	` $��  	` $����p, $�D��p,      G   , %#����� %#�  	` %/�  	` %/����� %#�����      G   , %j4��� %j4  	` %u�  	` %u���� %j4���      G   , %����� %��  	` %�<  	` %�<��� %�����      G   , %����p, %��  	` &�  	` &���p, %����p,      G   , &�t���� &�t  	` &�,  	` &�,���� &�t����      G   , &����� &��  	` &�|  	` &�|��� &�����      G   , '��� '  	` '�  	` '���� '���      G   , 'Vd��p, 'Vd  	` 'b  	` 'b��p, 'Vd��p,      G   , '����� '�  	` '�  	` '����� '�����      G   , ()T��� ()T  	` (5  	` (5��� ()T���      G   , (o���� (o�  	` ({\  	` ({\��� (o����      G   , (����p, (��  	` (��  	` (����p, (����p,      G   , )B����� )B�  	` )NL  	` )NL���� )B�����      G   , )����� )��  	` )��  	` )����� )�����      G   , )�4��� )�4  	` )��  	` )����� )�4���      G   , *���p, *�  	` *!<  	` *!<��p, *���p,      G   , *�$���� *�$  	` *��  	` *������ *�$����      G   , *�t��� *�t  	` *�,  	` *�,��� *�t���      G   , +.���� +.�  	` +:|  	` +:|��� +.����      G   , +u��p, +u  	` +��  	` +����p, +u��p,      G   , ,����� ,�  	` ,l  	` ,l���� ,�����      G   , ,H��� ,H  	` ,S�  	` ,S���� ,H���      G   , O��� O  	` Z�  	` Z���� O���      G   , �T��� �T  	` �  	` ���� �T���      G   , ۤ��p, ۤ  	` �\  	` �\��p, ۤ��p,      G   , hD���� hD  	` s�  	` s����� hD����      G   , ����� ��  	` �L  	` �L��� �����      G   , ����� ��  	`  �  	`  ���� �����      G   , ;4��p, ;4  	` F�  	` F���p, ;4��p,      G   , ������ ��  	` ӌ  	` ӌ���� ������      G  , , -, (�  -, (�  -	L (�  -	L (�  -, (�       G  , , (�@ 6@H (�@ 6Ch (�` 6Ch (�` 6@H (�@ 6@H      G  , , +y` 6@H +y` 6Ch +|� 6Ch +|� 6@H +y` 6@H      G  , , -* 6@H -* 6Ch --< 6Ch --< 6@H -* 6@H      G  , , (�@ 6: (�@ 6=( (�` 6=( (�` 6: (�@ 6:      G  , , +y` 6: +y` 6=( +|� 6=( +|� 6: +y` 6:      G  , , -* 6: -* 6=( --< 6=( --< 6: -* 6:      G  , , *� 6.P *� 61p *� 61p *� 6.P *� 6.P      G  , , -$ 6.P -$ 61p -D 61p -D 6.P -$ 6.P      G  , , *� 6( *� 6+0 *� 6+0 *� 6( *� 6(      G  , , -$ 6( -$ 6+0 -D 6+0 -D 6( -$ 6(      G  , , (s� 6X (s� 6x (w 6x (w 6X (s� 6X      G  , , +3 6X +3 6x +60 6x +60 6X +3 6X      G  , , -, 6X -, 6x -	L 6x -	L 6X -, 6X      G  , , (s� 6 (s� 68 (w 68 (w 6 (s� 6      G  , , +3 6 +3 68 +60 68 +60 6 +3 6      G  , , -, 6 -, 68 -	L 68 -	L 6 -, 6      G  , , )Ӏ 6
` )Ӏ 6� )֠ 6� )֠ 6
` )Ӏ 6
`      G  , , ,�4 6
` ,�4 6� ,�T 6� ,�T 6
` ,�4 6
`      G  , , )Ӏ 6  )Ӏ 6@ )֠ 6@ )֠ 6  )Ӏ 6       G  , , ,�4 6  ,�4 6@ ,�T 6@ ,�T 6  ,�4 6       G  , , (-� 5�h (-� 5�� (0� 5�� (0� 5�h (-� 5�h      G  , , *�� 5�h *�� 5�� *�� 5�� *�� 5�h *�� 5�h      G  , , ,�< 5�h ,�< 5�� ,�\ 5�� ,�\ 5�h ,�< 5�h      G  , , (-� 5�( (-� 5�H (0� 5�H (0� 5�( (-� 5�(      G  , , *�� 5�( *�� 5�H *�� 5�H *�� 5�( *�� 5�(      G  , , ,�< 5�( ,�< 5�H ,�\ 5�H ,�\ 5�( ,�< 5�(      G  , , )�0 5�p )�0 5� )�P 5� )�P 5�p )�0 5�p      G  , , ,LP 5�p ,LP 5� ,Op 5� ,Op 5�p ,LP 5�p      G  , , ,�D 5�p ,�D 5� ,�d 5� ,�d 5�p ,�D 5�p      G  , , )�0 5�0 )�0 5�P )�P 5�P )�P 5�0 )�0 5�0      G  , , ,LP 5�0 ,LP 5�P ,Op 5�P ,Op 5�0 ,LP 5�0      G  , , ,�D 5�0 ,�D 5�P ,�d 5�P ,�d 5�0 ,�D 5�0      G  , , '�P 5�x '�P 5ט '�p 5ט '�p 5�x '�P 5�x      G  , , *�p 5�x *�p 5ט *�� 5ט *�� 5�x *�p 5�x      G  , , ,�L 5�x ,�L 5ט ,�l 5ט ,�l 5�x ,�L 5�x      G  , , '�P 5�8 '�P 5�X '�p 5�X '�p 5�8 '�P 5�8      G  , , *�p 5�8 *�p 5�X *�� 5�X *�� 5�8 *�p 5�8      G  , , ,�L 5�8 ,�L 5�X ,�l 5�X ,�l 5�8 ,�L 5�8      G  , , )F� 5 )F� 5Š )J  5Š )J  5 )F� 5      G  , , ,  5 ,  5Š ,	  5Š ,	  5 ,  5      G  , , ,�T 5 ,�T 5Š ,�t 5Š ,�t 5 ,�T 5      G  , , )F� 5�@ )F� 5�` )J  5�` )J  5�@ )F� 5�@      G  , , ,  5�@ ,  5�` ,	  5�` ,	  5�@ ,  5�@      G  , , ,�T 5�@ ,�T 5�` ,�t 5�` ,�t 5�@ ,�T 5�@      G  , , -$ 5.` -$ 51� -D 51� -D 5.` -$ 5.`      G  , , -$ 5(  -$ 5+@ -D 5+@ -D 5(  -$ 5(       G  , , ,�4 4� ,�4 4�0 ,�T 4�0 ,�T 4� ,�4 4�      G  , , ,�4 4�� ,�4 4�� ,�T 4�� ,�T 4�� ,�4 4��      G  , , ,�D 4�� ,�D 4�� ,�d 4�� ,�d 4�� ,�D 4��      G  , , ,�D 4�� ,�D 4�� ,�d 4�� ,�d 4�� ,�D 4��      G  , , ,�T 4[p ,�T 4^� ,�t 4^� ,�t 4[p ,�T 4[p      G  , , ,�T 4U0 ,�T 4XP ,�t 4XP ,�t 4U0 ,�T 4U0      G  , , -* 3�� -* 3�� --< 3�� --< 3�� -* 3��      G  , , -* 3Ȑ -* 3˰ --< 3˰ --< 3Ȑ -* 3Ȑ      G  , , -, 3�� -, 3�� -	L 3�� -	L 3�� -, 3��      G  , , -, 3�@ -, 3�` -	L 3�` -	L 3�@ -, 3�@      G  , , ,�< 3B0 ,�< 3EP ,�\ 3EP ,�\ 3B0 ,�< 3B0      G  , , ,�< 3;� ,�< 3? ,�\ 3? ,�\ 3;� ,�< 3;�      G  , , ,�L 2�� ,�L 2�  ,�l 2�  ,�l 2�� ,�L 2��      G  , , ,�L 2�� ,�L 2�� ,�l 2�� ,�l 2�� ,�L 2��      G  , , -$ 2o@ -$ 2r` -D 2r` -D 2o@ -$ 2o@      G  , , -$ 2i  -$ 2l  -D 2l  -D 2i  -$ 2i       G  , , ,�4 2(� ,�4 2, ,�T 2, ,�T 2(� ,�4 2(�      G  , , ,�4 2"� ,�4 2%� ,�T 2%� ,�T 2"� ,�4 2"�      G  , , ,�D 1� ,�D 1�� ,�d 1�� ,�d 1� ,�D 1�      G  , , ,�D 1�` ,�D 1߀ ,�d 1߀ ,�d 1�` ,�D 1�`      G  , , ,�T 1�P ,�T 1�p ,�t 1�p ,�t 1�P ,�T 1�P      G  , , ,�T 1� ,�T 1�0 ,�t 1�0 ,�t 1� ,�T 1�      G  , , -* 1� -* 1� --< 1� --< 1� -* 1�      G  , , -* 1	p -* 1� --< 1� --< 1	p -* 1	p      G  , , -, 0�` -, 0̀ -	L 0̀ -	L 0�` -, 0�`      G  , , -, 0�  -, 0�@ -	L 0�@ -	L 0�  -, 0�       G  , , ,�< 0� ,�< 0�0 ,�\ 0�0 ,�\ 0� ,�< 0�      G  , , ,�< 0|� ,�< 0� ,�\ 0� ,�\ 0|� ,�< 0|�      G  , , ,�L 0<� ,�L 0?� ,�l 0?� ,�l 0<� ,�L 0<�      G  , , ,�L 06� ,�L 09� ,�l 09� ,�l 06� ,�L 06�      G  , , -$ /�  -$ /�@ -D /�@ -D /�  -$ /�       G  , , -$ /�� -$ /�  -D /�  -D /�� -$ /��      G  , , ,�4 /i� ,�4 /l� ,�T /l� ,�T /i� ,�4 /i�      G  , , %�� 6 %�� 68 %�� 68 %�� 6 %�� 6      G  , , $� 5�p $� 5� $ 5� $ 5�p $� 5�p      G  , , &� 5�p &� 5� &�0 5� &�0 5�p &� 5�p      G  , , #<  6: #<  6=( #?  6=( #?  6: #<  6:      G  , , !�p 6( !�p 6+0 !ߐ 6+0 !ߐ 6( !�p 6(      G  , , $�� 6( $�� 6+0 $�� 6+0 $�� 6( $�� 6(      G  , , $� 5�0 $� 5�P $ 5�P $ 5�0 $� 5�0      G  , , &� 5�0 &� 5�P &�0 5�P &�0 5�0 &� 5�0      G  , , $U@ 6
` $U@ 6� $X` 6� $X` 6
` $U@ 6
`      G  , , '` 6
` '` 6� '� 6� '� 6
` '` 6
`      G  , , 'Z� 6( 'Z� 6+0 ']� 6+0 ']� 6( 'Z� 6(      G  , , "i 5�x "i 5ט "l0 5ט "l0 5�x "i 5�x      G  , , %(0 5�x %(0 5ט %+P 5ט %+P 5�x %(0 5�x      G  , , %�  6: %�  6=( %�@ 6=( %�@ 6: %�  6:      G  , , $U@ 6  $U@ 6@ $X` 6@ $X` 6  $U@ 6       G  , , '` 6  '` 6@ '� 6@ '� 6  '` 6       G  , , "i 5�8 "i 5�X "l0 5�X "l0 5�8 "i 5�8      G  , , %(0 5�8 %(0 5�X %+P 5�X %+P 5�8 %(0 5�8      G  , , !�p 6.P !�p 61p !ߐ 61p !ߐ 6.P !�p 6.P      G  , , "�� 6X "�� 6x "�� 6x "�� 6X "�� 6X      G  , , "�` 5�h "�` 5�� "�� 5�� "�� 5�h "�` 5�h      G  , , #Ƞ 5 #Ƞ 5Š #�� 5Š #�� 5 #Ƞ 5      G  , , &�� 5 &�� 5Š &�� 5Š &�� 5 &�� 5      G  , , %n� 5�h %n� 5�� %q� 5�� %q� 5�h %n� 5�h      G  , , %�� 6X %�� 6x %�� 6x %�� 6X %�� 6X      G  , , $�� 6.P $�� 61p $�� 61p $�� 6.P $�� 6.P      G  , , #Ƞ 5�@ #Ƞ 5�` #�� 5�` #�� 5�@ #Ƞ 5�@      G  , , &�� 5�@ &�� 5�` &�� 5�` &�� 5�@ &�� 5�@      G  , , 'Z� 6.P 'Z� 61p ']� 61p ']� 6.P 'Z� 6.P      G  , , "�` 5�( "�` 5�H "�� 5�H "�� 5�( "�` 5�(      G  , , %n� 5�( %n� 5�H %q� 5�H %q� 5�( %n� 5�(      G  , , %�  6@H %�  6Ch %�@ 6Ch %�@ 6@H %�  6@H      G  , , "�� 6 "�� 68 "�� 68 "�� 6 "�� 6      G  , , #<  6@H #<  6Ch #?  6Ch #?  6@H #<  6@H      G  , , ,�D /#� ,�D /&� ,�d /&� ,�d /#� ,�D /#�      G  , , ,�D /@ ,�D / ` ,�d / ` ,�d /@ ,�D /@      G  , , ,�T .�0 ,�T .�P ,�t .�P ,�t .�0 ,�T .�0      G  , , ,�T .�� ,�T .� ,�t .� ,�t .�� ,�T .��      G  , , -* .P� -* .S� --< .S� --< .P� -* .P�      G  , , -* .JP -* .Mp --< .Mp --< .JP -* .JP      G  , , -, .
@ -, .` -	L .` -	L .
@ -, .
@      G  , , -, .  -, .  -	L .  -	L .  -, .       G  , , ,�< -�� ,�< -� ,�\ -� ,�\ -�� ,�< -��      G  , , ,�< -�� ,�< -�� ,�\ -�� ,�\ -�� ,�< -��      G  , , ,�L -}� ,�L -�� ,�l -�� ,�l -}� ,�L -}�      G  , , ,�L -w` ,�L -z� ,�l -z� ,�l -w` ,�L -w`      G  , , -$ ,�  -$ ,�  -D ,�  -D ,�  -$ ,�       G  , , -$ ,�� -$ ,�� -D ,�� -D ,�� -$ ,��      G  , , ,�4 ,�� ,�4 ,�� ,�T ,�� ,�T ,�� ,�4 ,��      G  , , ,�4 ,�p ,�4 ,�� ,�T ,�� ,�T ,�p ,�4 ,�p      G  , , ,�D ,d` ,�D ,g� ,�d ,g� ,�d ,d` ,�D ,d`      G  , , ,�D ,^  ,�D ,a@ ,�d ,a@ ,�d ,^  ,�D ,^       G  , , ,�T , ,�T ,!0 ,�t ,!0 ,�t , ,�T ,      G  , , ,�T ,� ,�T ,� ,�t ,� ,�t ,� ,�T ,�      G  , , -* +�p -* +�� --< +�� --< +�p -* +�p      G  , , -* +�0 -* +�P --< +�P --< +�0 -* +�0      G  , , -, +K  -, +N@ -	L +N@ -	L +K  -, +K       G  , , -, +D� -, +H  -	L +H  -	L +D� -, +D�      G  , , ,�< +� ,�< +� ,�\ +� ,�\ +� ,�< +�      G  , , ,�< *�� ,�< +� ,�\ +� ,�\ *�� ,�< *��      G  , , ,�L *�� ,�L *�� ,�l *�� ,�l *�� ,�L *��      G  , , ,�L *�@ ,�L *�` ,�l *�` ,�l *�@ ,�L *�@      G  , , -$ *1� -$ *5  -D *5  -D *1� -$ *1�      G  , , -$ *+� -$ *.� -D *.� -D *+� -$ *+�      G  , , ,�4 )� ,�4 )� ,�T )� ,�T )� ,�4 )�      G  , , ,�4 )�P ,�4 )�p ,�T )�p ,�T )�P ,�4 )�P      G  , , ,�D )�@ ,�D )�` ,�d )�` ,�d )�@ ,�D )�@      G  , , ,�D )�  ,�D )�  ,�d )�  ,�d )�  ,�D )�       G  , , ,�T )^� ,�T )b ,�t )b ,�t )^� ,�T )^�      G  , , ,�T )X� ,�T )[� ,�t )[� ,�t )X� ,�T )X�      G  , , -* (�P -* (�p --< (�p --< (�P -* (�P      G  , , -* (� -* (�0 --< (�0 --< (� -* (�      G  , , ,�4 /c� ,�4 /f� ,�T /f� ,�T /c� ,�4 /c�      G  , , �� 6: �� 6=( �� 6=( �� 6: �� 6:      G  , ,  |� 6:  |� 6=(  �  6=(  �  6:  |� 6:      G  , , �0 6 �0 68 �P 68 �P 6 �0 6      G  , , �P 6 �P 68 �p 68 �p 6 �P 6      G  , , wp 6 wp 68 z� 68 z� 6 wp 6      G  , , SP 5�p SP 5� Vp 5� Vp 5�p SP 5�p      G  , , p 5�p p 5� � 5� � 5�p p 5�p      G  , , ѐ 5�p ѐ 5� ԰ 5� ԰ 5�p ѐ 5�p      G  , , �� 5�p �� 5� �� 5� �� 5�p �� 5�p      G  , , !O� 5�p !O� 5� !R� 5� !R� 5�p !O� 5�p      G  , ,  6� 6  6� 68  9� 68  9� 6  6� 6      G  , , �� 6@H �� 6Ch � 6Ch � 6@H �� 6@H      G  , , �� 6@H �� 6Ch �� 6Ch �� 6@H �� 6@H      G  , , �� 6( �� 6+0 � 6+0 � 6( �� 6(      G  , , � 6( � 6+0 �0 6+0 �0 6( � 6(      G  , , SP 5�0 SP 5�P Vp 5�P Vp 5�0 SP 5�0      G  , , p 5�0 p 5�P � 5�P � 5�0 p 5�0      G  , , ѐ 5�0 ѐ 5�P ԰ 5�P ԰ 5�0 ѐ 5�0      G  , , �� 5�0 �� 5�P �� 5�P �� 5�0 �� 5�0      G  , , !O� 5�0 !O� 5�P !R� 5�P !R� 5�0 !O� 5�0      G  , , ^0 6( ^0 6+0 aP 6+0 aP 6( ^0 6(      G  , , �� 6
` �� 6� �� 6� �� 6
` �� 6
`      G  , , X� 6
` X� 6� [� 6� [� 6
` X� 6
`      G  , , � 6
` � 6�   6�   6
` � 6
`      G  , , �  6
` �  6� �  6� �  6
` �  6
`      G  , , l� 5�x l� 5ט o� 5ט o� 5�x l� 5�x      G  , , +� 5�x +� 5ט .� 5ט .� 5�x +� 5�x      G  , , �� 5�x �� 5ט �� 5ט �� 5�x �� 5�x      G  , , �� 5�x �� 5ט � 5ט � 5�x �� 5�x      G  , , !�  6
` !�  6� !�@ 6� !�@ 6
` !�  6
`      G  , , P 6( P 6+0  p 6+0  p 6( P 6(      G  , ,  |� 6@H  |� 6Ch  �  6Ch  �  6@H  |� 6@H      G  , , ?� 6@H ?� 6Ch B� 6Ch B� 6@H ?� 6@H      G  , , ?� 6: ?� 6=( B� 6=( B� 6: ?� 6:      G  , , l� 5�8 l� 5�X o� 5�X o� 5�8 l� 5�8      G  , , +� 5�8 +� 5�X .� 5�X .� 5�8 +� 5�8      G  , , �� 5�8 �� 5�X �� 5�X �� 5�8 �� 5�8      G  , , �� 5�8 �� 5�X � 5�X � 5�8 �� 5�8      G  , , �� 6  �� 6@ �� 6@ �� 6  �� 6       G  , , X� 6  X� 6@ [� 6@ [� 6  X� 6       G  , , � 6  � 6@   6@   6  � 6       G  , , �  6  �  6@ �  6@ �  6  �  6       G  , , !�  6  !�  6@ !�@ 6@ !�@ 6  !�  6       G  , , �  5 �  5Š �@ 5Š �@ 5 �  5      G  , , �@ 5 �@ 5Š �` 5Š �` 5 �@ 5      G  , , J` 5 J` 5Š M� 5Š M� 5 J` 5      G  , , !	� 5 !	� 5Š !� 5Š !� 5 !	� 5      G  , , �� 6.P �� 61p � 61p � 6.P �� 6.P      G  , , � 6.P � 61p �0 61p �0 6.P � 6.P      G  , , �0 6X �0 6x �P 6x �P 6X �0 6X      G  , , �P 6X �P 6x �p 6x �p 6X �P 6X      G  , , �� 5�h �� 5�� �  5�� �  5�h �� 5�h      G  , , �  5�@ �  5�` �@ 5�` �@ 5�@ �  5�@      G  , , �@ 5�@ �@ 5�` �` 5�` �` 5�@ �@ 5�@      G  , , J` 5�@ J` 5�` M� 5�` M� 5�@ J` 5�@      G  , , !	� 5�@ !	� 5�` !� 5�` !� 5�@ !	� 5�@      G  , , r  5�h r  5�� u  5�� u  5�h r  5�h      G  , , 1  5�h 1  5�� 4@ 5�� 4@ 5�h 1  5�h      G  , , �@ 5�h �@ 5�� �` 5�� �` 5�h �@ 5�h      G  , , wp 6X wp 6x z� 6x z� 6X wp 6X      G  , ,  6� 6X  6� 6x  9� 6x  9� 6X  6� 6X      G  , , ^0 6.P ^0 61p aP 61p aP 6.P ^0 6.P      G  , , P 6.P P 61p  p 61p  p 6.P P 6.P      G  , , �� 6: �� 6=( � 6=( � 6: �� 6:      G  , , �� 5�( �� 5�H �  5�H �  5�( �� 5�(      G  , , r  5�( r  5�H u  5�H u  5�( r  5�(      G  , , 1  5�( 1  5�H 4@ 5�H 4@ 5�( 1  5�(      G  , , �@ 5�( �@ 5�H �` 5�H �` 5�( �@ 5�(      G  , , -, (�� -, (�� -	L (�� -	L (�� -, (��      G  , , ,�< (E� ,�< (H� ,�\ (H� ,�\ (E� ,�< (E�      G  , , ,�< (?p ,�< (B� ,�\ (B� ,�\ (?p ,�< (?p      G  , , ,�L '�` ,�L (� ,�l (� ,�l '�` ,�L '�`      G  , , ,�L '�  ,�L '�@ ,�l '�@ ,�l '�  ,�L '�       G  , , -$ 'r� -$ 'u� -D 'u� -D 'r� -$ 'r�      G  , , -$ 'l� -$ 'o� -D 'o� -D 'l� -$ 'l�      G  , , ,�4 ',p ,�4 '/� ,�T '/� ,�T ',p ,�4 ',p      G  , , ,�4 '&0 ,�4 ')P ,�T ')P ,�T '&0 ,�4 '&0      G  , , ,�D &�  ,�D &�@ ,�d &�@ ,�d &�  ,�D &�       G  , , ,�D &�� ,�D &�  ,�d &�  ,�d &�� ,�D &��      G  , , ,�T &�� ,�T &�� ,�t &�� ,�t &�� ,�T &��      G  , , ,�T &�� ,�T &�� ,�t &�� ,�t &�� ,�T &��      G  , , -* &0 -* &P --< &P --< &0 -* &0      G  , , -* &� -* & --< & --< &� -* &�      G  , , -, %�� -, %�  -	L %�  -	L %�� -, %��      G  , , -, %Ơ -, %�� -	L %�� -	L %Ơ -, %Ơ      G  , , ,�< %�� ,�< %�� ,�\ %�� ,�\ %�� ,�< %��      G  , , ,�< %�P ,�< %�p ,�\ %�p ,�\ %�P ,�< %�P      G  , , ,�L %@@ ,�L %C` ,�l %C` ,�l %@@ ,�L %@@      G  , , ,�L %:  ,�L %=  ,�l %=  ,�l %:  ,�L %:       G  , , -$ $�� -$ $�� -D $�� -D $�� -$ $��      G  , , -$ $�` -$ $�� -D $�� -D $�` -$ $�`      G  , , ,�4 $mP ,�4 $pp ,�T $pp ,�T $mP ,�4 $mP      G  , , ,�4 $g ,�4 $j0 ,�T $j0 ,�T $g ,�4 $g      G  , , ,�D $'  ,�D $*  ,�d $*  ,�d $'  ,�D $'       G  , , ,�D $ � ,�D $#� ,�d $#� ,�d $ � ,�D $ �      G  , , ,�T #� ,�T #�� ,�t #�� ,�t #� ,�T #�      G  , , ,�T #�p ,�T #ݐ ,�t #ݐ ,�t #�p ,�T #�p      G  , , -* #T -* #W0 --< #W0 --< #T -* #T      G  , , -* #M� -* #P� --< #P� --< #M� -* #M�      G  , , -, #� -, #� -	L #� -	L #� -, #�      G  , , -, #� -, #
� -	L #
� -	L #� -, #�      G  , , ,�< "�p ,�< "ʐ ,�\ "ʐ ,�\ "�p ,�< "�p      G  , , ,�< "�0 ,�< "�P ,�\ "�P ,�\ "�0 ,�< "�0      G  , , ,�L "�  ,�L "�@ ,�l "�@ ,�l "�  ,�L "�       G  , , ,�L "z� ,�L "~  ,�l "~  ,�l "z� ,�L "z�      G  , , -$ !� -$ !�� -D !�� -D !� -$ !�      G  , , -$ !�@ -$ !�` -D !�` -D !�@ -$ !�@      G  , , ,�4 !�0 ,�4 !�P ,�T !�P ,�T !�0 ,�4 !�0      G  , , ,�4 !�� ,�4 !� ,�T !� ,�T !�� ,�4 !��      G  , , ,�D !g� ,�D !k  ,�d !k  ,�d !g� ,�D !g�      G  , , ,�D !a� ,�D !d� ,�d !d� ,�d !a� ,�D !a�      G  , , ,�T !!� ,�T !$� ,�t !$� ,�t !!� ,�T !!�      G  , , ,�T !P ,�T !p ,�t !p ,�t !P ,�T !P      G  , , -*  �� -*  � --<  � --<  �� -*  ��      G  , , -*  �� -*  �� --<  �� --<  �� -*  ��      G  , , -,  N� -,  Q� -	L  Q� -	L  N� -,  N�      G  , , -,  H` -,  K� -	L  K� -	L  H` -,  H`      G  , , ,�<  P ,�<  p ,�\  p ,�\  P ,�<  P      G  , , ,�<   ,�<  0 ,�\  0 ,�\   ,�<        G  , , ,�L �  ,�L �  ,�l �  ,�l �  ,�L �       G  , , ,�L �� ,�L �� ,�l �� ,�l �� ,�L ��      G  , , -$ 5` -$ 8� -D 8� -D 5` -$ 5`      G  , , -$ /  -$ 2@ -D 2@ -D /  -$ /       G  , , ,�4 � ,�4 �0 ,�T �0 ,�T � ,�4 �      G  , , ,�4 �� ,�4 �� ,�T �� ,�T �� ,�4 ��      G  , , ,�D �� ,�D �� ,�d �� ,�d �� ,�D ��      G  , , ,�D �� ,�D �� ,�d �� ,�d �� ,�D ��      G  , , ,�T bp ,�T e� ,�t e� ,�t bp ,�T bp      G  , , ,�T \0 ,�T _P ,�t _P ,�t \0 ,�T \0      G  , , -* �� -* �� --< �� --< �� -* ��      G  , , -* ϐ -* Ұ --< Ұ --< ϐ -* ϐ      G  , , -, �� -, �� -	L �� -	L �� -, ��      G  , , -, �@ -, �` -	L �` -	L �@ -, �@      G  , , ,�< I0 ,�< LP ,�\ LP ,�\ I0 ,�< I0      G  , , ,�< B� ,�< F ,�\ F ,�\ B� ,�< B�      G  , , ,�L � ,�L   ,�l   ,�l � ,�L �      G  , , ,�L �� ,�L �� ,�l �� ,�l �� ,�L ��      G  , , -$ v@ -$ y` -D y` -D v@ -$ v@      G  , , -$ p  -$ s  -D s  -D p  -$ p       G  , , ,�4 /� ,�4 3 ,�T 3 ,�T /� ,�4 /�      G  , , ,�4 )� ,�4 ,� ,�T ,� ,�T )� ,�4 )�      G  , , ,�D � ,�D �� ,�d �� ,�d � ,�D �      G  , , ,�D �` ,�D � ,�d � ,�d �` ,�D �`      G  , , ,�T �P ,�T �p ,�t �p ,�t �P ,�T �P      G  , , ,�T � ,�T �0 ,�t �0 ,�t � ,�T �      G  , , -* � -* � --< � --< � -* �      G  , , -* p -* � --< � --< p -* p      G  , ,���x (� ���x (� ���� (� ���� (� ���x (�       G  , , 4� 5�h 4� 5�� 7� 5�� 7� 5�h 4� 5�h      G  , , �� 5�h �� 5�� �� 5�� �� 5�h �� 5�h      G  , , �� 6X �� 6x �� 6x �� 6X �� 6X      G  , , �� 6X �� 6x �� 6x �� 6X �� 6X      G  , , z� 6X z� 6x ~ 6x ~ 6X z� 6X      G  , , : 6X : 6x =0 6x =0 6X : 6X      G  , , �` 5�( �` 5�H �� 5�H �� 5�( �` 5�(      G  , , u� 5�( u� 5�H x� 5�H x� 5�( u� 5�(      G  , , 4� 5�( 4� 5�H 7� 5�H 7� 5�( 4� 5�(      G  , , �� 5�( �� 5�H �� 5�H �� 5�( �� 5�(      G  , , �p 6.P �p 61p � 61p � 6.P �p 6.P      G  , , �� 6.P �� 61p �� 61p �� 6.P �� 6.P      G  , , a� 6.P a� 61p d� 61p d� 6.P a� 6.P      G  , ,  � 6.P  � 61p #� 61p #� 6.P  � 6.P      G  , , V� 5�p V� 5� Y� 5� Y� 5�p V� 5�p      G  , , � 5�p � 5�  5�  5�p � 5�p      G  , , � 5�p � 5� �0 5� �0 5�p � 5�p      G  , , �0 5�p �0 5� �P 5� �P 5�p �0 5�p      G  , , �� 6 �� 68 �� 68 �� 6 �� 6      G  , , �� 6 �� 68 �� 68 �� 6 �� 6      G  , , z� 6 z� 68 ~ 68 ~ 6 z� 6      G  , , : 6 : 68 =0 68 =0 6 : 6      G  , , V� 5�0 V� 5�P Y� 5�P Y� 5�0 V� 5�0      G  , , � 5�0 � 5�P  5�P  5�0 � 5�0      G  , , � 5�0 � 5�P �0 5�P �0 5�0 � 5�0      G  , , �0 5�0 �0 5�P �P 5�P �P 5�0 �0 5�0      G  , , C  6: C  6=( F  6=( F  6: C  6:      G  , ,   6:   6=( @ 6=( @ 6:   6:      G  , , �@ 6: �@ 6=( �` 6=( �` 6: �@ 6:      G  , , �` 6: �` 6=( �� 6=( �� 6: �` 6:      G  , , u� 5�h u� 5�� x� 5�� x� 5�h u� 5�h      G  , , p 5�x p 5ט s0 5ט s0 5�x p 5�x      G  , , /0 5�x /0 5ט 2P 5ט 2P 5�x /0 5�x      G  , , �P 5�x �P 5ט �p 5ט �p 5�x �P 5�x      G  , , �p 5�x �p 5ט �� 5ט �� 5�x �p 5�x      G  , , �  6
` �  6� �@ 6� �@ 6
` �  6
`      G  , , \@ 6
` \@ 6� _` 6� _` 6
` \@ 6
`      G  , , ` 6
` ` 6� � 6� � 6
` ` 6
`      G  , , ڀ 6
` ڀ 6� ݠ 6� ݠ 6
` ڀ 6
`      G  , , p 5�8 p 5�X s0 5�X s0 5�8 p 5�8      G  , , /0 5�8 /0 5�X 2P 5�X 2P 5�8 /0 5�8      G  , , �P 5�8 �P 5�X �p 5�X �p 5�8 �P 5�8      G  , , �p 5�8 �p 5�X �� 5�X �� 5�8 �p 5�8      G  , , �p 6( �p 6+0 � 6+0 � 6( �p 6(      G  , , �� 6( �� 6+0 �� 6+0 �� 6( �� 6(      G  , , a� 6( a� 6+0 d� 6+0 d� 6( a� 6(      G  , ,  � 6(  � 6+0 #� 6+0 #� 6(  � 6(      G  , , � 5 � 5Š � 5Š � 5 � 5      G  , , Ϡ 5 Ϡ 5Š �� 5Š �� 5 Ϡ 5      G  , , �� 5 �� 5Š �� 5Š �� 5 �� 5      G  , , M� 5 M� 5Š Q  5Š Q  5 M� 5      G  , ,   5   5Š   5Š   5   5      G  , , �  6  �  6@ �@ 6@ �@ 6  �  6       G  , , \@ 6  \@ 6@ _` 6@ _` 6  \@ 6       G  , , ` 6  ` 6@ � 6@ � 6  ` 6       G  , , ڀ 6  ڀ 6@ ݠ 6@ ݠ 6  ڀ 6       G  , , � 5�@ � 5�` � 5�` � 5�@ � 5�@      G  , , Ϡ 5�@ Ϡ 5�` �� 5�` �� 5�@ Ϡ 5�@      G  , , �� 5�@ �� 5�` �� 5�` �� 5�@ �� 5�@      G  , , M� 5�@ M� 5�` Q  5�` Q  5�@ M� 5�@      G  , ,   5�@   5�`   5�`   5�@   5�@      G  , , C  6@H C  6Ch F  6Ch F  6@H C  6@H      G  , ,   6@H   6Ch @ 6Ch @ 6@H   6@H      G  , , �@ 6@H �@ 6Ch �` 6Ch �` 6@H �@ 6@H      G  , , �` 6@H �` 6Ch �� 6Ch �� 6@H �` 6@H      G  , , �` 5�h �` 5�� �� 5�� �� 5�h �` 5�h      G  , , ؐ 5�p ؐ 5� ۰ 5� ۰ 5�p ؐ 5�p      G  , , �� 5�p �� 5� �� 5� �� 5�p �� 5�p      G  , , 
=� 6X 
=� 6x 
@� 6x 
@� 6X 
=� 6X      G  , , ~p 6 ~p 68 �� 68 �� 6 ~p 6      G  , , 
=� 6 
=� 68 
@� 68 
@� 6 
=� 6      G  , , ؐ 5�0 ؐ 5�P ۰ 5�P ۰ 5�0 ؐ 5�0      G  , , �� 5�0 �� 5�P �� 5�P �� 5�0 �� 5�0      G  , , �� 6: �� 6=( �� 6=( �� 6: �� 6:      G  , , 
�� 6: 
�� 6=( 
�  6=( 
�  6: 
�� 6:      G  , , 8  5�( 8  5�H ;@ 5�H ;@ 5�( 8  5�(      G  , , �� 5�x �� 5ט �� 5ט �� 5�x �� 5�x      G  , , 	�� 5�x 	�� 5ט 	� 5ט 	� 5�x 	�� 5�x      G  , , 	�@ 5�( 	�@ 5�H 	�` 5�H 	�` 5�( 	�@ 5�(      G  , , � 6
` � 6� "  6� "  6
` � 6
`      G  , , �  6
` �  6� �  6� �  6
` �  6
`      G  , , �� 5�8 �� 5�X �� 5�X �� 5�8 �� 5�8      G  , , 	�� 5�8 	�� 5�X 	� 5�X 	� 5�8 	�� 5�8      G  , , e0 6( e0 6+0 hP 6+0 hP 6( e0 6(      G  , , 	$P 6( 	$P 6+0 	'p 6+0 	'p 6( 	$P 6(      G  , , �@ 5 �@ 5Š �` 5Š �` 5 �@ 5      G  , , Q` 5 Q` 5Š T� 5Š T� 5 Q` 5      G  , , e0 6.P e0 61p hP 61p hP 6.P e0 6.P      G  , , 	$P 6.P 	$P 61p 	'p 61p 	'p 6.P 	$P 6.P      G  , , � 6  � 6@ "  6@ "  6  � 6       G  , , �  6  �  6@ �  6@ �  6  �  6       G  , , �@ 5�@ �@ 5�` �` 5�` �` 5�@ �@ 5�@      G  , , Q` 5�@ Q` 5�` T� 5�` T� 5�@ Q` 5�@      G  , , ~p 6X ~p 6x �� 6x �� 6X ~p 6X      G  , , �� 6@H �� 6Ch �� 6Ch �� 6@H �� 6@H      G  , , 
�� 6@H 
�� 6Ch 
�  6Ch 
�  6@H 
�� 6@H      G  , , 8  5�h 8  5�� ;@ 5�� ;@ 5�h 8  5�h      G  , , 	�@ 5�h 	�@ 5�� 	�` 5�� 	�` 5�h 	�@ 5�h      G  , ,���p 2"����p 2%����� 2%����� 2"����p 2"�      G  , ,���p 6
`���p 6����� 6����� 6
`���p 6
`      G  , ,  �� 6
`  �� 6�  �� 6�  �� 6
`  �� 6
`      G  , ,���X 5�x���X 5ט���x 5ט���x 5�x���X 5�x      G  , , s� 5�x s� 5ט v� 5ט v� 5�x s� 5�x      G  , ,���h 3B0���h 3EP���� 3EP���� 3B0���h 3B0      G  , , 2� 5�x 2� 5ט 5� 5ט 5� 5�x 2� 5�x      G  , ,���` 4�����` 4������ 4������ 4�����` 4��      G  , ,���P 4[p���P 4^����p 4^����p 4[p���P 4[p      G  , ,���` 1����` 1������ 1������ 1����` 1�      G  , ,���X 2�����X 2� ���x 2� ���x 2�����X 2��      G  , ,���` 1�`���` 1߀���� 1߀���� 1�`���` 1�`      G  , ,���x 6X���x 6x���� 6x���� 6X���x 6X      G  , , _� 6
` _� 6� b� 6� b� 6
` _� 6
`      G  , ,���` 4�����` 4������ 4������ 4�����` 4��      G  , ,���X 2�����X 2�����x 2�����x 2�����X 2��      G  , ,���P 1�P���P 1�p���p 1�p���p 1�P���P 1�P      G  , ,��_� 3����_� 3����b� 3����b� 3����_� 3��      G  , ,���P 1����P 1�0���p 1�0���p 1����P 1�      G  , ,  0 6X  0 6x P 6x P 6X  0 6X      G  , ,��q� 6(��q� 6+0��t� 6+0��t� 6(��q� 6(      G  , ,  �� 6(  �� 6+0  � 6+0  � 6(  �� 6(      G  , ,���X 5�8���X 5�X���x 5�X���x 5�8���X 5�8      G  , , s� 5�8 s� 5�X v� 5�X v� 5�8 s� 5�8      G  , , 2� 5�8 2� 5�X 5� 5�X 5� 5�8 2� 5�8      G  , ,��_� 6:��_� 6=(��b� 6=(��b� 6:��_� 6:      G  , ,���` 5�0���` 5�P���� 5�P���� 5�0���` 5�0      G  , ,��_� 1���_� 1���b� 1���b� 1���_� 1�      G  , ,��_� 3Ȑ��_� 3˰��b� 3˰��b� 3Ȑ��_� 3Ȑ      G  , ,��_� 1	p��_� 1���b� 1���b� 1	p��_� 1	p      G  , ,��q� 6.P��q� 61p��t� 61p��t� 6.P��q� 6.P      G  , , � 6( � 6+0 �0 6+0 �0 6( � 6(      G  , ,  ZP 5�0  ZP 5�P  ]p 5�P  ]p 5�0  ZP 5�0      G  , , p 5�0 p 5�P � 5�P � 5�0 p 5�0      G  , ,���x 0�`���x 0̀���� 0̀���� 0�`���x 0�`      G  , ,  �� 6.P  �� 61p  � 61p  � 6.P  �� 6.P      G  , ,���x 0� ���x 0�@���� 0�@���� 0� ���x 0�       G  , , � 6.P � 61p �0 61p �0 6.P � 6.P      G  , ,���p 6 ���p 6@���� 6@���� 6 ���p 6       G  , ,  �� 6   �� 6@  �� 6@  �� 6   �� 6       G  , ,���P 5���P 5Š���p 5Š���p 5���P 5      G  , ,    5    5Š    5Š    5    5      G  , , �  5 �  5Š �@ 5Š �@ 5 �  5      G  , ,���h 3;����h 3?���� 3?���� 3;����h 3;�      G  , ,���x 6���x 68���� 68���� 6���x 6      G  , ,���h 0����h 0�0���� 0�0���� 0����h 0�      G  , ,���P 4U0���P 4XP���p 4XP���p 4U0���P 4U0      G  , ,���h 0|����h 0����� 0����� 0|����h 0|�      G  , ,��q� 2o@��q� 2r`��t� 2r`��t� 2o@��q� 2o@      G  , ,���X 0<����X 0?����x 0?����x 0<����X 0<�      G  , , _� 6  _� 6@ b� 6@ b� 6  _� 6       G  , ,���h 5�(���h 5�H���� 5�H���� 5�(���h 5�(      G  , ,��q� 2i ��q� 2l ��t� 2l ��t� 2i ��q� 2i       G  , , �P 6X �P 6x �p 6x �p 6X �P 6X      G  , ,���X 06����X 09����x 09����x 06����X 06�      G  , ,���x 3�����x 3������ 3������ 3�����x 3��      G  , ,��q� /� ��q� /�@��t� /�@��t� /� ��q� /�       G  , ,��_� 6@H��_� 6Ch��b� 6Ch��b� 6@H��_� 6@H      G  , , F� 6@H F� 6Ch I� 6Ch I� 6@H F� 6@H      G  , ,���P 5�@���P 5�`���p 5�`���p 5�@���P 5�@      G  , ,    5�@    5�`    5�`    5�@    5�@      G  , , �  5�@ �  5�` �@ 5�` �@ 5�@ �  5�@      G  , , F� 6: F� 6=( I� 6=( I� 6: F� 6:      G  , , � 6: � 6=( � 6=( � 6: � 6:      G  , ,  0 6  0 68 P 68 P 6  0 6      G  , ,��q� /����q� /� ��t� /� ��t� /����q� /��      G  , ,���x 3�@���x 3�`���� 3�`���� 3�@���x 3�@      G  , ,���p /i����p /l����� /l����� /i����p /i�      G  , ,���` 5�p���` 5����� 5����� 5�p���` 5�p      G  , , � 6@H � 6Ch � 6Ch � 6@H � 6@H      G  , , �P 6 �P 68 �p 68 �p 6 �P 6      G  , , �� 5�( �� 5�H �  5�H �  5�( �� 5�(      G  , ,  ZP 5�p  ZP 5�  ]p 5�  ]p 5�p  ZP 5�p      G  , , p 5�p p 5� � 5� � 5�p p 5�p      G  , ,���h 5�h���h 5������ 5������ 5�h���h 5�h      G  , , �� 5�h �� 5�� �  5�� �  5�h �� 5�h      G  , ,��q� 5.`��q� 51���t� 51���t� 5.`��q� 5.`      G  , , y  5�h y  5�� |  5�� |  5�h y  5�h      G  , ,��q� 5( ��q� 5+@��t� 5+@��t� 5( ��q� 5(       G  , ,���p 2(����p 2,���� 2,���� 2(����p 2(�      G  , ,���p 4����p 4�0���� 4�0���� 4����p 4�      G  , , y  5�( y  5�H |  5�H |  5�( y  5�(      G  , ,���p 4�����p 4������ 4������ 4�����p 4��      G  , ,���x +D����x +H ���� +H ���� +D����x +D�      G  , ,���x . ���x . ���� . ���� . ���x .       G  , ,���h +����h +����� +����� +����h +�      G  , ,��q� ,����q� ,����t� ,����t� ,����q� ,��      G  , ,���h *�����h +����� +����� *�����h *��      G  , ,���P .�����P .����p .����p .�����P .��      G  , ,���X *�����X *�����x *�����x *�����X *��      G  , ,���p ,�����p ,������ ,������ ,�����p ,��      G  , ,���X *�@���X *�`���x *�`���x *�@���X *�@      G  , ,���h -�����h -����� -����� -�����h -��      G  , ,��q� *1���q� *5 ��t� *5 ��t� *1���q� *1�      G  , ,���p ,�p���p ,������ ,������ ,�p���p ,�p      G  , ,��q� *+���q� *.���t� *.���t� *+���q� *+�      G  , ,��_� .JP��_� .Mp��b� .Mp��b� .JP��_� .JP      G  , ,���p )����p )����� )����� )����p )�      G  , ,���` ,d`���` ,g����� ,g����� ,d`���` ,d`      G  , ,���p )�P���p )�p���� )�p���� )�P���p )�P      G  , ,���h -�����h -������ -������ -�����h -��      G  , ,���` )�@���` )�`���� )�`���� )�@���` )�@      G  , ,���` ,^ ���` ,a@���� ,a@���� ,^ ���` ,^       G  , ,���` )� ���` )� ���� )� ���� )� ���` )�       G  , ,���P .�0���P .�P���p .�P���p .�0���P .�0      G  , ,���P )^����P )b���p )b���p )^����P )^�      G  , ,���P ,���P ,!0���p ,!0���p ,���P ,      G  , ,���P )X����P )[����p )[����p )X����P )X�      G  , ,���p /c����p /f����� /f����� /c����p /c�      G  , ,���X -}����X -�����x -�����x -}����X -}�      G  , ,���` /#����` /&����� /&����� /#����` /#�      G  , ,��_� (�P��_� (�p��b� (�p��b� (�P��_� (�P      G  , ,���P ,����P ,����p ,����p ,����P ,�      G  , ,��_� (���_� (�0��b� (�0��b� (���_� (�      G  , ,���x .
@���x .`���� .`���� .
@���x .
@      G  , ,��_� +�p��_� +����b� +����b� +�p��_� +�p      G  , ,���X -w`���X -z����x -z����x -w`���X -w`      G  , ,��_� +�0��_� +�P��b� +�P��b� +�0��_� +�0      G  , ,��_� .P���_� .S���b� .S���b� .P���_� .P�      G  , ,���x +K ���x +N@���� +N@���� +K ���x +K       G  , ,��q� ,� ��q� ,� ��t� ,� ��t� ,� ��q� ,�       G  , ,���` /@���` / `���� / `���� /@���` /@      G  , ,���h (?p���h (B����� (B����� (?p���h (?p      G  , ,���p !�����p !����� !����� !�����p !��      G  , ,���X %: ���X %= ���x %= ���x %: ���X %:       G  , ,���` !g����` !k ���� !k ���� !g����` !g�      G  , ,���` &�����` &� ���� &� ���� &�����` &��      G  , ,���` !a����` !d����� !d����� !a����` !a�      G  , ,��q� $����q� $����t� $����t� $����q� $��      G  , ,���P !!����P !$����p !$����p !!����P !!�      G  , ,��q� 'r���q� 'u���t� 'u���t� 'r���q� 'r�      G  , ,���P !P���P !p���p !p���p !P���P !P      G  , ,��q� $�`��q� $����t� $����t� $�`��q� $�`      G  , ,��_�  ����_�  ���b�  ���b�  ����_�  ��      G  , ,���P &�����P &�����p &�����p &�����P &��      G  , ,��_�  ����_�  ����b�  ����b�  ����_�  ��      G  , ,���p $mP���p $pp���� $pp���� $mP���p $mP      G  , ,���x  N����x  Q�����  Q�����  N����x  N�      G  , ,���h (E����h (H����� (H����� (E����h (E�      G  , ,���x  H`���x  K�����  K�����  H`���x  H`      G  , ,���p $g���p $j0���� $j0���� $g���p $g      G  , ,���h  P���h  p����  p����  P���h  P      G  , ,���P &�����P &�����p &�����p &�����P &��      G  , ,���h  ���h  0����  0����  ���h        G  , ,���` $' ���` $* ���� $* ���� $' ���` $'       G  , ,���X � ���X � ���x � ���x � ���X �       G  , ,��q� 'l���q� 'o���t� 'o���t� 'l���q� 'l�      G  , ,���X �����X �����x �����x �����X ��      G  , ,���` $ ����` $#����� $#����� $ ����` $ �      G  , ,��q� 5`��q� 8���t� 8���t� 5`��q� 5`      G  , ,��_� &0��_� &P��b� &P��b� &0��_� &0      G  , ,��q� / ��q� 2@��t� 2@��t� / ��q� /       G  , ,���P #����P #�����p #�����p #����P #�      G  , ,���p ����p �0���� �0���� ����p �      G  , ,���X '�`���X (����x (����x '�`���X '�`      G  , ,���p �����p ������ ������ �����p ��      G  , ,���P #�p���P #ݐ���p #ݐ���p #�p���P #�p      G  , ,���` �����` ������ ������ �����` ��      G  , ,��_� &���_� &��b� &��b� &���_� &�      G  , ,���` �����` ������ ������ �����` ��      G  , ,��_� #T��_� #W0��b� #W0��b� #T��_� #T      G  , ,���P bp���P e����p e����p bp���P bp      G  , ,���p ',p���p '/����� '/����� ',p���p ',p      G  , ,���P \0���P _P���p _P���p \0���P \0      G  , ,��_� #M���_� #P���b� #P���b� #M���_� #M�      G  , ,��_� ����_� ����b� ����b� ����_� ��      G  , ,���x %�����x %� ���� %� ���� %�����x %��      G  , ,��_� ϐ��_� Ұ��b� Ұ��b� ϐ��_� ϐ      G  , ,���x #����x #����� #����� #����x #�      G  , ,���x �����x ������ ������ �����x ��      G  , ,���x (�����x (������ (������ (�����x (��      G  , ,���x �@���x �`���� �`���� �@���x �@      G  , ,���x #����x #
����� #
����� #����x #�      G  , ,���h I0���h LP���� LP���� I0���h I0      G  , ,���x %Ơ���x %������ %������ %Ơ���x %Ơ      G  , ,���h B����h F���� F���� B����h B�      G  , ,���h "�p���h "ʐ���� "ʐ���� "�p���h "�p      G  , ,���X ����X  ���x  ���x ����X �      G  , ,���p '&0���p ')P���� ')P���� '&0���p '&0      G  , ,���X �����X �����x �����x �����X ��      G  , ,���h "�0���h "�P���� "�P���� "�0���h "�0      G  , ,��q� v@��q� y`��t� y`��t� v@��q� v@      G  , ,���h %�����h %������ %������ %�����h %��      G  , ,��q� p ��q� s ��t� s ��t� p ��q� p       G  , ,���X "� ���X "�@���x "�@���x "� ���X "�       G  , ,���p /����p 3���� 3���� /����p /�      G  , ,���X '� ���X '�@���x '�@���x '� ���X '�       G  , ,���p )����p ,����� ,����� )����p )�      G  , ,���X "z����X "~ ���x "~ ���x "z����X "z�      G  , ,���` ����` ������ ������ ����` �      G  , ,���h %�P���h %�p���� %�p���� %�P���h %�P      G  , ,���` �`���` ����� ����� �`���` �`      G  , ,��q� !���q� !����t� !����t� !���q� !�      G  , ,���P �P���P �p���p �p���p �P���P �P      G  , ,���` &� ���` &�@���� &�@���� &� ���` &�       G  , ,���P ����P �0���p �0���p ����P �      G  , ,��q� !�@��q� !�`��t� !�`��t� !�@��q� !�@      G  , ,��_� ���_� ���b� ���b� ���_� �      G  , ,���X %@@���X %C`���x %C`���x %@@���X %@@      G  , ,��_� p��_� ���b� ���b� p��_� p      G  , ,���p !�0���p !�P���� !�P���� !�0���p !�0      G  , ,���x �`���x Ӏ���� Ӏ���� �`���x �`      G  , ,���x � ���x �@���� �@���� � ���x �       G  , ,���h ����h �0���� �0���� ����h �      G  , ,���h �����h ������ ������ �����h ��      G  , ,���X C����X F����x F����x C����X C�      G  , ,���X =����X @����x @����x =����X =�      G  , ,��q� � ��q� �@��t� �@��t� � ��q� �       G  , ,��q� ����q� � ��t� � ��t� ����q� ��      G  , ,���p p����p s����� s����� p����p p�      G  , ,���p j����p m����� m����� j����p j�      G  , ,���` *����` -����� -����� *����` *�      G  , ,���` $@���` '`���� '`���� $@���` $@      G  , ,���P �0���P �P���p �P���p �0���P �0      G  , ,���P �����P ����p ����p �����P ��      G  , ,��_� W���_� Z���b� Z���b� W���_� W�      G  , ,��_� QP��_� Tp��b� Tp��b� QP��_� QP      G  , ,���x @���x `���� `���� @���x @      G  , ,���x  ���x  ����  ����  ���x        G  , ,���h �����h ����� ����� �����h ��      G  , ,���h İ���h ������ ������ İ���h İ      G  , ,���X �����X �����x �����x �����X ��      G  , ,���X ~`���X �����x �����x ~`���X ~`      G  , ,��q� � ��q� � ��t� � ��t� � ��q� �       G  , ,��q� ����q� ����t� ����t� ����q� ��      G  , ,���p �����p ������ ������ �����p ��      G  , ,���p �p���p ������ ������ �p���p �p      G  , ,���` k`���` n����� n����� k`���` k`      G  , ,���` e ���` h@���� h@���� e ���` e       G  , ,���P %���P (0���p (0���p %���P %      G  , ,���P ����P !����p !����p ����P �      G  , ,��_� �p��_� ����b� ����b� �p��_� �p      G  , ,��_� �0��_� �P��b� �P��b� �0��_� �0      G  , ,���x R ���x U@���� U@���� R ���x R       G  , ,���x K����x O ���� O ���� K����x K�      G  , ,���h ����h ����� ����� ����h �      G  , ,���h ����h ����� ����� ����h �      G  , ,���X ŀ���X Ƞ���x Ƞ���x ŀ���X ŀ      G  , ,���X �@���X �`���x �`���x �@���X �@      G  , ,��q� 8���q� < ��t� < ��t� 8���q� 8�      G  , ,��q� 2���q� 5���t� 5���t� 2���q� 2�      G  , ,���p ����p ������ ������ ����p �      G  , ,���p �P���p �p���� �p���� �P���p �P      G  , ,���` �@���` �`���� �`���� �@���` �@      G  , ,���` � ���` � ���� � ���� � ���` �       G  , ,���P e����P i���p i���p e����P e�      G  , ,���P _����P b����p b����p _����P _�      G  , ,��_� �P��_� �p��b� �p��b� �P��_� �P      G  , ,��_� ���_� �0��b� �0��b� ���_� �      G  , ,���x � ���x � ���� � ���� � ���x �       G  , ,���x �����x ������ ������ �����x ��      G  , ,���h L����h O����� O����� L����h L�      G  , ,���h Fp���h I����� I����� Fp���h Fp      G  , ,���X `���X 	����x 	����x `���X `      G  , ,���X   ���X @���x @���x   ���X         G  , ,��q� y���q� |���t� |���t� y���q� y�      G  , ,��q� s���q� v���t� v���t� s���q� s�      G  , ,���p 3p���p 6����� 6����� 3p���p 3p      G  , ,���p -0���p 0P���� 0P���� -0���p -0      G  , ,���` � ���` �@���� �@���� � ���` �       G  , ,���` �����` � ���� � ���� �����` ��      G  , ,���P �����P �����p �����p �����P ��      G  , ,���P �����P �����p �����p �����P ��      G  , ,��_� 0��_� P��b� P��b� 0��_� 0      G  , ,��_� ���_� ��b� ��b� ���_� �      G  , ,���x �����x � ���� � ���� �����x ��      G  , ,���x ͠���x ������ ������ ͠���x ͠      G  , ,���h �����h ������ ������ �����h ��      G  , ,���h �P���h �p���� �p���� �P���h �P      G  , ,���X G@���X J`���x J`���x G@���X G@      G  , ,���X A ���X D ���x D ���x A ���X A       G  , ,��q� ����q� ����t� ����t� ����q� ��      G  , ,��q� �`��q� ����t� ����t� �`��q� �`      G  , ,���p tP���p wp���� wp���� tP���p tP      G  , ,���p n���p q0���� q0���� n���p n      G  , ,���` . ���` 1 ���� 1 ���� . ���` .       G  , ,���` '����` *����� *����� '����` '�      G  , ,���P ����P �����p �����p ����P �      G  , ,���P �p���P ����p ����p �p���P �p      G  , ,��_� [��_� ^0��b� ^0��b� [��_� [      G  , ,��_� T���_� W���b� W���b� T���_� T�      G  , ,���x ����x ����� ����� ����x �      G  , ,���x ����x ����� ����� ����x �      G  , ,���h �p���h ѐ���� ѐ���� �p���h �p      G  , ,���h �0���h �P���� �P���� �0���h �0      G  , ,���X � ���X �@���x �@���x � ���X �       G  , ,���X �����X � ���x � ���x �����X ��      G  , ,��q� ����q� ����t� ����t� ����q� ��      G  , ,��q� �@��q� �`��t� �`��t� �@��q� �@      G  , ,���p �0���p �P���� �P���� �0���p �0      G  , ,���p �����p ����� ����� �����p ��      G  , ,���` n����` r ���� r ���� n����` n�      G  , ,���` h����` k����� k����� h����` h�      G  , ,���P (����P +����p +����p (����P (�      G  , ,���P "P���P %p���p %p���p "P���P "P      G  , ,��_� 
����_� 
���b� 
���b� 
����_� 
��      G  , ,��_� 
����_� 
����b� 
����b� 
����_� 
��      G  , ,���x 
U����x 
X����� 
X����� 
U����x 
U�      G  , ,���x 
O`���x 
R����� 
R����� 
O`���x 
O`      G  , ,���h 
P���h 
p���� 
p���� 
P���h 
P      G  , ,���h 
	���h 
0���� 
0���� 
	���h 
	      G  , ,���X 	� ���X 	� ���x 	� ���x 	� ���X 	�       G  , ,���X 	�����X 	�����x 	�����x 	�����X 	��      G  , ,��q� 	<`��q� 	?���t� 	?���t� 	<`��q� 	<`      G  , ,��q� 	6 ��q� 	9@��t� 	9@��t� 	6 ��q� 	6       G  , ,���p ����p �0���� �0���� ����p �      G  , ,���p �����p ������ ������ �����p ��      G  , ,���` �����` ������ ������ �����` ��      G  , ,���` �����` ������ ������ �����` ��      G  , ,���P ip���P l����p l����p ip���P ip      G  , ,���P c0���P fP���p fP���p c0���P c0      G  , ,��_� ����_� ����b� ����b� ����_� ��      G  , ,��_� ֐��_� ٰ��b� ٰ��b� ֐��_� ֐      G  , ,���x �����x ������ ������ �����x ��      G  , ,���x �@���x �`���� �`���� �@���x �@      G  , ,���h P0���h SP���� SP���� P0���h P0      G  , ,���h I����h M���� M���� I����h I�      G  , ,���X 	����X  ���x  ���x 	����X 	�      G  , ,���X ����X ����x ����x ����X �      G  , ,��q� }@��q� �`��t� �`��t� }@��q� }@      G  , ,��q� w ��q� z ��t� z ��t� w ��q� w       G  , ,���p 6����p :���� :���� 6����p 6�      G  , ,���p 0����p 3����� 3����� 0����p 0�      G  , ,���` ����` ������ ������ ����` �      G  , ,���` �`���` ����� ����� �`���` �`      G  , ,���P �P���P �p���p �p���p �P���P �P      G  , ,���P ����P �0���p �0���p ����P �      G  , ,��_� ���_�  ���b�  ���b� ���_� �      G  , ,��_� p��_� ���b� ���b� p��_� p      G  , ,���x �`���x ڀ���� ڀ���� �`���x �`      G  , ,���x � ���x �@���� �@���� � ���x �       G  , ,���h ����h �0���� �0���� ����h �      G  , ,���h �����h ������ ������ �����h ��      G  , ,���X J����X M����x M����x J����X J�      G  , ,���X D����X G����x G����x D����X D�      G  , ,��q� � ��q� �@��t� �@��t� � ��q� �       G  , ,��q� ����q� � ��t� � ��t� ����q� ��      G  , ,���p w����p z����� z����� w����p w�      G  , ,���p q����p t����� t����� q����p q�      G  , ,���` 1����` 4����� 4����� 1����` 1�      G  , ,���` +@���` .`���� .`���� +@���` +@      G  , ,���P �0���P �P���p �P���p �0���P �0      G  , ,���P �����P ����p ����p �����P ��      G  , ,��_� ^���_� a���b� a���b� ^���_� ^�      G  , ,��_� XP��_� [p��b� [p��b� XP��_� XP      G  , ,���x @���x `���� `���� @���x @      G  , ,���x  ���x  ����  ����  ���x        G  , ,���h �����h ����� ����� �����h ��      G  , ,���h ˰���h ������ ������ ˰���h ˰      G  , ,���X �����X �����x �����x �����X ��      G  , ,���X �`���X �����x �����x �`���X �`      G  , ,��q�  � ��q�  ��t�  ��t�  � ��q�  �       G  , ,��q�  ����q�  ����t�  ����t�  ����q�  ��      G  , ,���p  �����p  ������  ������  �����p  ��      G  , ,���p  �p���p  ������  ������  �p���p  �p      G  , ,���`  r`���`  u�����  u�����  r`���`  r`      G  , ,���`  l ���`  o@����  o@����  l ���`  l       G  , ,���P  ,���P  /0���p  /0���p  ,���P  ,      G  , ,���P  %����P  (����p  (����p  %����P  %�      G  , ,���P���`���P�������p�������p���`���P���`      G  , ,   ���`   ����   ����   ���`   ���`      G  , , � ���` � ���� �@���� �@���` � ���`      G  , ,���P��� ���P���@���p���@���p��� ���P���       G  , ,   ���    ���@   ���@   ���    ���       G  , , � ���  � ���@ �@���@ �@���  � ���       G  , ,���X���h���X������x������x���h���X���h      G  , , s����h s���� v���� v����h s����h      G  , , 2����h 2���� 5���� 5����h 2����h      G  , ,���X���(���X���H���x���H���x���(���X���(      G  , , s����( s����H v����H v����( s����(      G  , , 2����( 2����H 5����H 5����( 2����(      G  , ,���`���p���`��Ԑ������Ԑ�������p���`���p      G  , ,  ZP���p  ZP��Ԑ  ]p��Ԑ  ]p���p  ZP���p      G  , , p���p p��Ԑ ���Ԑ ����p p���p      G  , ,���`���0���`���P�������P�������0���`���0      G  , ,  ZP���0  ZP���P  ]p���P  ]p���0  ZP���0      G  , , p���0 p���P ����P ����0 p���0      G  , ,���h���x���h���������������x���h���x      G  , , �����x ���� � �� � ���x �����x      G  , , y ���x y �� | �� | ���x y ���x      G  , ,���h���8���h���X�������X�������8���h���8      G  , , �����8 �����X � ���X � ���8 �����8      G  , , y ���8 y ���X | ���X | ���8 y ���8      G  , ,���p�������p�����������������������p����      G  , ,  ������  ������  ������  ������  ������      G  , , _����� _����� b����� b����� _�����      G  , ,���p���@���p���`�������`�������@���p���@      G  , ,  �����@  �����`  �����`  �����@  �����@      G  , , _����@ _����` b����` b����@ _����@      G  , ,���x�������x�����������������������x����      G  , ,  0����  0���� P���� P����  0����      G  , , �P���� �P���� �p���� �p���� �P����      G  , ,���x���H���x���h�������h�������H���x���H      G  , ,  0���H  0���h P���h P���H  0���H      G  , , �P���H �P���h �p���h �p���H �P���H      G  , ,��q�������q�������t�������t�������q�����      G  , ,  ������  ������  �����  �����  ������      G  , , ����� ����� �0���� �0���� �����      G  , ,��q����P��q����p��t����p��t����P��q����P      G  , ,  �����P  �����p  ����p  ����P  �����P      G  , , ����P ����p �0���p �0���P ����P      G  , ,��_���w���_���z���b���z���b���w���_���w�      G  , , F���w� F���z� I���z� I���w� F���w�      G  , , ���w� ���z� ���z� ���w� ���w�      G  , ,��_���qX��_���tx��b���tx��b���qX��_���qX      G  , , F���qX F���tx I���tx I���qX F���qX      G  , , ���qX ���tx ���tx ���qX ���qX      G  , , ����@ ����` " ���` " ���@ ����@      G  , , � ���@ � ���` � ���` � ���@ � ���@      G  , , �����( �����H �����H �����( �����(      G  , , 	�����( 	�����H 	����H 	����( 	�����(      G  , , �@���  �@���@ �`���@ �`���  �@���       G  , , ~p���� ~p���� ������ ������ ~p����      G  , , 
=����� 
=����� 
@����� 
@����� 
=�����      G  , , 8 ���x 8 �� ;@�� ;@���x 8 ���x      G  , , 	�@���x 	�@�� 	�`�� 	�`���x 	�@���x      G  , , �����h ����� ����� �����h �����h      G  , , ~p���H ~p���h �����h �����H ~p���H      G  , , 
=����H 
=����h 
@����h 
@����H 
=����H      G  , , 	�����h 	����� 	���� 	����h 	�����h      G  , , ؐ���p ؐ��Ԑ ۰��Ԑ ۰���p ؐ���p      G  , , 8 ���8 8 ���X ;@���X ;@���8 8 ���8      G  , , e0���� e0���� hP���� hP���� e0����      G  , , 	$P���� 	$P���� 	'p���� 	'p���� 	$P����      G  , , 	�@���8 	�@���X 	�`���X 	�`���8 	�@���8      G  , , �����p ����Ԑ ����Ԑ �����p �����p      G  , , Q`���  Q`���@ T����@ T����  Q`���       G  , , e0���P e0���p hP���p hP���P e0���P      G  , , 	$P���P 	$P���p 	'p���p 	'p���P 	$P���P      G  , , Q`���` Q`���� T����� T����` Q`���`      G  , , ����� ����� " ���� " ���� �����      G  , , � ���� � ���� � ���� � ���� � ����      G  , , ����w� ����z� ����z� ����w� ����w�      G  , , 
����w� 
����z� 
� ��z� 
� ��w� 
����w�      G  , , �@���` �@���� �`���� �`���` �@���`      G  , , ؐ���0 ؐ���P ۰���P ۰���0 ؐ���0      G  , , �����0 �����P �����P �����0 �����0      G  , , ����qX ����tx ����tx ����qX ����qX      G  , , 
����qX 
����tx 
� ��tx 
� ��qX 
����qX      G  , , \@���� \@���� _`���� _`���� \@����      G  , , `���� `���� ����� ����� `����      G  , , ڀ���� ڀ���� ݠ���� ݠ���� ڀ����      G  , , ����p ���Ԑ �0��Ԑ �0���p ����p      G  , , �0���p �0��Ԑ �P��Ԑ �P���p �0���p      G  , , p���h p��� s0��� s0���h p���h      G  , , /0���h /0��� 2P��� 2P���h /0���h      G  , , �P���h �P��� �p��� �p���h �P���h      G  , , � ���@ � ���` �@���` �@���@ � ���@      G  , , \@���@ \@���` _`���` _`���@ \@���@      G  , , `���@ `���` ����` ����@ `���@      G  , , ڀ���@ ڀ���` ݠ���` ݠ���@ ڀ���@      G  , , �p���h �p��� ����� �����h �p���h      G  , , ����  ����@ ����@ ����  ����       G  , , V����0 V����P Y����P Y����0 V����0      G  , , ����0 ����P ���P ���0 ����0      G  , , ����0 ����P �0���P �0���0 ����0      G  , , ������ ������ ������ ������ ������      G  , , ������ ������ ������ ������ ������      G  , , z����� z����� ~���� ~���� z�����      G  , , :���� :���� =0���� =0���� :����      G  , , �0���0 �0���P �P���P �P���0 �0���0      G  , , Ϡ���  Ϡ���@ �����@ �����  Ϡ���       G  , , �����  �����@ �����@ �����  �����       G  , , M����  M����@ Q ���@ Q ���  M����       G  , ,  ���   ���@  ���@  ���   ���       G  , , �����H �����h �����h �����H �����H      G  , , �����H �����h �����h �����H �����H      G  , , z����H z����h ~���h ~���H z����H      G  , , :���H :���h =0���h =0���H :���H      G  , , p���( p���H s0���H s0���( p���(      G  , , �`���x �`�� ���� �����x �`���x      G  , , u����x u��� x��� x����x u����x      G  , , 4����x 4��� 7��� 7����x 4����x      G  , , �����x ���� ���� �����x �����x      G  , , �p���� �p���� ����� ����� �p����      G  , , ������ ������ ������ ������ ������      G  , , a����� a����� d����� d����� a�����      G  , ,  �����  ����� #����� #�����  �����      G  , , /0���( /0���H 2P���H 2P���( /0���(      G  , , �P���( �P���H �p���H �p���( �P���(      G  , , �p���( �p���H �����H �����( �p���(      G  , , ����` ����� ����� ����` ����`      G  , , Ϡ���` Ϡ���� ������ �����` Ϡ���`      G  , , �p���P �p���p ����p ����P �p���P      G  , , �����P �����p �����p �����P �����P      G  , , a����P a����p d����p d����P a����P      G  , ,  ����P  ����p #����p #����P  ����P      G  , , �`���8 �`���X �����X �����8 �`���8      G  , , u����8 u����X x����X x����8 u����8      G  , , 4����8 4����X 7����X 7����8 4����8      G  , , �����8 �����X �����X �����8 �����8      G  , , �����` ������ ������ �����` �����`      G  , , C ��w� C ��z� F ��z� F ��w� C ��w�      G  , ,  ��w�  ��z� @��z� @��w�  ��w�      G  , , �@��w� �@��z� �`��z� �`��w� �@��w�      G  , , �`��w� �`��z� ����z� ����w� �`��w�      G  , , M����` M����� Q ���� Q ���` M����`      G  , ,  ���`  ����  ����  ���`  ���`      G  , , V����p V���Ԑ Y���Ԑ Y����p V����p      G  , , ����p ���Ԑ ��Ԑ ���p ����p      G  , , � ���� � ���� �@���� �@���� � ����      G  , , C ��qX C ��tx F ��tx F ��qX C ��qX      G  , ,  ��qX  ��tx @��tx @��qX  ��qX      G  , , �@��qX �@��tx �`��tx �`��qX �@��qX      G  , , �`��qX �`��tx ����tx ����qX �`��qX      G  , , ,�4 j� ,�4 m� ,�T m� ,�T j� ,�4 j�      G  , , ,�T � ,�T �� ,�t �� ,�t � ,�T �      G  , , -$ 8� -$ <  -D <  -D 8� -$ 8�      G  , , ,�T �p ,�T � ,�t � ,�t �p ,�T �p      G  , , ,�< İ ,�< �� ,�\ �� ,�\ İ ,�< İ      G  , , -* [ -* ^0 --< ^0 --< [ -* [      G  , , -$ 2� -$ 5� -D 5� -D 2� -$ 2�      G  , , -* T� -* W� --< W� --< T� -* T�      G  , , ,�< � ,�< �0 ,�\ �0 ,�\ � ,�< �      G  , , ,�4 � ,�4 �� ,�T �� ,�T � ,�4 �      G  , , ,�L �� ,�L �� ,�l �� ,�l �� ,�L ��      G  , , ,�4 �P ,�4 �p ,�T �p ,�T �P ,�4 �P      G  , , ,�D *� ,�D -� ,�d -� ,�d *� ,�D *�      G  , , ,�D �@ ,�D �` ,�d �` ,�d �@ ,�D �@      G  , , ,�L ~` ,�L �� ,�l �� ,�l ~` ,�L ~`      G  , , ,�D �  ,�D �  ,�d �  ,�d �  ,�D �       G  , , ,�L =� ,�L @� ,�l @� ,�l =� ,�L =�      G  , , ,�T e� ,�T i ,�t i ,�t e� ,�T e�      G  , , -$ �  -$ �  -D �  -D �  -$ �       G  , , ,�T _� ,�T b� ,�t b� ,�t _� ,�T _�      G  , , ,�D $@ ,�D '` ,�d '` ,�d $@ ,�D $@      G  , , -* �P -* �p --< �p --< �P -* �P      G  , , -$ �� -$ �� -D �� -D �� -$ ��      G  , , -* � -* �0 --< �0 --< � -* �      G  , , -, �  -, �@ -	L �@ -	L �  -, �       G  , , -, �  -, �  -	L �  -	L �  -, �       G  , , ,�4 �� ,�4 �� ,�T �� ,�T �� ,�4 ��      G  , , -, �� -, �� -	L �� -	L �� -, ��      G  , , ,�T �0 ,�T �P ,�t �P ,�t �0 ,�T �0      G  , , ,�< L� ,�< O� ,�\ O� ,�\ L� ,�< L�      G  , , ,�4 �p ,�4 �� ,�T �� ,�T �p ,�4 �p      G  , , ,�< Fp ,�< I� ,�\ I� ,�\ Fp ,�< Fp      G  , , -$ �  -$ �@ -D �@ -D �  -$ �       G  , , ,�L ` ,�L 	� ,�l 	� ,�l ` ,�L `      G  , , ,�D k` ,�D n� ,�d n� ,�d k` ,�D k`      G  , , ,�L    ,�L @ ,�l @ ,�l    ,�L         G  , , ,�T �� ,�T � ,�t � ,�t �� ,�T ��      G  , , -$ y� -$ |� -D |� -D y� -$ y�      G  , , ,�D e  ,�D h@ ,�d h@ ,�d e  ,�D e       G  , , -$ s� -$ v� -D v� -D s� -$ s�      G  , , ,�< �� ,�< �� ,�\ �� ,�\ �� ,�< ��      G  , , ,�4 3p ,�4 6� ,�T 6� ,�T 3p ,�4 3p      G  , , ,�T % ,�T (0 ,�t (0 ,�t % ,�T %      G  , , ,�4 -0 ,�4 0P ,�T 0P ,�T -0 ,�4 -0      G  , , -* W� -* Z� --< Z� --< W� -* W�      G  , , ,�D �  ,�D �@ ,�d �@ ,�d �  ,�D �       G  , , ,�T � ,�T !� ,�t !� ,�t � ,�T �      G  , , ,�D �� ,�D �  ,�d �  ,�d �� ,�D ��      G  , , -$ �� -$ �  -D �  -D �� -$ ��      G  , , ,�T �� ,�T �� ,�t �� ,�t �� ,�T ��      G  , , -* �p -* �� --< �� --< �p -* �p      G  , , ,�T �� ,�T �� ,�t �� ,�t �� ,�T ��      G  , , -* QP -* Tp --< Tp --< QP -* QP      G  , , -* 0 -* P --< P --< 0 -* 0      G  , , -* �0 -* �P --< �P --< �0 -* �0      G  , , -* � -*  --<  --< � -* �      G  , , -, �` -, Ӏ -	L Ӏ -	L �` -, �`      G  , , -, �� -, �  -	L �  -	L �� -, ��      G  , , -, R  -, U@ -	L U@ -	L R  -, R       G  , , -, ͠ -, �� -	L �� -	L ͠ -, ͠      G  , , -, @ -, ` -	L ` -	L @ -, @      G  , , ,�< �� ,�< �� ,�\ �� ,�\ �� ,�< ��      G  , , -, K� -, O  -	L O  -	L K� -, K�      G  , , ,�< �P ,�< �p ,�\ �p ,�\ �P ,�< �P      G  , , ,�4 p� ,�4 s� ,�T s� ,�T p� ,�4 p�      G  , , ,�L G@ ,�L J` ,�l J` ,�l G@ ,�L G@      G  , , ,�< � ,�< � ,�\ � ,�\ � ,�< �      G  , , ,�L A  ,�L D  ,�l D  ,�l A  ,�L A       G  , , -,   -,   -	L   -	L   -,        G  , , -$ �� -$ �� -D �� -D �� -$ ��      G  , , ,�< � ,�< � ,�\ � ,�\ � ,�< �      G  , , -$ �` -$ �� -D �� -D �` -$ �`      G  , , ,�L C� ,�L F� ,�l F� ,�l C� ,�L C�      G  , , ,�4 tP ,�4 wp ,�T wp ,�T tP ,�4 tP      G  , , ,�L ŀ ,�L Ƞ ,�l Ƞ ,�l ŀ ,�L ŀ      G  , , ,�4 n ,�4 q0 ,�T q0 ,�T n ,�4 n      G  , , ,�< �� ,�< � ,�\ � ,�\ �� ,�< ��      G  , , ,�D .  ,�D 1  ,�d 1  ,�d .  ,�D .       G  , , ,�L �@ ,�L �` ,�l �` ,�l �@ ,�L �@      G  , , ,�D '� ,�D *� ,�d *� ,�d '� ,�D '�      G  , , l����h l���� o���� o����h l����h      G  , , SP���p SP��Ԑ Vp��Ԑ Vp���p SP���p      G  , , p���p p��Ԑ ���Ԑ ����p p���p      G  , , ������ ������ ������ ������ ������      G  , , X����� X����� [����� [����� X�����      G  , , ����� �����  ����  ���� �����      G  , , � ���� � ���� � ���� � ���� � ����      G  , , !� ���� !� ���� !�@���� !�@���� !� ����      G  , , ѐ���p ѐ��Ԑ ԰��Ԑ ԰���p ѐ���p      G  , , �����p ����Ԑ ����Ԑ �����p �����p      G  , , !O����p !O���Ԑ !R���Ԑ !R����p !O����p      G  , , +����h +���� .���� .����h +����h      G  , , �����@ �����` �����` �����@ �����@      G  , , X����@ X����` [����` [����@ X����@      G  , , ����@ ����`  ���`  ���@ ����@      G  , , � ���@ � ���` � ���` � ���@ � ���@      G  , , !� ���@ !� ���` !�@���` !�@���@ !� ���@      G  , , �����h ����� ����� �����h �����h      G  , , �����h ����� ���� ����h �����h      G  , , �@���  �@���@ �`���@ �`���  �@���       G  , , SP���0 SP���P Vp���P Vp���0 SP���0      G  , , p���0 p���P ����P ����0 p���0      G  , , �0���� �0���� �P���� �P���� �0����      G  , , �P���� �P���� �p���� �p���� �P����      G  , , wp���� wp���� z����� z����� wp����      G  , ,  6�����  6�����  9�����  9�����  6�����      G  , , ѐ���0 ѐ���P ԰���P ԰���0 ѐ���0      G  , , �����0 �����P �����P �����0 �����0      G  , , !O����0 !O����P !R����P !R����0 !O����0      G  , , J`���  J`���@ M����@ M����  J`���       G  , , �0���H �0���h �P���h �P���H �0���H      G  , , �P���H �P���h �p���h �p���H �P���H      G  , , wp���H wp���h z����h z����H wp���H      G  , ,  6����H  6����h  9����h  9����H  6����H      G  , , !	����  !	����@ !����@ !����  !	����       G  , , �@���` �@���� �`���� �`���` �@���`      G  , , l����( l����H o����H o����( l����(      G  , , +����( +����H .����H .����( +����(      G  , , �����x ���� � �� � ���x �����x      G  , , ������ ������ ����� ����� ������      G  , , ����� ����� �0���� �0���� �����      G  , , ^0���� ^0���� aP���� aP���� ^0����      G  , , P���� P����  p����  p���� P����      G  , , r ���x r �� u �� u ���x r ���x      G  , , 1 ���x 1 �� 4@�� 4@���x 1 ���x      G  , , �@���x �@�� �`�� �`���x �@���x      G  , , �����( �����H �����H �����( �����(      G  , , �����P �����p ����p ����P �����P      G  , , ����P ����p �0���p �0���P ����P      G  , , ^0���P ^0���p aP���p aP���P ^0���P      G  , , P���P P���p  p���p  p���P P���P      G  , , �����( �����H ����H ����( �����(      G  , , J`���` J`���� M����� M����` J`���`      G  , , !	����` !	����� !����� !����` !	����`      G  , , �����8 �����X � ���X � ���8 �����8      G  , , r ���8 r ���X u ���X u ���8 r ���8      G  , , ?���w� ?���z� B���z� B���w� ?���w�      G  , , ����w� ����z� ���z� ���w� ����w�      G  , , ����w� ����z� ����z� ����w� ����w�      G  , ,  |���w�  |���z�  � ��z�  � ��w�  |���w�      G  , , 1 ���8 1 ���X 4@���X 4@���8 1 ���8      G  , , �@���8 �@���X �`���X �`���8 �@���8      G  , , � ���` � ���� �@���� �@���` � ���`      G  , , � ���  � ���@ �@���@ �@���  � ���       G  , , ?���qX ?���tx B���tx B���qX ?���qX      G  , , ����qX ����tx ���tx ���qX ����qX      G  , , ����qX ����tx ����tx ����qX ����qX      G  , ,  |���qX  |���tx  � ��tx  � ��qX  |���qX      G  , , ,�< P0 ,�< SP ,�\ SP ,�\ P0 ,�< P0      G  , , -$ �� -$ �� -D �� -D �� -$ ��      G  , , ,�< I� ,�< M ,�\ M ,�\ I� ,�< I�      G  , , -, 
U� -, 
X� -	L 
X� -	L 
U� -, 
U�      G  , , ,�< �p ,�< ѐ ,�\ ѐ ,�\ �p ,�< �p      G  , , -, 
O` -, 
R� -	L 
R� -	L 
O` -, 
O`      G  , , -$ �@ -$ �` -D �` -D �@ -$ �@      G  , , ,�L 	� ,�L   ,�l   ,�l 	� ,�L 	�      G  , , ,�4 �0 ,�4 �P ,�T �P ,�T �0 ,�4 �0      G  , , ,�L � ,�L � ,�l � ,�l � ,�L �      G  , , ,�< �0 ,�< �P ,�\ �P ,�\ �0 ,�< �0      G  , , -$ }@ -$ �` -D �` -D }@ -$ }@      G  , , -$ w  -$ z  -D z  -D w  -$ w       G  , , ,�< 
P ,�< 
p ,�\ 
p ,�\ 
P ,�< 
P      G  , , ,�< 
	 ,�< 
0 ,�\ 
0 ,�\ 
	 ,�< 
	      G  , , ,�L 	�  ,�L 	�  ,�l 	�  ,�l 	�  ,�L 	�       G  , , ,�L 	�� ,�L 	�� ,�l 	�� ,�l 	�� ,�L 	��      G  , , -, � -, � -	L � -	L � -, �      G  , , ,�4 �� ,�4 � ,�T � ,�T �� ,�4 ��      G  , , -$ 	<` -$ 	?� -D 	?� -D 	<` -$ 	<`      G  , , -$ 	6  -$ 	9@ -D 	9@ -D 	6  -$ 	6       G  , , ,�D n� ,�D r  ,�d r  ,�d n� ,�D n�      G  , , ,�4 � ,�4 �0 ,�T �0 ,�T � ,�4 �      G  , , ,�4 �� ,�4 �� ,�T �� ,�T �� ,�4 ��      G  , , ,�D h� ,�D k� ,�d k� ,�d h� ,�D h�      G  , , ,�D �� ,�D �� ,�d �� ,�d �� ,�D ��      G  , , ,�T (� ,�T +� ,�t +� ,�t (� ,�T (�      G  , , ,�L �  ,�L �@ ,�l �@ ,�l �  ,�L �       G  , , ,�D �� ,�D �� ,�d �� ,�d �� ,�D ��      G  , , -, � -, � -	L � -	L � -, �      G  , , ,�T ip ,�T l� ,�t l� ,�t ip ,�T ip      G  , , ,�T c0 ,�T fP ,�t fP ,�t c0 ,�T c0      G  , , -* �� -* �� --< �� --< �� -* ��      G  , , ,�T "P ,�T %p ,�t %p ,�t "P ,�T "P      G  , , ,�L �� ,�L �  ,�l �  ,�l �� ,�L ��      G  , , -* ֐ -* ٰ --< ٰ --< ֐ -* ֐      G  , , -* 
�� -* 
� --< 
� --< 
�� -* 
��      G  , , -, �� -, �� -	L �� -	L �� -, ��      G  , , -, �@ -, �` -	L �` -	L �@ -, �@      G  , , -* 
�� -* 
�� --< 
�� --< 
�� -* 
��      G  , , &�����  &�����@ &�����@ &�����  &�����       G  , , $U@���@ $U@���` $X`���` $X`���@ $U@���@      G  , , "�����H "�����h "�����h "�����H "�����H      G  , , %�����H %�����h %�����h %�����H %�����H      G  , , '`���@ '`���` '����` '����@ '`���@      G  , , $����0 $����P $���P $���0 $����0      G  , , &����0 &����P &�0���P &�0���0 &����0      G  , , !�p���� !�p���� !ߐ���� !ߐ���� !�p����      G  , , $������ $������ $������ $������ $������      G  , , 'Z����� 'Z����� ']����� ']����� 'Z�����      G  , , "�`���8 "�`���X "�����X "�����8 "�`���8      G  , , $U@���� $U@���� $X`���� $X`���� $U@����      G  , , $����p $���Ԑ $��Ԑ $���p $����p      G  , , &����p &���Ԑ &�0��Ԑ &�0���p &����p      G  , , "i���h "i��� "l0��� "l0���h "i���h      G  , , '`���� '`���� '����� '����� '`����      G  , , %(0���h %(0��� %+P��� %+P���h %(0���h      G  , , !�p���P !�p���p !ߐ���p !ߐ���P !�p���P      G  , , $�����P $�����p $�����p $�����P $�����P      G  , , 'Z����P 'Z����p ']����p ']����P 'Z����P      G  , , "������ "������ "������ "������ "������      G  , , %������ %������ %������ %������ %������      G  , , #Ƞ���` #Ƞ���� #������ #�����` #Ƞ���`      G  , , "�`���x "�`�� "���� "�����x "�`���x      G  , , %n����x %n��� %q��� %q����x %n����x      G  , , #< ��w� #< ��z� #? ��z� #? ��w� #< ��w�      G  , , %� ��w� %� ��z� %�@��z� %�@��w� %� ��w�      G  , , "i���( "i���H "l0���H "l0���( "i���(      G  , , %n����8 %n����X %q����X %q����8 %n����8      G  , , #Ƞ���  #Ƞ���@ #�����@ #�����  #Ƞ���       G  , , &�����` &������ &������ &�����` &�����`      G  , , %(0���( %(0���H %+P���H %+P���( %(0���(      G  , , #< ��qX #< ��tx #? ��tx #? ��qX #< ��qX      G  , , %� ��qX %� ��tx %�@��tx %�@��qX %� ��qX      G  , , ,�L D� ,�L G� ,�l G� ,�l D� ,�L D�      G  , , ,�T �P ,�T �p ,�t �p ,�t �P ,�T �P      G  , , *�p���( *�p���H *�����H *�����( *�p���(      G  , , ,�L���( ,�L���H ,�l���H ,�l���( ,�L���(      G  , , ,�4  �p ,�4  �� ,�T  �� ,�T  �p ,�4  �p      G  , , )F����  )F����@ )J ���@ )J ���  )F����       G  , , , ���  , ���@ ,	 ���@ ,	 ���  , ���       G  , , (s����H (s����h (w���h (w���H (s����H      G  , , +3���H +3���h +60���h +60���H +3���H      G  , , -,���H -,���h -	L���h -	L���H -,���H      G  , , )F����` )F����� )J ���� )J ���` )F����`      G  , , -$ �  -$ �@ -D �@ -D �  -$ �       G  , , (-����8 (-����X (0����X (0����8 (-����8      G  , , -$ �� -$ �  -D �  -D �� -$ ��      G  , , , ���` , ���� ,	 ���� ,	 ���` , ���`      G  , , ,�4 w� ,�4 z� ,�T z� ,�T w� ,�4 w�      G  , , ,�T���` ,�T���� ,�t���� ,�t���` ,�T���`      G  , , ,�4 q� ,�4 t� ,�T t� ,�T q� ,�4 q�      G  , , ,�T  , ,�T  /0 ,�t  /0 ,�t  , ,�T  ,      G  , , *�����8 *�����X *�����X *�����8 *�����8      G  , , )Ӏ���@ )Ӏ���` )֠���` )֠���@ )Ӏ���@      G  , , )�0���0 )�0���P )�P���P )�P���0 )�0���0      G  , , ,LP���0 ,LP���P ,Op���P ,Op���0 ,LP���0      G  , , ,�4���@ ,�4���` ,�T���` ,�T���@ ,�4���@      G  , , ,�T���  ,�T���@ ,�t���@ ,�t���  ,�T���       G  , , ,�T � ,�T �0 ,�t �0 ,�t � ,�T �      G  , , *����� *����� *����� *����� *�����      G  , , -$���� -$���� -D���� -D���� -$����      G  , , ,�D 1� ,�D 4� ,�d 4� ,�d 1� ,�D 1�      G  , , ,�D���0 ,�D���P ,�d���P ,�d���0 ,�D���0      G  , , ,�D +@ ,�D .` ,�d .` ,�d +@ ,�D +@      G  , , ,�<���8 ,�<���X ,�\���X ,�\���8 ,�<���8      G  , , ,�T �0 ,�T �P ,�t �P ,�t �0 ,�T �0      G  , , -* � -*  � --<  � --< � -* �      G  , , ,�T �� ,�T � ,�t � ,�t �� ,�T ��      G  , , )Ӏ���� )Ӏ���� )֠���� )֠���� )Ӏ����      G  , , -* ^� -* a� --< a� --< ^� -* ^�      G  , , -* p -* � --< � --< p -* p      G  , , ,�4���� ,�4���� ,�T���� ,�T���� ,�4����      G  , , -, �` -, ڀ -	L ڀ -	L �` -, �`      G  , , ,�4 6� ,�4 : ,�T : ,�T 6� ,�4 6�      G  , , )�0���p )�0��Ԑ )�P��Ԑ )�P���p )�0���p      G  , , ,LP���p ,LP��Ԑ ,Op��Ԑ ,Op���p ,LP���p      G  , , ,�D���p ,�D��Ԑ ,�d��Ԑ ,�d���p ,�D���p      G  , , *����P *����p *����p *����P *����P      G  , , -$���P -$���p -D���p -D���P -$���P      G  , , ,�D  l  ,�D  o@ ,�d  o@ ,�d  l  ,�D  l       G  , , -* XP -* [p --< [p --< XP -* XP      G  , , '�P���h '�P��� '�p��� '�p���h '�P���h      G  , , -, @ -, ` -	L ` -	L @ -, @      G  , , *�p���h *�p��� *����� *�����h *�p���h      G  , , -,   -,   -	L   -	L   -,        G  , , ,�L���h ,�L��� ,�l��� ,�l���h ,�L���h      G  , , ,�< �� ,�< � ,�\ � ,�\ �� ,�< ��      G  , , ,�4 0� ,�4 3� ,�T 3� ,�T 0� ,�4 0�      G  , , ,�T  %� ,�T  (� ,�t  (� ,�t  %� ,�T  %�      G  , , (s����� (s����� (w���� (w���� (s�����      G  , , +3���� +3���� +60���� +60���� +3����      G  , , (-����x (-��� (0��� (0����x (-����x      G  , , -,���� -,���� -	L���� -	L���� -,����      G  , , -, �  -, �@ -	L �@ -	L �  -, �       G  , , (�@��w� (�@��z� (�`��z� (�`��w� (�@��w�      G  , , +y`��w� +y`��z� +|���z� +|���w� +y`��w�      G  , , -*��w� -*��z� --<��z� --<��w� -*��w�      G  , , ,�< ˰ ,�< �� ,�\ �� ,�\ ˰ ,�< ˰      G  , , *�����x *���� *���� *�����x *�����x      G  , , ,�L �� ,�L �� ,�l �� ,�l �� ,�L ��      G  , , ,�<���x ,�<�� ,�\�� ,�\���x ,�<���x      G  , , ,�L �` ,�L �� ,�l �� ,�l �` ,�L �`      G  , , ,�D � ,�D �� ,�d �� ,�d � ,�D �      G  , , -$  �  -$   -D   -D  �  -$  �       G  , , ,�< � ,�< �0 ,�\ �0 ,�\ � ,�< �      G  , , -$  �� -$  �� -D  �� -D  �� -$  ��      G  , , ,�4  �� ,�4  �� ,�T  �� ,�T  �� ,�4  ��      G  , , ,�D  r` ,�D  u� ,�d  u� ,�d  r` ,�D  r`      G  , , ,�< �� ,�< �� ,�\ �� ,�\ �� ,�< ��      G  , , ,�D �` ,�D � ,�d � ,�d �` ,�D �`      G  , , ,�L J� ,�L M� ,�l M� ,�l J� ,�L J�      G  , , '�P���( '�P���H '�p���H '�p���( '�P���(      G  , , (�@��qX (�@��tx (�`��tx (�`��qX (�@��qX      G  , , +y`��qX +y`��tx +|���tx +|���qX +y`��qX      G  , , -*��qX -*��tx --<��tx --<��qX -*��qX   	   H   !       $ ,�0 �� +�. �� +�. �� +�� ��      H   ,��[< 68���[< 6D� -1� 6D� -1� 68���[< 68�      H   ,��m4 6&���m4 62� -� 62� -� 6&���m4 6&�      H   ,��, 6���, 6 � -� 6 � -� 6���, 6�      H   ,���$ 6����$ 6� ,�� 6� ,�� 6����$ 6�      H   ,��� 5����� 5�� ,� 5�� ,� 5����� 5��      H   ,��� 5���� 5� ,װ 5� ,װ 5���� 5�      H   ,��� 5���� 5�� ,Ÿ 5�� ,Ÿ 5���� 5�      H   ,��� 5���� 5�� ,�� 5�� ,�� 5���� 5�      H   ,�������������� ,������ ,�������������      H   ,������������� ,Ÿ��� ,Ÿ�����������      H   ,�����������ռ ,װ��ռ ,װ���������      H   ,������������� ,����� ,����������      H   ,���$������$���� ,������ ,��������$���      H   ,��,�����,���� -����� -������,���      H   ,��m4���$��m4���� -����� -����$��m4���$      H   ,��[<��p,��[<��{� -1���{� -1���p,��[<��p,      H   , ,�� (�� ,�� (�L -� (�L -� (�� ,�� (��      H   , ,�� /bd ,�� /n -� /n -� /bd ,�� /bd      H   , -%� 68� -%� 68� -1� 68� -1� 68� -%� 68�      H   , *� 62� *� 62� *!< 62� *!< 62� *� 62�      H   , -� 62� -� 62� -� 62� -� 62� -� 62�      H   , *� 6&� *� 6&� *!< 6&� *!< 6&� *� 6&�      H   , -� 6&� -� 6&� -� 6&� -� 6&� -� 6&�      H   , (o� 6 � (o� 6 � ({\ 6 � ({\ 6 � (o� 6 �      H   , +.� 6 � +.� 6 � +:| 6 � +:| 6 � +.� 6 �      H   , -� 6 � -� 6 � -� 6 � -� 6 � -� 6 �      H   , (o� 6� (o� 6� ({\ 6� ({\ 6� (o� 6�      H   , +.� 6� +.� 6� +:| 6� +:| 6� +.� 6�      H   , -� 6� -� 6� -� 6� -� 6� -� 6�      H   , )�4 6� )�4 6� )�� 6� )�� 6� )�4 6�      H   , ,�� 6� ,�� 6� ,�� 6� ,�� 6� ,�� 6�      H   , )�4 6� )�4 6� )�� 6� )�� 6� )�4 6�      H   , ,�� 6� ,�� 6� ,�� 6� ,�� 6� ,�� 6�      H   , ()T 5�� ()T 5�� (5 5�� (5 5�� ()T 5��      H   , *�t 5�� *�t 5�� *�, 5�� *�, 5�� *�t 5��      H   , ,�� 5�� ,�� 5�� ,� 5�� ,� 5�� ,�� 5��      H   , ()T 5�� ()T 5�� (5 5�� (5 5�� ()T 5��      H   , *�t 5�� *�t 5�� *�, 5�� *�, 5�� *�t 5��      H   , ,�� 5�� ,�� 5�� ,� 5�� ,� 5�� ,�� 5��      H   , )�� 5� )�� 5�� )�� 5�� )�� 5� )�� 5�      H   , ,H 5� ,H 5�� ,S� 5�� ,S� 5� ,H 5�      H   , ,�� 5� ,�� 5�� ,װ 5�� ,װ 5� ,�� 5�      H   , )�� 5�� )�� 5� )�� 5� )�� 5�� )�� 5��      H   , ,H 5�� ,H 5� ,S� 5� ,S� 5�� ,H 5��      H   , ,�� 5�� ,�� 5� ,װ 5� ,װ 5�� ,�� 5��      H   , '� 5�� '� 5�� '� 5�� '� 5�� '� 5��      H   , *�$ 5�� *�$ 5�� *�� 5�� *�� 5�� *�$ 5��      H   , ,�  5�� ,�  5�� ,Ÿ 5�� ,Ÿ 5�� ,�  5��      H   , (�� 6D� (�� 6D� (�� 6D� (�� 6D� (�� 6D�      H   , '� 5� '� 5� '� 5� '� 5� '� 5�      H   , *�$ 5� *�$ 5� *�� 5� *�� 5� *�$ 5�      H   , ,�  5� ,�  5� ,Ÿ 5� ,Ÿ 5� ,�  5�      H   , )B� 5�� )B� 5�� )NL 5�� )NL 5�� )B� 5��      H   , ,� 5�� ,� 5�� ,l 5�� ,l 5�� ,� 5��      H   , ,� 5�� ,� 5�� ,�� 5�� ,�� 5�� ,� 5��      H   , +u 6D� +u 6D� +�� 6D� +�� 6D� +u 6D�      H   , )B� 5�
 )B� 5� )NL 5� )NL 5�
 )B� 5�
      H   , ,� 5�
 ,� 5� ,l 5� ,l 5�
 ,� 5�
      H   , ,� 5�
 ,� 5� ,�� 5� ,�� 5�
 ,� 5�
      H   , -� 52� -� 52� -� 52� -� 52� -� 52�      H   , ,�� 5&� ,�� 52� -1� 52� -1� 5&� ,�� 5&�      H   , -� 5&� -� 5&� -� 5&� -� 5&� -� 5&�      H   , ,�� 4�\ ,�� 4�f ,�� 4�f ,�� 4�\ ,�� 4�\      H   , ,�� 4� ,�� 4�\ -� 4�\ -� 4� ,�� 4�      H   , ,�� 4�� ,�� 4� ,�� 4� ,�� 4�� ,�� 4��      H   , ,�� 4� ,�� 4� ,װ 4� ,װ 4� ,�� 4�      H   , ,�� 4�T ,�� 4� ,� 4� ,� 4�T ,�� 4�T      H   , ,�� 4�J ,�� 4�T ,װ 4�T ,װ 4�J ,�� 4�J      H   , ,� 4_� ,� 4_� ,�� 4_� ,�� 4_� ,� 4_�      H   , ,�� 4T ,�� 4_� ,Ÿ 4_� ,Ÿ 4T ,�� 4T      H   , ,� 4S� ,� 4T ,�� 4T ,�� 4S� ,� 4S�      H   , -%� 3� -%� 3�& -1� 3�& -1� 3� -%� 3�      H   , ,�� 3�d ,�� 3� -1� 3� -1� 3�d ,�� 3�d      H   , -%� 3�Z -%� 3�d -1� 3�d -1� 3�Z -%� 3�Z      H   , -� 3�� -� 3�� -� 3�� -� 3�� -� 3��      H   , ,�� 3� ,�� 3�� -� 3�� -� 3� ,�� 3�      H   , -� 3�
 -� 3� -� 3� -� 3�
 -� 3�
      H   , ,�� 3F| ,�� 3F� ,� 3F� ,� 3F| ,�� 3F|      H   , ,�� 3:� ,�� 3F| ,� 3F| ,� 3:� ,�� 3:�      H   , ,�� 3:� ,�� 3:� ,� 3:� ,� 3:� ,�� 3:�      H   , ,�  3 , ,�  3 6 ,Ÿ 3 6 ,Ÿ 3 , ,�  3 ,      H   , ,�� 2�t ,�� 3 , ,Ÿ 3 , ,Ÿ 2�t ,�� 2�t      H   , ,�  2�j ,�  2�t ,Ÿ 2�t ,Ÿ 2�j ,�  2�j      H   , -� 2s� -� 2s� -� 2s� -� 2s� -� 2s�      H   , ,�� 2g� ,�� 2s� -1� 2s� -1� 2g� ,�� 2g�      H   , -� 2g� -� 2g� -� 2g� -� 2g� -� 2g�      H   , ,�� 2-< ,�� 2-F ,�� 2-F ,�� 2-< ,�� 2-<      H   , ,�� 2!� ,�� 2-< -� 2-< -� 2!� ,�� 2!�      H   , ,�� 2!z ,�� 2!� ,�� 2!� ,�� 2!z ,�� 2!z      H   , ,�� 1�� ,�� 1�� ,װ 1�� ,װ 1�� ,�� 1��      H   , ,�� 1�4 ,�� 1�� ,� 1�� ,� 1�4 ,�� 1�4      H   , ,�� 1�* ,�� 1�4 ,װ 1�4 ,װ 1�* ,�� 1�*      H   , ,� 1�� ,� 1�� ,�� 1�� ,�� 1�� ,� 1��      H   , ,�� 1�� ,�� 1�� ,Ÿ 1�� ,Ÿ 1�� ,�� 1��      H   , ,� 1�� ,� 1�� ,�� 1�� ,�� 1�� ,� 1��      H   , -%� 1� -%� 1 -1� 1 -1� 1� -%� 1�      H   , ,�� 1D ,�� 1� -1� 1� -1� 1D ,�� 1D      H   , -%� 1: -%� 1D -1� 1D -1� 1: -%� 1:      H   , -� 0ͬ -� 0Ͷ -� 0Ͷ -� 0ͬ -� 0ͬ      H   , ,�� 0�� ,�� 0ͬ -� 0ͬ -� 0�� ,�� 0��      H   , -� 0�� -� 0�� -� 0�� -� 0�� -� 0��      H   , ,�� 0�\ ,�� 0�f ,� 0�f ,� 0�\ ,�� 0�\      H   , ,�� 0{� ,�� 0�\ ,� 0�\ ,� 0{� ,�� 0{�      H   , ,�� 0{� ,�� 0{� ,� 0{� ,� 0{� ,�� 0{�      H   , ,�  0A ,�  0A ,Ÿ 0A ,Ÿ 0A ,�  0A      H   , ,�� 05T ,�� 0A ,Ÿ 0A ,Ÿ 05T ,�� 05T      H   , ,�  05J ,�  05T ,Ÿ 05T ,Ÿ 05J ,�  05J      H   , -� /�l -� /�v -� /�v -� /�l -� /�l      H   , ,�� /�� ,�� /�l -1� /�l -1� /�� ,�� /��      H   , -� /�� -� /�� -� /�� -� /�� -� /��      H   , ,�� /n ,�� /n& ,�� /n& ,�� /n ,�� /n      H   , +u 68� +u 68� +�� 68� +�� 68� +u 68�      H   , (�� 68� (�� 68� (�� 68� (�� 68� (�� 68�      H   , -%� 6D� -%� 6D� -1� 6D� -1� 6D� -%� 6D�      H   , #7� 6D� #7� 6D� #Cl 6D� #Cl 6D� #7� 6D�      H   , "� 5�� "� 5�� "�� 5�� "�� 5�� "� 5��      H   , %j4 5�� %j4 5�� %u� 5�� %u� 5�� %j4 5��      H   , 'Vd 6&� 'Vd 6&� 'b 6&� 'b 6&� 'Vd 6&�      H   , #�T 5�
 #�T 5� #� 5� #� 5�
 #�T 5�
      H   , &�t 5�
 &�t 5� &�, 5� &�, 5�
 &�t 5�
      H   , 'Vd 62� 'Vd 62� 'b 62� 'b 62� 'Vd 62�      H   , !�$ 62� !�$ 62� !�� 62� !�� 62� !�$ 62�      H   , $
� 5� $
� 5�� $\ 5�� $\ 5� $
� 5�      H   , &�� 5� &�� 5�� &�| 5�� &�| 5� &�� 5�      H   , $P� 6� $P� 6� $\� 6� $\� 6� $P� 6�      H   , ' 6� ' 6� '� 6� '� 6� ' 6�      H   , "�d 6 � "�d 6 � "� 6 � "� 6 � "�d 6 �      H   , %�� 6D� %�� 6D� &� 6D� &� 6D� %�� 6D�      H   , $
� 5�� $
� 5� $\ 5� $\ 5�� $
� 5��      H   , &�� 5�� &�� 5� &�| 5� &�| 5�� &�� 5��      H   , %�� 6 � %�� 6 � %�< 6 � %�< 6 � %�� 6 �      H   , $P� 6� $P� 6� $\� 6� $\� 6� $P� 6�      H   , ' 6� ' 6� '� 6� '� 6� ' 6�      H   , "d� 5�� "d� 5�� "p| 5�� "p| 5�� "d� 5��      H   , %#� 5�� %#� 5�� %/� 5�� %/� 5�� %#� 5��      H   , $�D 62� $�D 62� $�� 62� $�� 62� $�D 62�      H   , !�$ 6&� !�$ 6&� !�� 6&� !�� 6&� !�$ 6&�      H   , "� 5�� "� 5�� "�� 5�� "�� 5�� "� 5��      H   , %j4 5�� %j4 5�� %u� 5�� %u� 5�� %j4 5��      H   , "d� 5� "d� 5� "p| 5� "p| 5� "d� 5�      H   , %#� 5� %#� 5� %/� 5� %/� 5� %#� 5�      H   , $�D 6&� $�D 6&� $�� 6&� $�� 6&� $�D 6&�      H   , "�d 6� "�d 6� "� 6� "� 6� "�d 6�      H   , %�� 6� %�� 6� %�< 6� %�< 6� %�� 6�      H   , #�T 5�� #�T 5�� #� 5�� #� 5�� #�T 5��      H   , &�t 5�� &�t 5�� &�, 5�� &�, 5�� &�t 5��      H   , #7� 68� #7� 68� #Cl 68� #Cl 68� #7� 68�      H   , %�� 68� %�� 68� &� 68� &� 68� %�� 68�      H   , ,� .�| ,� .� ,�� .� ,�� .�| ,� .�|      H   , ,�� .�� ,�� .�| ,Ÿ .�| ,Ÿ .�� ,�� .��      H   , ,� .պ ,� .�� ,�� .�� ,�� .պ ,� .պ      H   , -%� .T� -%� .T� -1� .T� -1� .T� -%� .T�      H   , ,�� .I$ ,�� .T� -1� .T� -1� .I$ ,�� .I$      H   , -%� .I -%� .I$ -1� .I$ -1� .I -%� .I      H   , -� .� -� .� -� .� -� .� -� .�      H   , ,�� .� ,�� .� -� .� -� .� ,�� .�      H   , -� .� -� .� -� .� -� .� -� .�      H   , ,�� -�< ,�� -�F ,� -�F ,� -�< ,�� -�<      H   , ,�� -�� ,�� -�< ,� -�< ,� -�� ,�� -��      H   , ,�� -�z ,�� -�� ,� -�� ,� -�z ,�� -�z      H   , ,�  -�� ,�  -�� ,Ÿ -�� ,Ÿ -�� ,�  -��      H   , ,�� -v4 ,�� -�� ,Ÿ -�� ,Ÿ -v4 ,�� -v4      H   , ,�  -v* ,�  -v4 ,Ÿ -v4 ,Ÿ -v* ,�  -v*      H   , -� ,�L -� ,�V -� ,�V -� ,�L -� ,�L      H   , ,�� ,� ,�� ,�L -1� ,�L -1� ,� ,�� ,�      H   , -� ,� -� ,� -� ,� -� ,� -� ,�      H   , ,�� ,�� ,�� ,� ,�� ,� ,�� ,�� ,�� ,��      H   , ,�� ,�D ,�� ,�� -� ,�� -� ,�D ,�� ,�D      H   , ,�� ,�: ,�� ,�D ,�� ,�D ,�� ,�: ,�� ,�:      H   , ,�� ,h� ,�� ,h� ,װ ,h� ,װ ,h� ,�� ,h�      H   , ,�� ,\� ,�� ,h� ,� ,h� ,� ,\� ,�� ,\�      H   , ,�� ,\� ,�� ,\� ,װ ,\� ,װ ,\� ,�� ,\�      H   , ,� ,"\ ,� ,"f ,�� ,"f ,�� ,"\ ,� ,"\      H   , ,�� ,� ,�� ,"\ ,Ÿ ,"\ ,Ÿ ,� ,�� ,�      H   , ,� ,� ,� ,� ,�� ,� ,�� ,� ,� ,�      H   , -%� +�� -%� +�� -1� +�� -1� +�� -%� +��      H   , ,�� +� ,�� +�� -1� +�� -1� +� ,�� +�      H   , -%� +�� -%� +� -1� +� -1� +�� -%� +��      H   , -� +Ol -� +Ov -� +Ov -� +Ol -� +Ol      H   , ,�� +C� ,�� +Ol -� +Ol -� +C� ,�� +C�      H   , -� +C� -� +C� -� +C� -� +C� -� +C�      H   , ,�� +	 ,�� +	& ,� +	& ,� +	 ,�� +	      H   , ,�� *�d ,�� +	 ,� +	 ,� *�d ,�� *�d      H   , ,�� *�Z ,�� *�d ,� *�d ,� *�Z ,�� *�Z      H   , ,�  *�� ,�  *�� ,Ÿ *�� ,Ÿ *�� ,�  *��      H   , ,�� *� ,�� *�� ,Ÿ *�� ,Ÿ *� ,�� *�      H   , ,�  *�
 ,�  *� ,Ÿ *� ,Ÿ *�
 ,�  *�
      H   , -� *6, -� *66 -� *66 -� *6, -� *6,      H   , ,�� **t ,�� *6, -1� *6, -1� **t ,�� **t      H   , -� **j -� **t -� **t -� **j -� **j      H   , ,�� )�� ,�� )�� ,�� )�� ,�� )�� ,�� )��      H   , ,�� )�$ ,�� )�� -� )�� -� )�$ ,�� )�$      H   , ,�� )� ,�� )�$ ,�� )�$ ,�� )� ,�� )�      H   , ,�� )�� ,�� )�� ,װ )�� ,װ )�� ,�� )��      H   , ,�� )�� ,�� )�� ,� )�� ,� )�� ,�� )��      H   , ,�� )�� ,�� )�� ,װ )�� ,װ )�� ,�� )��      H   , ,� )c< ,� )cF ,�� )cF ,�� )c< ,� )c<      H   , ,�� )W� ,�� )c< ,Ÿ )c< ,Ÿ )W� ,�� )W�      H   , ,� )Wz ,� )W� ,�� )W� ,�� )Wz ,� )Wz      H   , -%� (֜ -%� (֦ -1� (֦ -1� (֜ -%� (֜      H   , ,�� (�� ,�� (֜ -1� (֜ -1� (�� ,�� (��      H   , -%� (�� -%� (�� -1� (�� -1� (�� -%� (��      H   , -� (�L -� (�V -� (�V -� (�L -� (�L      H   , ,�� /bZ ,�� /bd ,�� /bd ,�� /bZ ,�� /bZ      H   , ,�� /'� ,�� /'� ,װ /'� ,װ /'� ,�� /'�      H   , ,�� / ,�� /'� ,� /'� ,� / ,�� /      H   , ,�� /
 ,�� / ,װ / ,װ /
 ,�� /
      H   , Y� 62� Y� 62� e� 62� e� 62� Y� 62�      H   , �� 5�
 �� 5� ӌ 5� ӌ 5�
 �� 5�
      H   , �� 5�
 �� 5� �� 5� �� 5�
 �� 5�
      H   , F 5�
 F 5� Q� 5� Q� 5�
 F 5�
      H   , !4 5�
 !4 5� !� 5� !� 5�
 !4 5�
      H   , �� 5�� �� 5�� �L 5�� �L 5�� �� 5��      H   , m� 5�� m� 5�� yl 5�� yl 5�� m� 5��      H   , ,� 5�� ,� 5�� 8� 5�� 8� 5�� ,� 5��      H   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      H   ,  62�  62� $� 62� $� 62�  62�      H   , ۤ 62� ۤ 62� �\ 62� �\ 62� ۤ 62�      H   , �T 6D� �T 6D�  6D�  6D� �T 6D�      H   , �� 6 � �� 6 �  � 6 �  � 6 � �� 6 �      H   , �T 6� �T 6� � 6� � 6� �T 6�      H   , O 5� O 5�� Z� 5�� Z� 5� O 5�      H   , $ 5� $ 5�� � 5�� � 5� $ 5�      H   , �D 5� �D 5�� �� 5�� �� 5� �D 5�      H   , �d 5� �d 5�� � 5�� � 5� �d 5�      H   , !K� 5� !K� 5�� !W< 5�� !W< 5� !K� 5�      H   , Tt 6� Tt 6� `, 6� `, 6� Tt 6�      H   , � 6� � 6� L 6� L 6� � 6�      H   , Ҵ 6� Ҵ 6� �l 6� �l 6� Ҵ 6�      H   , !�� 6� !�� 6� !�� 6� !�� 6� !�� 6�      H   , � 6 � � 6 � �� 6 � �� 6 � � 6 �      H   , s$ 6 � s$ 6 � ~� 6 � ~� 6 � s$ 6 �      H   , O 5�� O 5� Z� 5� Z� 5�� O 5��      H   , $ 5�� $ 5� � 5� � 5�� $ 5��      H   , �D 5�� �D 5� �� 5� �� 5�� �D 5��      H   , �d 5�� �d 5� � 5� � 5�� �d 5��      H   , !K� 5�� !K� 5� !W< 5� !W< 5�� !K� 5��      H   ,  2D 6 �  2D 6 �  =� 6 �  =� 6 �  2D 6 �      H   , ۤ 6&� ۤ 6&� �\ 6&� �\ 6&� ۤ 6&�      H   ,  x� 6D�  x� 6D�  �L 6D�  �L 6D�  x� 6D�      H   , �T 6� �T 6� � 6� � 6� �T 6�      H   , Tt 6� Tt 6� `, 6� `, 6� Tt 6�      H   , hD 5�� hD 5�� s� 5�� s� 5�� hD 5��      H   , 'd 5�� 'd 5�� 3 5�� 3 5�� 'd 5��      H   , � 5�� � 5�� �< 5�� �< 5�� � 5��      H   , �� 5�� �� 5�� �\ 5�� �\ 5�� �� 5��      H   , � 6� � 6� L 6� L 6� � 6�      H   , Ҵ 6� Ҵ 6� �l 6� �l 6� Ҵ 6�      H   , !�� 6� !�� 6� !�� 6� !�� 6� !�� 6�      H   , �� 6&� �� 6&� �| 6&� �| 6&� �� 6&�      H   , Y� 6&� Y� 6&� e� 6&� e� 6&� Y� 6&�      H   ,  6&�  6&� $� 6&� $� 6&�  6&�      H   , hD 5� hD 5� s� 5� s� 5� hD 5�      H   , 'd 5� 'd 5� 3 5� 3 5� 'd 5�      H   , � 5� � 5� �< 5� �< 5� � 5�      H   , �� 5� �� 5� �\ 5� �\ 5� �� 5�      H   , �� 62� �� 62� �| 62� �| 62� �� 62�      H   , �� 5�� �� 5�� �L 5�� �L 5�� �� 5��      H   , m� 5�� m� 5�� yl 5�� yl 5�� m� 5��      H   , ,� 5�� ,� 5�� 8� 5�� 8� 5�� ,� 5��      H   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      H   , �� 5�� �� 5�� ӌ 5�� ӌ 5�� �� 5��      H   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      H   , F 5�� F 5�� Q� 5�� Q� 5�� F 5��      H   , !4 5�� !4 5�� !� 5�� !� 5�� !4 5��      H   , �t 6D� �t 6D� �, 6D� �, 6D� �t 6D�      H   , �� 6� �� 6�  � 6�  � 6� �� 6�      H   , � 6� � 6� �� 6� �� 6� � 6�      H   , ;4 6D� ;4 6D� F� 6D� F� 6D� ;4 6D�      H   , ;4 68� ;4 68� F� 68� F� 68� ;4 68�      H   , �T 68� �T 68�  68�  68� �T 68�      H   , �t 68� �t 68� �, 68� �, 68� �t 68�      H   ,  x� 68�  x� 68�  �L 68�  �L 68�  x� 68�      H   , s$ 6� s$ 6� ~� 6� ~� 6� s$ 6�      H   ,  2D 6�  2D 6�  =� 6�  =� 6�  2D 6�      H   , ,�� 'kT ,�� 'w -1� 'w -1� 'kT ,�� 'kT      H   , -� 'kJ -� 'kT -� 'kT -� 'kJ -� 'kJ      H   , ,�� '0� ,�� '0� ,�� '0� ,�� '0� ,�� '0�      H   , ,�� '% ,�� '0� -� '0� -� '% ,�� '%      H   , ,�� '$� ,�� '% ,�� '% ,�� '$� ,�� '$�      H   , ,�� &�l ,�� &�v ,װ &�v ,װ &�l ,�� &�l      H   , ,�� &޴ ,�� &�l ,� &�l ,� &޴ ,�� &޴      H   , ,�� &ު ,�� &޴ ,װ &޴ ,װ &ު ,�� &ު      H   , ,� &� ,� &�& ,�� &�& ,�� &� ,� &�      H   , ,�� &�d ,�� &� ,Ÿ &� ,Ÿ &�d ,�� &�d      H   , ,� &�Z ,� &�d ,�� &�d ,�� &�Z ,� &�Z      H   , -%� &| -%� &� -1� &� -1� &| -%� &|      H   , ,�� &� ,�� &| -1� &| -1� &� ,�� &�      H   , -%� &� -%� &� -1� &� -1� &� -%� &�      H   , -� %�, -� %�6 -� %�6 -� %�, -� %�,      H   , ,�� %�t ,�� %�, -� %�, -� %�t ,�� %�t      H   , -� %�j -� %�t -� %�t -� %�j -� %�j      H   , ,�� %�� ,�� %�� ,� %�� ,� %�� ,�� %��      H   , ,�� %$ ,�� %�� ,� %�� ,� %$ ,�� %$      H   , ,�� % ,�� %$ ,� %$ ,� % ,�� %      H   , ,�  %D� ,�  %D� ,Ÿ %D� ,Ÿ %D� ,�  %D�      H   , ,�� %8� ,�� %D� ,Ÿ %D� ,Ÿ %8� ,�� %8�      H   , ,�  %8� ,�  %8� ,Ÿ %8� ,Ÿ %8� ,�  %8�      H   , -� $�� -� $�� -� $�� -� $�� -� $��      H   , ,�� $�4 ,�� $�� -1� $�� -1� $�4 ,�� $�4      H   , -� $�* -� $�4 -� $�4 -� $�* -� $�*      H   , ,�� $q� ,�� $q� ,�� $q� ,�� $q� ,�� $q�      H   , ,�� $e� ,�� $q� -� $q� -� $e� ,�� $e�      H   , ,�� $e� ,�� $e� ,�� $e� ,�� $e� ,�� $e�      H   , ,�� $+L ,�� $+V ,װ $+V ,װ $+L ,�� $+L      H   , ,�� $� ,�� $+L ,� $+L ,� $� ,�� $�      H   , ,�� $� ,�� $� ,װ $� ,װ $� ,�� $�      H   , ,� #�� ,� #� ,�� #� ,�� #�� ,� #��      H   , ,�� #�D ,�� #�� ,Ÿ #�� ,Ÿ #�D ,�� #�D      H   , ,� #�: ,� #�D ,�� #�D ,�� #�: ,� #�:      H   , -%� #X\ -%� #Xf -1� #Xf -1� #X\ -%� #X\      H   , ,�� #L� ,�� #X\ -1� #X\ -1� #L� ,�� #L�      H   , -%� #L� -%� #L� -1� #L� -1� #L� -%� #L�      H   , -� # -� # -� # -� # -� #      H   , ,�� #T ,�� # -� # -� #T ,�� #T      H   , -� #J -� #T -� #T -� #J -� #J      H   , ,�� "˼ ,�� "�� ,� "�� ,� "˼ ,�� "˼      H   , ,�� "� ,�� "˼ ,� "˼ ,� "� ,�� "�      H   , ,�� "�� ,�� "� ,� "� ,� "�� ,�� "��      H   , ,�  "�l ,�  "�v ,Ÿ "�v ,Ÿ "�l ,�  "�l      H   , ,�� "y� ,�� "�l ,Ÿ "�l ,Ÿ "y� ,�� "y�      H   , ,�  "y� ,�  "y� ,Ÿ "y� ,Ÿ "y� ,�  "y�      H   , -� !�� -� !�� -� !�� -� !�� -� !��      H   , ,�� !� ,�� !�� -1� !�� -1� !� ,�� !�      H   , -� !�
 -� !� -� !� -� !�
 -� !�
      H   , -� (�� -� (�� -� (�� -� (�� -� (��      H   , ,�� (I� ,�� (J ,� (J ,� (I� ,�� (I�      H   , ,�� (>D ,�� (I� ,� (I� ,� (>D ,�� (>D      H   , ,�� (>: ,�� (>D ,� (>D ,� (>: ,�� (>:      H   , ,�  (� ,�  (� ,Ÿ (� ,Ÿ (� ,�  (�      H   , ,�� '�� ,�� (� ,Ÿ (� ,Ÿ '�� ,�� '��      H   , ,�  '�� ,�  '�� ,Ÿ '�� ,Ÿ '�� ,�  '��      H   , -� 'w -� 'w -� 'w -� 'w -� 'w      H   , ,� ! ,� !$ ,�� !$ ,�� ! ,� !      H   , -%�  �< -%�  �F -1�  �F -1�  �< -%�  �<      H   , ,��  �� ,��  �< -1�  �< -1�  �� ,��  ��      H   , -%�  �z -%�  �� -1�  �� -1�  �z -%�  �z      H   , -�  R� -�  R� -�  R� -�  R� -�  R�      H   , ,��  G4 ,��  R� -�  R� -�  G4 ,��  G4      H   , -�  G* -�  G4 -�  G4 -�  G* -�  G*      H   , ,��  � ,��  � ,�  � ,�  � ,��  �      H   , ,��   � ,��  � ,�  � ,�   � ,��   �      H   , ,��   � ,��   � ,�   � ,�   � ,��   �      H   , ,�  �L ,�  �V ,Ÿ �V ,Ÿ �L ,�  �L      H   , ,�� �� ,�� �L ,Ÿ �L ,Ÿ �� ,�� ��      H   , ,�  �� ,�  �� ,Ÿ �� ,Ÿ �� ,�  ��      H   , -� 9� -� 9� -� 9� -� 9� -� 9�      H   , ,�� -� ,�� 9� -1� 9� -1� -� ,�� -�      H   , -� -� -� -� -� -� -� -� -� -�      H   , ,�� �\ ,�� �f ,�� �f ,�� �\ ,�� �\      H   , ,�� � ,�� �\ -� �\ -� � ,�� �      H   , ,�� � ,�� � ,�� � ,�� � ,�� �      H   , ,�� � ,�� � ,װ � ,װ � ,�� �      H   , ,�� �T ,�� � ,� � ,� �T ,�� �T      H   , ,�� �J ,�� �T ,װ �T ,װ �J ,�� �J      H   , ,� f� ,� f� ,�� f� ,�� f� ,� f�      H   , ,�� [ ,�� f� ,Ÿ f� ,Ÿ [ ,�� [      H   , ,� Z� ,� [ ,�� [ ,�� Z� ,� Z�      H   , -%� � -%� �& -1� �& -1� � -%� �      H   , ,�� �d ,�� � -1� � -1� �d ,�� �d      H   , -%� �Z -%� �d -1� �d -1� �Z -%� �Z      H   , -� �� -� �� -� �� -� �� -� ��      H   , ,�� � ,�� �� -� �� -� � ,�� �      H   , -� �
 -� � -� � -� �
 -� �
      H   , ,�� M| ,�� M� ,� M� ,� M| ,�� M|      H   , ,�� A� ,�� M| ,� M| ,� A� ,�� A�      H   , ,�� A� ,�� A� ,� A� ,� A� ,�� A�      H   , ,�  , ,�  6 ,Ÿ 6 ,Ÿ , ,�  ,      H   , ,�� �t ,�� , ,Ÿ , ,Ÿ �t ,�� �t      H   , ,�  �j ,�  �t ,Ÿ �t ,Ÿ �j ,�  �j      H   , -� z� -� z� -� z� -� z� -� z�      H   , ,�� n� ,�� z� -1� z� -1� n� ,�� n�      H   , -� n� -� n� -� n� -� n� -� n�      H   , ,�� 4< ,�� 4F ,�� 4F ,�� 4< ,�� 4<      H   , ,�� (� ,�� 4< -� 4< -� (� ,�� (�      H   , ,�� (z ,�� (� ,�� (� ,�� (z ,�� (z      H   , ,�� �� ,�� �� ,װ �� ,װ �� ,�� ��      H   , ,�� �4 ,�� �� ,� �� ,� �4 ,�� �4      H   , ,�� �* ,�� �4 ,װ �4 ,װ �* ,�� �*      H   , ,� �� ,� �� ,�� �� ,�� �� ,� ��      H   , ,�� �� ,�� �� ,Ÿ �� ,Ÿ �� ,�� ��      H   , ,� �� ,� �� ,�� �� ,�� �� ,� ��      H   , -%� � -%�  -1�  -1� � -%� �      H   , ,�� D ,�� � -1� � -1� D ,�� D      H   , -%� : -%� D -1� D -1� : -%� :      H   , ,�� !�| ,�� !�� ,�� !�� ,�� !�| ,�� !�|      H   , ,�� !�� ,�� !�| -� !�| -� !�� ,�� !��      H   , ,�� !�� ,�� !�� ,�� !�� ,�� !�� ,�� !��      H   , ,�� !l, ,�� !l6 ,װ !l6 ,װ !l, ,�� !l,      H   , ,�� !`t ,�� !l, ,� !l, ,� !`t ,�� !`t      H   , ,�� !`j ,�� !`t ,װ !`t ,װ !`j ,�� !`j      H   , ,� !%� ,� !%� ,�� !%� ,�� !%� ,� !%�      H   , ,�� !$ ,�� !%� ,Ÿ !%� ,Ÿ !$ ,�� !$      H   ,��, (����, (�L  	` (�L  	` (����, (��      H   , >� 68� >� 68� Jl 68� Jl 68� >� 68�      H   , R� 5�� R� 5� ^< 5� ^< 5�� R� 5��      H   , � 5�� � 5� \ 5� \ 5�� � 5��      H   , �� 5�� �� 5� �| 5� �| 5�� �� 5��      H   , �� 5�� �� 5� �� 5� �� 5�� �� 5��      H   , �� 68� �� 68� 	� 68� 	� 68� �� 68�      H   , �� 68� �� 68� Ȭ 68� Ȭ 68� �� 68�      H   , | 68� | 68� �� 68� �� 68� | 68�      H   , k� 5�� k� 5�� w| 5�� w| 5�� k� 5��      H   , *� 5�� *� 5�� 6� 5�� 6� 5�� *� 5��      H   , � 5�� � 5�� �� 5�� �� 5�� � 5��      H   , �$ 5�� �$ 5�� �� 5�� �� 5�� �$ 5��      H   , �� 6� �� 6� �� 6� �� 6� �� 6�      H   , W� 6� W� 6� c� 6� c� 6� W� 6�      H   ,  6�  6� "� 6� "� 6�  6�      H   , �4 6� �4 6� �� 6� �� 6� �4 6�      H   , �$ 6&� �$ 6&� �� 6&� �� 6&� �$ 6&�      H   , �D 6&� �D 6&� �� 6&� �� 6&� �D 6&�      H   , k� 5� k� 5� w| 5� w| 5� k� 5�      H   , *� 5� *� 5� 6� 5� 6� 5� *� 5�      H   , � 5� � 5� �� 5� �� 5� � 5�      H   , �$ 5� �$ 5� �� 5� �� 5� �$ 5�      H   , ]d 6&� ]d 6&� i 6&� i 6&� ]d 6&�      H   , � 6&� � 6&� (< 6&� (< 6&� � 6&�      H   , 5� 6� 5� 6� A| 6� A| 6� 5� 6�      H   , 4 5�� 4 5�� � 5�� � 5�� 4 5��      H   , �T 5�� �T 5�� � 5�� � 5�� �T 5��      H   , �t 5�� �t 5�� �, 5�� �, 5�� �t 5��      H   , I� 5�� I� 5�� UL 5�� UL 5�� I� 5��      H   , � 5�� � 5�� l 5�� l 5�� � 5��      H   , �� 6� �� 6� �� 6� �� 6� �� 6�      H   , W� 6� W� 6� c� 6� c� 6� W� 6�      H   ,  6�  6� "� 6� "� 6�  6�      H   , �4 6� �4 6� �� 6� �� 6� �4 6�      H   , >� 6D� >� 6D� Jl 6D� Jl 6D� >� 6D�      H   , �� 6D� �� 6D� 	� 6D� 	� 6D� �� 6D�      H   , �� 6D� �� 6D� Ȭ 6D� Ȭ 6D� �� 6D�      H   , | 6D� | 6D� �� 6D� �� 6D� | 6D�      H   , 4 5�
 4 5� � 5� � 5�
 4 5�
      H   , �T 5�
 �T 5� � 5� � 5�
 �T 5�
      H   , �t 5�
 �t 5� �, 5� �, 5�
 �t 5�
      H   , I� 5�
 I� 5� UL 5� UL 5�
 I� 5�
      H   , � 5�
 � 5� l 5� l 5�
 � 5�
      H   , � 5�� � 5�� �� 5�� �� 5�� � 5��      H   , q4 5�� q4 5�� |� 5�� |� 5�� q4 5��      H   , 0T 5�� 0T 5�� < 5�� < 5�� 0T 5��      H   , �t 5�� �t 5�� �, 5�� �, 5�� �t 5��      H   , �d 6 � �d 6 �  6 �  6 � �d 6 �      H   , �� 6 � �� 6 � �< 6 � �< 6 � �� 6 �      H   , v� 6 � v� 6 � �\ 6 � �\ 6 � v� 6 �      H   , 5� 6 � 5� 6 � A| 6 � A| 6 � 5� 6 �      H   , � 5�� � 5�� �� 5�� �� 5�� � 5��      H   , q4 5�� q4 5�� |� 5�� |� 5�� q4 5��      H   , 0T 5�� 0T 5�� < 5�� < 5�� 0T 5��      H   , �t 5�� �t 5�� �, 5�� �, 5�� �t 5��      H   , �$ 62� �$ 62� �� 62� �� 62� �$ 62�      H   , �D 62� �D 62� �� 62� �� 62� �D 62�      H   , ]d 62� ]d 62� i 62� i 62� ]d 62�      H   , � 62� � 62� (< 62� (< 62� � 62�      H   , R� 5� R� 5�� ^< 5�� ^< 5� R� 5�      H   , � 5� � 5�� \ 5�� \ 5� � 5�      H   , �� 5� �� 5�� �| 5�� �| 5� �� 5�      H   , �� 5� �� 5�� �� 5�� �� 5� �� 5�      H   , �d 6� �d 6�  6�  6� �d 6�      H   , �� 6� �� 6� �< 6� �< 6� �� 6�      H   , v� 6� v� 6� �\ 6� �\ 6� v� 6�      H   ,��, /bd��, /n  	` /n  	` /bd��, /bd      H   , `� 6&� `� 6&� l� 6&� l� 6&� `� 6&�      H   , 	  6&� 	  6&� 	+� 6&� 	+� 6&� 	  6&�      H   , �d 5�� �d 5� � 5� � 5�� �d 5��      H   , � 5� � 5� �< 5� �< 5� � 5�      H   , 	�� 5� 	�� 5� 	�\ 5� 	�\ 5� 	�� 5�      H   , �t 68� �t 68� �, 68� �, 68� �t 68�      H   , �t 6D� �t 6D� �, 6D� �, 6D� �t 6D�      H   , � 6� � 6� &L 6� &L 6� � 6�      H   , ٴ 6� ٴ 6� �l 6� �l 6� ٴ 6�      H   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      H   , M 5�� M 5�� X� 5�� X� 5�� M 5��      H   , 
� 68� 
� 68� 
�L 68� 
�L 68� 
� 68�      H   , 
� 6D� 
� 6D� 
�L 6D� 
�L 6D� 
� 6D�      H   , �� 5�
 �� 5� �� 5� �� 5�
 �� 5�
      H   , M 5�
 M 5� X� 5� X� 5�
 M 5�
      H   , 3� 5�� 3� 5�� ?� 5�� ?� 5�� 3� 5��      H   , 	�� 5�� 	�� 5�� 	�� 5�� 	�� 5�� 	�� 5��      H   , � 6� � 6� &L 6� &L 6� � 6�      H   , ٴ 6� ٴ 6� �l 6� �l 6� ٴ 6�      H   , z$ 6 � z$ 6 � �� 6 � �� 6 � z$ 6 �      H   , 
9D 6 � 
9D 6 � 
D� 6 � 
D� 6 � 
9D 6 �      H   , `� 62� `� 62� l� 62� l� 62� `� 62�      H   , 3� 5�� 3� 5�� ?� 5�� ?� 5�� 3� 5��      H   , 	�� 5�� 	�� 5�� 	�� 5�� 	�� 5�� 	�� 5��      H   , � 5�� � 5�� �< 5�� �< 5�� � 5��      H   , 	  62� 	  62� 	+� 62� 	+� 62� 	  62�      H   , 	�� 5�� 	�� 5�� 	�\ 5�� 	�\ 5�� 	�� 5��      H   , �D 5� �D 5�� �� 5�� �� 5� �D 5�      H   , �d 5� �d 5�� � 5�� � 5� �d 5�      H   , �D 5�� �D 5� �� 5� �� 5�� �D 5��      H   , z$ 6� z$ 6� �� 6� �� 6� z$ 6�      H   , 
9D 6� 
9D 6� 
D� 6� 
D� 6� 
9D 6�      H   ,��m4 6&���m4 6&���x� 6&���x� 6&���m4 6&�      H   ,���$ 6����$ 6����� 6����� 6����$ 6�      H   ,��[< 6D���[< 6D���f� 6D���f� 6D���[< 6D�      H   ,��� 5�
��� 5���� 5���� 5�
��� 5�
      H   ,  � 5�
  � 5�  l 5�  l 5�
  � 5�
      H   , �� 5�
 �� 5� ڌ 5� ڌ 5�
 �� 5�
      H   , �� 6&� �� 6&� �| 6&� �| 6&� �� 6&�      H   , T 6D� T 6D�  6D�  6D� T 6D�      H   ,  �T 6�  �T 6�  � 6�  � 6�  �T 6�      H   , [t 6� [t 6� g, 6� g, 6� [t 6�      H   ,��m4 62���m4 62���x� 62���x� 62���m4 62�      H   ,��, 6 ���, 6 ����� 6 ����� 6 ���, 6 �      H   , �� 6 � �� 6 � � 6 � � 6 � �� 6 �      H   ,��� 5����� 5������ 5������ 5����� 5��      H   , �� 5�� �� 5�� �L 5�� �L 5�� �� 5��      H   , t� 5�� t� 5�� �l 5�� �l 5�� t� 5��      H   ,��� 5���� 5����� 5����� 5���� 5�      H   ,���$ 6����$ 6����� 6����� 6����$ 6�      H   ,  �T 6�  �T 6�  � 6�  � 6�  �T 6�      H   ,��m4 52���m4 52���x� 52���x� 52���m4 52�      H   ,��[< 5&���[< 52�  	` 52�  	` 5&���[< 5&�      H   , [t 6� [t 6� g, 6� g, 6� [t 6�      H   ,��m4 5&���m4 5&���x� 5&���x� 5&���m4 5&�      H   ,���$ 4�\���$ 4�f���� 4�f���� 4�\���$ 4�\      H   , � 6 � � 6 � Ƽ 6 � Ƽ 6 � � 6 �      H   ,��, 4���, 4�\  	` 4�\  	` 4���, 4�      H   , oD 5� oD 5� z� 5� z� 5� oD 5�      H   ,���$ 4�����$ 4����� 4����� 4�����$ 4��      H   , .d 5� .d 5� : 5� : 5� .d 5�      H   ,��� 4���� 4����� 4����� 4���� 4�      H   ,��� 5����� 5������ 5������ 5����� 5��      H   ,��� 4�T��� 4�  	` 4�  	` 4�T��� 4�T      H   ,��� 4�J��� 4�T���� 4�T���� 4�J��� 4�J      H   , oD 5�� oD 5�� z� 5�� z� 5�� oD 5��      H   ,��� 4_���� 4_���� 4_���� 4_���� 4_�      H   ,��� 4T��� 4_�  	` 4_�  	` 4T��� 4T      H   ,  � 62�  � 62�  �\ 62�  �\ 62�  � 62�      H   ,��� 4S���� 4T��� 4T��� 4S���� 4S�      H   , �� 62� �� 62� �| 62� �| 62� �� 62�      H   ,��[< 3���[< 3�&��f� 3�&��f� 3���[< 3�      H   ,��� 5����� 5����� 5����� 5����� 5��      H   ,��[< 3�d��[< 3�  	` 3�  	` 3�d��[< 3�d      H   ,��� 5����� 5������ 5������ 5����� 5��      H   ,��[< 3�Z��[< 3�d��f� 3�d��f� 3�Z��[< 3�Z      H   , �� 5�� �� 5�� �L 5�� �L 5�� �� 5��      H   ,��, 3����, 3������ 3������ 3����, 3��      H   , t� 5�� t� 5�� �l 5�� �l 5�� t� 5��      H   ,��, 3���, 3��  	` 3��  	` 3���, 3�      H   ,  � 5��  � 5��  l 5��  l 5��  � 5��      H   ,��, 3�
��, 3����� 3����� 3�
��, 3�
      H   , �� 5�� �� 5�� ڌ 5�� ڌ 5�� �� 5��      H   ,��� 3F|��� 3F����� 3F����� 3F|��� 3F|      H   , .d 5�� .d 5�� : 5�� : 5�� .d 5��      H   ,��� 3:���� 3F|  	` 3F|  	` 3:���� 3:�      H   ,��� 3:���� 3:����� 3:����� 3:���� 3:�      H   , $ 5�� $ 5�  � 5�  � 5�� $ 5��      H   ,��� 3 ,��� 3 6���� 3 6���� 3 ,��� 3 ,      H   ,��� 2�t��� 3 ,  	` 3 ,  	` 2�t��� 2�t      H   ,  � 6&�  � 6&�  �\ 6&�  �\ 6&�  � 6&�      H   ,��� 2�j��� 2�t���� 2�t���� 2�j��� 2�j      H   ,��[< /����[< /�l  	` /�l  	` /����[< /��      H   ,��m4 2s���m4 2s���x� 2s���x� 2s���m4 2s�      H   ,��[< 2g���[< 2s�  	` 2s�  	` 2g���[< 2g�      H   ,���$ /n���$ /n&���� /n&���� /n���$ /n      H   ,��m4 2g���m4 2g���x� 2g���x� 2g���m4 2g�      H   ,���$ 2-<���$ 2-F���� 2-F���� 2-<���$ 2-<      H   ,��[< 68���[< 68���f� 68���f� 68���[< 68�      H   ,��, 2!���, 2-<  	` 2-<  	` 2!���, 2!�      H   , B4 68� B4 68� M� 68� M� 68� B4 68�      H   ,���$ 2!z���$ 2!����� 2!����� 2!z���$ 2!z      H   ,��, 6���, 6����� 6����� 6���, 6�      H   ,��� 1����� 1������ 1������ 1����� 1��      H   , �� 6� �� 6� � 6� � 6� �� 6�      H   ,��� 1�4��� 1��  	` 1��  	` 1�4��� 1�4      H   ,��� 5���� 5������ 5������ 5���� 5�      H   ,��� 1�*��� 1�4���� 1�4���� 1�*��� 1�*      H   ,  V 5�  V 5��  a� 5��  a� 5�  V 5�      H   ,��� 1����� 1����� 1����� 1����� 1��      H   , $ 5� $ 5��  � 5��  � 5� $ 5�      H   ,��� 1����� 1��  	` 1��  	` 1����� 1��      H   , T 68� T 68�  68�  68� T 68�      H   ,��� 1����� 1����� 1����� 1����� 1��      H   ,��m4 /����m4 /����x� /����x� /����m4 /��      H   ,��[< 1���[< 1��f� 1��f� 1���[< 1�      H   ,��� 5����� 5����� 5����� 5����� 5��      H   ,��[< 1D��[< 1�  	` 1�  	` 1D��[< 1D      H   ,��[< 1:��[< 1D��f� 1D��f� 1:��[< 1:      H   ,��� 05J��� 05T���� 05T���� 05J��� 05J      H   ,��, 0ͬ��, 0Ͷ���� 0Ͷ���� 0ͬ��, 0ͬ      H   ,��, 0����, 0ͬ  	` 0ͬ  	` 0����, 0��      H   , � 6� � 6� Ƽ 6� Ƽ 6� � 6�      H   ,��, 0����, 0������ 0������ 0����, 0��      H   , B4 6D� B4 6D� M� 6D� M� 6D� B4 6D�      H   ,��� 0�\��� 0�f���� 0�f���� 0�\��� 0�\      H   ,��m4 /�l��m4 /�v��x� /�v��x� /�l��m4 /�l      H   ,��� 0{���� 0�\  	` 0�\  	` 0{���� 0{�      H   ,  V 5��  V 5�  a� 5�  a� 5��  V 5��      H   ,��� 0{���� 0{����� 0{����� 0{���� 0{�      H   ,��� 0A��� 0A���� 0A���� 0A��� 0A      H   ,��� 05T��� 0A  	` 0A  	` 05T��� 05T      H   ,���$ )�����$ )������ )������ )�����$ )��      H   ,��, +Ol��, +Ov���� +Ov���� +Ol��, +Ol      H   ,��, )�$��, )��  	` )��  	` )�$��, )�$      H   ,��� -�<��� -�F���� -�F���� -�<��� -�<      H   ,��� /��� /'�  	` /'�  	` /��� /      H   ,��[< ,���[< ,�L  	` ,�L  	` ,���[< ,�      H   ,��� -����� -�<  	` -�<  	` -����� -��      H   ,���$ )����$ )�$���� )�$���� )����$ )�      H   ,��� -�z��� -������ -������ -�z��� -�z      H   ,��m4 ,���m4 ,���x� ,���x� ,���m4 ,�      H   ,��, +C���, +Ol  	` +Ol  	` +C���, +C�      H   ,��� )����� )������ )������ )����� )��      H   ,��� ,���� ,���� ,���� ,���� ,�      H   ,��� )����� )��  	` )��  	` )����� )��      H   ,��, +C���, +C����� +C����� +C���, +C�      H   ,���$ ,�����$ ,����� ,����� ,�����$ ,��      H   ,��� )����� )������ )������ )����� )��      H   ,��� ,"\��� ,"f��� ,"f��� ,"\��� ,"\      H   ,��� )c<��� )cF��� )cF��� )c<��� )c<      H   ,��, ,�D��, ,��  	` ,��  	` ,�D��, ,�D      H   ,��� +	��� +	&���� +	&���� +	��� +	      H   ,��� )W���� )c<  	` )c<  	` )W���� )W�      H   ,��� -����� -������ -������ -����� -��      H   ,��[< +����[< +����f� +����f� +����[< +��      H   ,��� )Wz��� )W���� )W���� )Wz��� )Wz      H   ,��� *�d��� +	  	` +	  	` *�d��� *�d      H   ,��� -v4��� -��  	` -��  	` -v4��� -v4      H   ,��[< (֜��[< (֦��f� (֦��f� (֜��[< (֜      H   ,��� /'���� /'����� /'����� /'���� /'�      H   ,��[< (����[< (֜  	` (֜  	` (����[< (��      H   ,��� *�Z��� *�d���� *�d���� *�Z��� *�Z      H   ,��[< (����[< (����f� (����f� (����[< (��      H   ,��[< +���[< +��  	` +��  	` +���[< +�      H   ,��, (�L��, (�V���� (�V���� (�L��, (�L      H   ,��� *����� *������ *������ *����� *��      H   ,��� .պ��� .����� .����� .պ��� .պ      H   ,��� -v*��� -v4���� -v4���� -v*��� -v*      H   ,��� ,���� ,"\  	` ,"\  	` ,���� ,�      H   ,��[< .T���[< .T���f� .T���f� .T���[< .T�      H   ,��� *���� *��  	` *��  	` *���� *�      H   ,��m4 ,�L��m4 ,�V��x� ,�V��x� ,�L��m4 ,�L      H   ,���$ ,�:���$ ,�D���� ,�D���� ,�:���$ ,�:      H   ,��[< .I$��[< .T�  	` .T�  	` .I$��[< .I$      H   ,��� /
��� /���� /���� /
��� /
      H   ,��[< .I��[< .I$��f� .I$��f� .I��[< .I      H   ,��� ,h���� ,h����� ,h����� ,h���� ,h�      H   ,��� *�
��� *����� *����� *�
��� *�
      H   ,��, .���, .����� .����� .���, .�      H   ,��[< +����[< +���f� +���f� +����[< +��      H   ,��m4 *6,��m4 *66��x� *66��x� *6,��m4 *6,      H   ,��, .���, .�  	` .�  	` .���, .�      H   ,��� .�|��� .���� .���� .�|��� .�|      H   ,��, .���, .����� .����� .���, .�      H   ,��[< **t��[< *6,  	` *6,  	` **t��[< **t      H   ,��� ,\���� ,\����� ,\����� ,\���� ,\�      H   ,��� ,\���� ,h�  	` ,h�  	` ,\���� ,\�      H   ,��m4 **j��m4 **t��x� **t��x� **j��m4 **j      H   ,���$ /bZ���$ /bd���� /bd���� /bZ���$ /bZ      H   ,��� .����� .�|  	` .�|  	` .����� .��      H   ,��, (����, (������ (������ (����, (��      H   ,��[< $�4��[< $��  	` $��  	` $�4��[< $�4      H   ,��� &���� &�&��� &�&��� &���� &�      H   ,��m4 $�*��m4 $�4��x� $�4��x� $�*��m4 $�*      H   ,��[< 'kT��[< 'w  	` 'w  	` 'kT��[< 'kT      H   ,���$ $q����$ $q����� $q����� $q����$ $q�      H   ,��� &�d��� &�  	` &�  	` &�d��� &�d      H   ,��, $e���, $q�  	` $q�  	` $e���, $e�      H   ,��� (���� (����� (����� (���� (�      H   ,���$ $e����$ $e����� $e����� $e����$ $e�      H   ,��� &�Z��� &�d��� &�d��� &�Z��� &�Z      H   ,��� $+L��� $+V���� $+V���� $+L��� $+L      H   ,��m4 'kJ��m4 'kT��x� 'kT��x� 'kJ��m4 'kJ      H   ,��� $���� $+L  	` $+L  	` $���� $�      H   ,��[< &|��[< &���f� &���f� &|��[< &|      H   ,��� $���� $����� $����� $���� $�      H   ,��� (>D��� (I�  	` (I�  	` (>D��� (>D      H   ,��� #����� #���� #���� #����� #��      H   ,��[< &���[< &|  	` &|  	` &���[< &�      H   ,��� #�D��� #��  	` #��  	` #�D��� #�D      H   ,���$ '0����$ '0����� '0����� '0����$ '0�      H   ,��� #�:��� #�D��� #�D��� #�:��� #�:      H   ,��[< &���[< &���f� &���f� &���[< &�      H   ,��[< #X\��[< #Xf��f� #Xf��f� #X\��[< #X\      H   ,��� '����� (�  	` (�  	` '����� '��      H   ,��[< #L���[< #X\  	` #X\  	` #L���[< #L�      H   ,��, %�,��, %�6���� %�6���� %�,��, %�,      H   ,��[< #L���[< #L���f� #L���f� #L���[< #L�      H   ,��, '%��, '0�  	` '0�  	` '%��, '%      H   ,��, #��, #���� #���� #��, #      H   ,��, %�t��, %�,  	` %�,  	` %�t��, %�t      H   ,��, #T��, #  	` #  	` #T��, #T      H   ,��� (I���� (J���� (J���� (I���� (I�      H   ,��, #J��, #T���� #T���� #J��, #J      H   ,��, %�j��, %�t���� %�t���� %�j��, %�j      H   ,��� "˼��� "������ "������ "˼��� "˼      H   ,���$ '$����$ '%���� '%���� '$����$ '$�      H   ,��� "���� "˼  	` "˼  	` "���� "�      H   ,��� %����� %������ %������ %����� %��      H   ,��� "����� "����� "����� "����� "��      H   ,��� '����� '������ '������ '����� '��      H   ,��� "�l��� "�v���� "�v���� "�l��� "�l      H   ,��� %$��� %��  	` %��  	` %$��� %$      H   ,��� "y���� "�l  	` "�l  	` "y���� "y�      H   ,��� &�l��� &�v���� &�v���� &�l��� &�l      H   ,��� "y���� "y����� "y����� "y���� "y�      H   ,��� %��� %$���� %$���� %��� %      H   ,��m4 !����m4 !����x� !����x� !����m4 !��      H   ,��� (>:��� (>D���� (>D���� (>:��� (>:      H   ,��[< !���[< !��  	` !��  	` !���[< !�      H   ,��� %D���� %D����� %D����� %D���� %D�      H   ,��m4 !�
��m4 !���x� !���x� !�
��m4 !�
      H   ,��� &޴��� &�l  	` &�l  	` &޴��� &޴      H   ,��� %8���� %D�  	` %D�  	` %8���� %8�      H   ,��m4 'w��m4 'w��x� 'w��x� 'w��m4 'w      H   ,��� %8���� %8����� %8����� %8���� %8�      H   ,��� &ު��� &޴���� &޴���� &ު��� &ު      H   ,��m4 $����m4 $����x� $����x� $����m4 $��      H   ,��[< �d��[< �  	` �  	` �d��[< �d      H   ,��,  R���,  R�����  R�����  R���,  R�      H   ,��[< �Z��[< �d��f� �d��f� �Z��[< �Z      H   ,��� ����� ������ ������ ����� ��      H   ,��, ����, ������ ������ ����, ��      H   ,��� !`j��� !`t���� !`t���� !`j��� !`j      H   ,��, ���, ��  	` ��  	` ���, �      H   ,��m4 9���m4 9���x� 9���x� 9���m4 9�      H   ,��, �
��, ����� ����� �
��, �
      H   ,��,  G4��,  R�  	`  R�  	`  G4��,  G4      H   ,��� M|��� M����� M����� M|��� M|      H   ,��[< -���[< 9�  	` 9�  	` -���[< -�      H   ,��� A���� M|  	` M|  	` A���� A�      H   ,��[<  �<��[<  �F��f�  �F��f�  �<��[<  �<      H   ,��� A���� A����� A����� A���� A�      H   ,��m4 -���m4 -���x� -���x� -���m4 -�      H   ,��� ,��� 6���� 6���� ,��� ,      H   ,��,  G*��,  G4����  G4����  G*��,  G*      H   ,��� �t��� ,  	` ,  	` �t��� �t      H   ,���$ �\���$ �f���� �f���� �\���$ �\      H   ,��� �j��� �t���� �t���� �j��� �j      H   ,��� !$��� !%�  	` !%�  	` !$��� !$      H   ,��m4 z���m4 z���x� z���x� z���m4 z�      H   ,��, ���, �\  	` �\  	` ���, �      H   ,��[< n���[< z�  	` z�  	` n���[< n�      H   ,���  ����  �����  �����  ����  �      H   ,��m4 n���m4 n���x� n���x� n���m4 n�      H   ,���$ ����$ ����� ����� ����$ �      H   ,���$ 4<���$ 4F���� 4F���� 4<���$ 4<      H   ,��[<  ����[<  �<  	`  �<  	`  ����[<  ��      H   ,��, (���, 4<  	` 4<  	` (���, (�      H   ,��� ���� ����� ����� ���� �      H   ,���$ (z���$ (����� (����� (z���$ (z      H   ,���   ����  �  	`  �  	`   ����   �      H   ,��� ����� ������ ������ ����� ��      H   ,��� �T��� �  	` �  	` �T��� �T      H   ,��� �4��� ��  	` ��  	` �4��� �4      H   ,��� !%���� !%���� !%���� !%���� !%�      H   ,��� �*��� �4���� �4���� �*��� �*      H   ,��� �J��� �T���� �T���� �J��� �J      H   ,��� ����� ����� ����� ����� ��      H   ,���   ����   �����   �����   ����   �      H   ,��� ����� ��  	` ��  	` ����� ��      H   ,��� f���� f���� f���� f���� f�      H   ,��� ����� ����� ����� ����� ��      H   ,��[<  �z��[<  ����f�  ����f�  �z��[<  �z      H   ,��[< ���[< ��f� ��f� ���[< �      H   ,��� [��� f�  	` f�  	` [��� [      H   ,��[< D��[< �  	` �  	` D��[< D      H   ,���$ !�|���$ !������ !������ !�|���$ !�|      H   ,��[< :��[< D��f� D��f� :��[< :      H   ,��� �L��� �V���� �V���� �L��� �L      H   ,��, !����, !�|  	` !�|  	` !����, !��      H   ,��� Z���� [��� [��� Z���� Z�      H   ,���$ !�����$ !������ !������ !�����$ !��      H   ,��� !��� !$��� !$��� !��� !      H   ,��� !l,��� !l6���� !l6���� !l,��� !l,      H   ,��[< ���[< �&��f� �&��f� ���[< �      H   ,��� !`t��� !l,  	` !l,  	` !`t��� !`t      H   ,��� ����� �L  	` �L  	` ����� ��      H   ,��� <J��� <T���� <T���� <J��� <J      H   ,��m4 �l��m4 �v��x� �v��x� �l��m4 �l      H   ,��[< ����[< �l  	` �l  	` ����[< ��      H   ,��m4 ����m4 ����x� ����x� ����m4 ��      H   ,���$ u���$ u&���� u&���� u���$ u      H   ,��, id��, u  	` u  	` id��, id      H   ,���$ iZ���$ id���� id���� iZ���$ iZ      H   ,��� .���� .����� .����� .���� .�      H   ,��� #��� .�  	` .�  	` #��� #      H   ,��� #
��� #���� #���� #
��� #
      H   ,��� �|��� ���� ���� �|��� �|      H   ,��� ����� �|  	` �|  	` ����� ��      H   ,��� ܺ��� ����� ����� ܺ��� ܺ      H   ,��[< [���[< [���f� [���f� [���[< [�      H   ,��[< P$��[< [�  	` [�  	` P$��[< P$      H   ,��[< P��[< P$��f� P$��f� P��[< P      H   ,��, ���, ����� ����� ���, �      H   ,��, 	���, �  	` �  	` 	���, 	�      H   ,��, 	���, 	����� 	����� 	���, 	�      H   ,��� �<��� �F���� �F���� �<��� �<      H   ,��� Ä��� �<  	` �<  	` Ä��� Ä      H   ,��� �z��� Ä���� Ä���� �z��� �z      H   ,��� ����� ������ ������ ����� ��      H   ,��� }4��� ��  	` ��  	` }4��� }4      H   ,��� }*��� }4���� }4���� }*��� }*      H   ,��m4 �L��m4 �V��x� �V��x� �L��m4 �L      H   ,��[< ���[< �L  	` �L  	` ���[< �      H   ,��m4 ����m4 ���x� ���x� ����m4 ��      H   ,���$ �����$ ����� ����� �����$ ��      H   ,��, �D��, ��  	` ��  	` �D��, �D      H   ,���$ �:���$ �D���� �D���� �:���$ �:      H   ,��� o���� o����� o����� o���� o�      H   ,��� c���� o�  	` o�  	` c���� c�      H   ,��� c���� c����� c����� c���� c�      H   ,��� )\��� )f��� )f��� )\��� )\      H   ,��� ���� )\  	` )\  	` ���� �      H   ,��� ���� ���� ���� ���� �      H   ,��[< ����[< ����f� ����f� ����[< ��      H   ,��[< ���[< ��  	` ��  	` ���[< �      H   ,��[< ����[< ���f� ���f� ����[< ��      H   ,��, Vl��, Vv���� Vv���� Vl��, Vl      H   ,��, J���, Vl  	` Vl  	` J���, J�      H   ,��, J���, J����� J����� J���, J�      H   ,��� ��� &���� &���� ���       H   ,��� d���   	`   	` d��� d      H   ,��� Z��� d���� d���� Z��� Z      H   ,��� ����� ������ ������ ����� ��      H   ,��� ���� ��  	` ��  	` ���� �      H   ,��� �
��� ����� ����� �
��� �
      H   ,��m4 =,��m4 =6��x� =6��x� =,��m4 =,      H   ,��[< 1t��[< =,  	` =,  	` 1t��[< 1t      H   ,��m4 1j��m4 1t��x� 1t��x� 1j��m4 1j      H   ,��, Ԭ��, Զ���� Զ���� Ԭ��, Ԭ      H   ,��, ����, Ԭ  	` Ԭ  	` ����, ��      H   ,��, ����, ������ ������ ����, ��      H   ,��� �\��� �f���� �f���� �\��� �\      H   ,��� ����� �\  	` �\  	` ����� ��      H   ,��� ����� ������ ������ ����� ��      H   ,��� H��� H���� H���� H��� H      H   ,��� <T��� H  	` H  	` <T��� <T      H   ,��� ^z��� ^���� ^���� ^z��� ^z      H   ,��[< ݜ��[< ݦ��f� ݦ��f� ݜ��[< ݜ      H   ,��[< ����[< ݜ  	` ݜ  	` ����[< ��      H   ,��[< ����[< ����f� ����f� ����[< ��      H   ,��, �L��, �V���� �V���� �L��, �L      H   ,��, ����, �L  	` �L  	` ����, ��      H   ,��, ����, ������ ������ ����, ��      H   ,��� P���� Q���� Q���� P���� P�      H   ,��� ED��� P�  	` P�  	` ED��� ED      H   ,��� E:��� ED���� ED���� E:��� E:      H   ,��� 
���� 
����� 
����� 
���� 
�      H   ,��� ����� 
�  	` 
�  	` ����� ��      H   ,��� ����� ������ ������ ����� ��      H   ,��m4 ~��m4 ~��x� ~��x� ~��m4 ~      H   ,��[< rT��[< ~  	` ~  	` rT��[< rT      H   ,��m4 rJ��m4 rT��x� rT��x� rJ��m4 rJ      H   ,���$ 7����$ 7����� 7����� 7����$ 7�      H   ,��, ,��, 7�  	` 7�  	` ,��, ,      H   ,���$ +����$ ,���� ,���� +����$ +�      H   ,��� �l��� �v���� �v���� �l��� �l      H   ,��� ���� �l  	` �l  	` ���� �      H   ,��� ���� ����� ����� ���� �      H   ,��� ���� �&��� �&��� ���� �      H   ,��� �d��� �  	` �  	` �d��� �d      H   ,��� �Z��� �d��� �d��� �Z��� �Z      H   ,��[< |��[< ���f� ���f� |��[< |      H   ,��[< ���[< |  	` |  	` ���[< �      H   ,��[< ���[< ���f� ���f� ���[< �      H   ,��, �,��, �6���� �6���� �,��, �,      H   ,��, �t��, �,  	` �,  	` �t��, �t      H   ,��, �j��, �t���� �t���� �j��, �j      H   ,��� ����� ������ ������ ����� ��      H   ,��� �$��� ��  	` ��  	` �$��� �$      H   ,��� ���� �$���� �$���� ���� �      H   ,��� K���� K����� K����� K���� K�      H   ,��� ?���� K�  	` K�  	` ?���� ?�      H   ,��� ?���� ?����� ?����� ?���� ?�      H   ,��m4 ����m4 ����x� ����x� ����m4 ��      H   ,��[< �4��[< ��  	` ��  	` �4��[< �4      H   ,��m4 �*��m4 �4��x� �4��x� �*��m4 �*      H   ,���$ x����$ x����� x����� x����$ x�      H   ,��, l���, x�  	` x�  	` l���, l�      H   ,���$ l����$ l����� l����� l����$ l�      H   ,��� 2L��� 2V���� 2V���� 2L��� 2L      H   ,��� &���� 2L  	` 2L  	` &���� &�      H   ,��� &���� &����� &����� &���� &�      H   ,��� ����� ���� ���� ����� ��      H   ,��� �D��� ��  	` ��  	` �D��� �D      H   ,��� �:��� �D��� �D��� �:��� �:      H   ,��[< _\��[< _f��f� _f��f� _\��[< _\      H   ,��[< S���[< _\  	` _\  	` S���[< S�      H   ,��[< S���[< S���f� S���f� S���[< S�      H   ,���$ �����$ ������ ������ �����$ ��      H   ,��, �$��, ��  	` ��  	` �$��, �$      H   ,���$ ����$ �$���� �$���� ����$ �      H   ,��� ����� ������ ������ ����� ��      H   ,��� ����� ��  	` ��  	` ����� ��      H   ,��� ����� ������ ������ ����� ��      H   ,��� j<��� jF��� jF��� j<��� j<      H   ,��� ^���� j<  	` j<  	` ^���� ^�      H   ,��� ����� ������ ������ ����� ��      H   ,��m4 ����m4 ����x� ����x� ����m4 ��      H   ,��[< ���[< ��  	` ��  	` ���[< �      H   ,��m4 �
��m4 ���x� ���x� �
��m4 �
      H   ,���$ �|���$ ������ ������ �|���$ �|      H   ,��, ����, �|  	` �|  	` ����, ��      H   ,���$ �����$ ������ ������ �����$ ��      H   ,��� s,��� s6���� s6���� s,��� s,      H   ,��� gt��� s,  	` s,  	` gt��� gt      H   ,��� gj��� gt���� gt���� gj��� gj      H   ,��� ,���� ,���� ,���� ,���� ,�      H   ,��� !$��� ,�  	` ,�  	` !$��� !$      H   ,��� !��� !$��� !$��� !��� !      H   ,��[< 
�<��[< 
�F��f� 
�F��f� 
�<��[< 
�<      H   ,��[< 
����[< 
�<  	` 
�<  	` 
����[< 
��      H   ,��[< 
�z��[< 
����f� 
����f� 
�z��[< 
�z      H   ,��, 
Y���, 
Y����� 
Y����� 
Y���, 
Y�      H   ,��, 
N4��, 
Y�  	` 
Y�  	` 
N4��, 
N4      H   ,��, 
N*��, 
N4���� 
N4���� 
N*��, 
N*      H   ,��� 
���� 
����� 
����� 
���� 
�      H   ,��� 
���� 
�  	` 
�  	` 
���� 
�      H   ,��� 
���� 
����� 
����� 
���� 
�      H   ,��� 	�L��� 	�V���� 	�V���� 	�L��� 	�L      H   ,��� 	����� 	�L  	` 	�L  	` 	����� 	��      H   ,��� 	����� 	������ 	������ 	����� 	��      H   ,��m4 	@���m4 	@���x� 	@���x� 	@���m4 	@�      H   ,��[< 	4���[< 	@�  	` 	@�  	` 	4���[< 	4�      H   ,��m4 	4���m4 	4���x� 	4���x� 	4���m4 	4�      H   ,���$ �\���$ �f���� �f���� �\���$ �\      H   ,��, ���, �\  	` �\  	` ���, �      H   ,���$ ����$ ����� ����� ����$ �      H   ,��� ���� ����� ����� ���� �      H   ,��� �T��� �  	` �  	` �T��� �T      H   ,��� �J��� �T���� �T���� �J��� �J      H   ,��� m���� m���� m���� m���� m�      H   ,��� b��� m�  	` m�  	` b��� b      H   ,��� a���� b��� b��� a���� a�      H   ,��[< ���[< �&��f� �&��f� ���[< �      H   ,��[< �d��[< �  	` �  	` �d��[< �d      H   ,��[< �Z��[< �d��f� �d��f� �Z��[< �Z      H   ,��, ����, ������ ������ ����, ��      H   ,��, ���, ��  	` ��  	` ���, �      H   ,��, �
��, ����� ����� �
��, �
      H   ,��� T|��� T����� T����� T|��� T|      H   ,��� H���� T|  	` T|  	` H���� H�      H   ,��� H���� H����� H����� H���� H�      H   ,��� ,��� 6���� 6���� ,��� ,      H   ,��� t��� ,  	` ,  	` t��� t      H   ,��� j��� t���� t���� j��� j      H   ,��m4 ����m4 ����x� ����x� ����m4 ��      H   ,��[< u���[< ��  	` ��  	` u���[< u�      H   ,��m4 u���m4 u���x� u���x� u���m4 u�      H   ,��, ��, ���� ���� ��,       H   ,��, T��,   	`   	` T��, T      H   ,��, J��, T���� T���� J��, J      H   ,��� Ҽ��� ������ ������ Ҽ��� Ҽ      H   ,��� ���� Ҽ  	` Ҽ  	` ���� �      H   ,��� ����� ����� ����� ����� ��      H   ,��� �l��� �v���� �v���� �l��� �l      H   ,��� ����� �l  	` �l  	` ����� ��      H   ,��� ����� ����� ����� ����� ��      H   ,��[< !���[< "��f� "��f� !���[< !�      H   ,��[< D��[< !�  	` !�  	` D��[< D      H   ,��[< :��[< D��f� D��f� :��[< :      H   ,��, ۬��, ۶���� ۶���� ۬��, ۬      H   ,��, ����, ۬  	` ۬  	` ����, ��      H   ,��, ����, ������ ������ ����, ��      H   ,��� �\��� �f���� �f���� �\��� �\      H   ,��� ����� �\  	` �\  	` ����� ��      H   ,��� ����� ������ ������ ����� ��      H   ,��� O��� O���� O���� O��� O      H   ,��� CT��� O  	` O  	` CT��� CT      H   ,��� CJ��� CT���� CT���� CJ��� CJ      H   ,��m4 �l��m4 �v��x� �v��x� �l��m4 �l      H   ,��[< ����[< �l  	` �l  	` ����[< ��      H   ,��m4 ����m4 ����x� ����x� ����m4 ��      H   ,���$ |���$ |&���� |&���� |���$ |      H   ,��, pd��, |  	` |  	` pd��, pd      H   ,���$ pZ���$ pd���� pd���� pZ���$ pZ      H   ,��� 5���� 5����� 5����� 5���� 5�      H   ,��� *��� 5�  	` 5�  	` *��� *      H   ,��� *
��� *���� *���� *
��� *
      H   ,��� �|��� ���� ���� �|��� �|      H   ,��� ����� �|  	` �|  	` ����� ��      H   ,��� ���� ����� ����� ���� �      H   ,���$ ;<���$ ;F���� ;F���� ;<���$ ;<      H   ,��, /���, ;<  	` ;<  	` /���, /�      H   ,���$ /z���$ /����� /����� /z���$ /z      H   ,��� ����� ������ ������ ����� ��      H   ,��� �4��� ��  	` ��  	` �4��� �4      H   ,��� �*��� �4���� �4���� �*��� �*      H   ,��� ����� ����� ����� ����� ��      H   ,��� ����� ��  	` ��  	` ����� ��      H   ,��� �z��� ʄ���� ʄ���� �z��� �z      H   ,��� ����� ������ ������ ����� ��      H   ,��� �4��� ��  	` ��  	` �4��� �4      H   ,��� �*��� �4���� �4���� �*��� �*      H   ,��m4 L��m4 V��x� V��x� L��m4 L      H   ,��[<  ����[< L  	` L  	`  ����[<  ��      H   ,��m4  ����m4  ����x�  ����x�  ����m4  ��      H   ,���$  �����$  �����  �����  �����$  ��      H   ,��,  �D��,  ��  	`  ��  	`  �D��,  �D      H   ,���$  �:���$  �D����  �D����  �:���$  �:      H   ,���  v����  v�����  v�����  v����  v�      H   ,���  j����  v�  	`  v�  	`  j����  j�      H   ,���  j����  j�����  j�����  j����  j�      H   ,���  0\���  0f���  0f���  0\���  0\      H   ,���  $����  0\  	`  0\  	`  $����  $�      H   ,���  $����  $����  $����  $����  $�      H   ,�����������������������������������      H   ,  �����  �����  l����  l����  �����      H   ,��[< b���[< b���f� b���f� b���[< b�      H   ,�����������������������������������      H   ,  �����  �����  l����  l����  �����      H   ,��������������������������������      H   , oD��� oD��� z���� z���� oD���      H   ,��[< W$��[< b�  	` b�  	` W$��[< W$      H   ,�������������������������������������      H   , oD���� oD���� z����� z����� oD����      H   ,�����ռ���������������������ռ�����ռ      H   ,  V��ռ  V����  a�����  a���ռ  V��ռ      H   ,��[< W��[< W$��f� W$��f� W��[< W      H   ,�����������������������������������      H   ,  V����  V���  a����  a�����  V����      H   ,�������������������������������������      H   , ������ ������ �L���� �L���� ������      H   ,��, ���, ����� ����� ���, �      H   ,��������������������������������      H   , ����� ����� �L��� �L��� �����      H   ,���$�������$�����������������������$����      H   ,  �T����  �T����  �����  �����  �T����      H   ,��, ���, �  	` �  	` ���, �      H   ,���$���
���$�����������������
���$���
      H   ,  �T���
  �T���  ����  ����
  �T���
      H   ,��,������,����������������������,����      H   , ������ ������ ����� ����� ������      H   ,��, ���, ����� ����� ���, �      H   ,��,�����,�������������������,���      H   , ����� ����� ���� ���� �����      H   ,��m4������m4������x�������x�������m4����      H   ,  �����  �����  �\����  �\����  �����      H   ,��� �<��� �F���� �F���� �<��� �<      H   ,��m4�����m4���$��x����$��x������m4���      H   ,  ����  ����$  �\���$  �\���  ����      H   ,��[<��{���[<��{���f���{���f���{���[<��{�      H   ,��� ʄ��� �<  	` �<  	` ʄ��� ʄ      H   ,��[<��p"��[<��p,��f���p,��f���p"��[<��p"      H   , t���� t���� �l��� �l��� t����      H   , $���� $���  ����  ����� $����      H   , ������ ������ ڌ���� ڌ���� ������      H   , ���� ���� Ƽ��� Ƽ��� ����      H   , [t���� [t���� g,���� g,���� [t����      H   , $��ռ $����  �����  ���ռ $��ռ      H   , ������ ������ �|���� �|���� ������      H   , t����� t����� �l���� �l���� t�����      H   , .d��� .d��� :��� :��� .d���      H   , [t���
 [t��� g,��� g,���
 [t���
      H   , ����� �����$ �|���$ �|��� �����      H   , .d���� .d���� :���� :���� .d����      H   , B4��{� B4��{� M���{� M���{� B4��{�      H   , T��{� T��{� ��{� ��{� T��{�      H   , ������ ������ ڌ���� ڌ���� ������      H   , ����� ����� Ƽ���� Ƽ���� �����      H   , B4��p" B4��p, M���p, M���p" B4��p"      H   , T��p" T��p, ��p, ��p" T��p"      H   , 3����� 3����� ?����� ?����� 3�����      H   , 	������ 	������ 	������ 	������ 	������      H   , z$���� z$���� ������ ������ z$����      H   , 
9D���� 
9D���� 
D����� 
D����� 
9D����      H   , M���� M���� X����� X����� M����      H   , �D��ռ �D���� ������ ����ռ �D��ռ      H   , �d��ռ �d���� ����� ���ռ �d��ռ      H   , ������ ������ ������ ������ ������      H   , z$��� z$��� ����� ����� z$���      H   , 
9D��� 
9D��� 
D���� 
D���� 
9D���      H   , 3���� 3���� ?���� ?���� 3����      H   , 	����� 	����� 	����� 	����� 	�����      H   , M���� M���� X����� X����� M����      H   , `����� `����� l����� l����� `�����      H   , 	 ���� 	 ���� 	+����� 	+����� 	 ����      H   , ������ ������ ������ ������ ������      H   , ����� ����� �<���� �<���� �����      H   , ����� ����� &L���� &L���� �����      H   , ٴ���� ٴ���� �l���� �l���� ٴ����      H   , `���� `����$ l����$ l���� `����      H   , 	 ��� 	 ���$ 	+����$ 	+���� 	 ���      H   , �D���� �D��� ����� ������ �D����      H   , �d���� �d��� ���� ����� �d����      H   , 	������ 	������ 	�\���� 	�\���� 	������      H   , �t��{� �t��{� �,��{� �,��{� �t��{�      H   , 
���{� 
���{� 
�L��{� 
�L��{� 
���{�      H   , ���� ���� �<��� �<��� ����      H   , ����
 ���� &L��� &L���
 ����
      H   , ٴ���
 ٴ��� �l��� �l���
 ٴ���
      H   , 	����� 	����� 	�\��� 	�\��� 	�����      H   , �t��p" �t��p, �,��p, �,��p" �t��p"      H   , 
���p" 
���p, 
�L��p, 
�L��p" 
���p"      H   , ���� ���� ����� ����� ����      H   , �$��� �$��� ����� ����� �$���      H   , 4���� 4���� ����� ����� 4����      H   , �T���� �T���� ����� ����� �T����      H   , �t���� �t���� �,���� �,���� �t����      H   , �����
 ����� ����� �����
 �����
      H   , W����
 W���� c���� c����
 W����
      H   , ���
 ��� "���� "����
 ���
      H   , �4���
 �4��� ����� �����
 �4���
      H   , R����� R���� ^<��� ^<���� R�����      H   , ����� ���� \��� \���� �����      H   , ������ ����� �|��� �|���� ������      H   , ������ ����� ����� ������ ������      H   , I����� I����� UL���� UL���� I�����      H   , �d���� �d���� ���� ���� �d����      H   , ������ ������ �<���� �<���� ������      H   , v����� v����� �\���� �\���� v�����      H   , 5����� 5����� A|���� A|���� 5�����      H   , ����� ����� l���� l���� �����      H   , �T���� �T���� ����� ����� �T����      H   , k����� k����� w|���� w|���� k�����      H   , *����� *����� 6����� 6����� *�����      H   , ����� ����� ������ ������ �����      H   , q4���� q4���� |����� |����� q4����      H   , �d��� �d��� ��� ��� �d���      H   , ����� ����� �<��� �<��� �����      H   , v���� v���� �\��� �\��� v����      H   , 5���� 5���� A|��� A|��� 5����      H   , 0T���� 0T���� <���� <���� 0T����      H   , �t���� �t���� �,���� �,���� �t����      H   , ����� ����� ������ ������ �����      H   , �$���� �$���� ������ ������ �$����      H   , �t���� �t���� �,���� �,���� �t����      H   , �$���� �$���� ������ ������ �$����      H   , �D���� �D���� ������ ������ �D����      H   , ]d���� ]d���� i���� i���� ]d����      H   , ����� ����� (<���� (<���� �����      H   , I����� I����� UL���� UL���� I�����      H   , ����� ����� l���� l���� �����      H   , 4���� 4���� ����� ����� 4����      H   , ���� ���� ����� ����� ����      H   , q4��� q4��� |���� |���� q4���      H   , 0T��� 0T��� <��� <��� 0T���      H   , �$��� �$���$ �����$ ����� �$���      H   , �D��� �D���$ �����$ ����� �D���      H   , ]d��� ]d���$ i���$ i��� ]d���      H   , ���� ����$ (<���$ (<��� ����      H   , �t��� �t��� �,��� �,��� �t���      H   , k���� k���� w|��� w|��� k����      H   , R���ռ R����� ^<���� ^<��ռ R���ռ      H   , ���ռ ����� \���� \��ռ ���ռ      H   , ����ռ ������ �|���� �|��ռ ����ռ      H   , >���{� >���{� Jl��{� Jl��{� >���{�      H   , ����{� ����{� 	���{� 	���{� ����{�      H   , ����{� ����{� Ȭ��{� Ȭ��{� ����{�      H   , |��{� |��{� ����{� ����{� |��{�      H   , ����ռ ������ ������ ����ռ ����ռ      H   , ������ ������ ������ ������ ������      H   , W����� W����� c����� c����� W�����      H   , ���� ���� "����� "����� ����      H   , �4���� �4���� ������ ������ �4����      H   , *���� *���� 6���� 6���� *����      H   , >���p" >���p, Jl��p, Jl��p" >���p"      H   , ����p" ����p, 	���p, 	���p" ����p"      H   , ����p" ����p, Ȭ��p, Ȭ��p" ����p"      H   , |��p" |��p, ����p, ����p" |��p"      H   , -� � -� � -� � -� � -� �      H   , ,�� J� ,�� Vl -� Vl -� J� ,�� J�      H   , ,�� u ,�� u& ,�� u& ,�� u ,�� u      H   , -� J� -� J� -� J� -� J� -� J�      H   , ,�� 	� ,�� � -� � -� 	� ,�� 	�      H   , ,��  ,�� & ,� & ,�  ,��       H   , ,�  H ,�  H ,Ÿ H ,Ÿ H ,�  H      H   , ,�� d ,��  ,�  ,� d ,�� d      H   , -� 	� -� 	� -� 	� -� 	� -� 	�      H   , ,�� Z ,�� d ,� d ,� Z ,�� Z      H   , ,�� id ,�� u -� u -� id ,�� id      H   , ,�  �� ,�  �� ,Ÿ �� ,Ÿ �� ,�  ��      H   , ,�� �< ,�� �F ,� �F ,� �< ,�� �<      H   , ,�� � ,�� �� ,Ÿ �� ,Ÿ � ,�� �      H   , ,�� �\ ,�� �f ,� �f ,� �\ ,�� �\      H   , ,�  �
 ,�  � ,Ÿ � ,Ÿ �
 ,�  �
      H   , ,�� Ä ,�� �< ,� �< ,� Ä ,�� Ä      H   , -� =, -� =6 -� =6 -� =, -� =,      H   , ,�� iZ ,�� id ,�� id ,�� iZ ,�� iZ      H   , ,�� 1t ,�� =, -1� =, -1� 1t ,�� 1t      H   , ,�� �z ,�� Ä ,� Ä ,� �z ,�� �z      H   , -� 1j -� 1t -� 1t -� 1j -� 1j      H   , ,�� <T ,�� H ,Ÿ H ,Ÿ <T ,�� <T      H   , ,�  �� ,�  �� ,Ÿ �� ,Ÿ �� ,�  ��      H   , ,�� .� ,�� .� ,װ .� ,װ .� ,�� .�      H   , ,�� }4 ,�� �� ,Ÿ �� ,Ÿ }4 ,�� }4      H   , -� Ԭ -� Զ -� Զ -� Ԭ -� Ԭ      H   , ,�  }* ,�  }4 ,Ÿ }4 ,Ÿ }* ,�  }*      H   , ,�� # ,�� .� ,� .� ,� # ,�� #      H   , -� �L -� �V -� �V -� �L -� �L      H   , ,�  <J ,�  <T ,Ÿ <T ,Ÿ <J ,�  <J      H   , ,�� � ,�� �L -1� �L -1� � ,�� �      H   , ,�� #
 ,�� # ,װ # ,װ #
 ,�� #
      H   , -� �� -� � -� � -� �� -� ��      H   , ,�� �� ,�� �\ ,� �\ ,� �� ,�� ��      H   , ,�� �� ,�� � ,�� � ,�� �� ,�� ��      H   , ,� �| ,� � ,�� � ,�� �| ,� �|      H   , ,�� �D ,�� �� -� �� -� �D ,�� �D      H   , -� �l -� �v -� �v -� �l -� �l      H   , ,�� �: ,�� �D ,�� �D ,�� �: ,�� �:      H   , ,�� �� ,�� �| ,Ÿ �| ,Ÿ �� ,�� ��      H   , ,�� o� ,�� o� ,װ o� ,װ o� ,�� o�      H   , -� �� -� �� -� �� -� �� -� ��      H   , ,�� c� ,�� o� ,� o� ,� c� ,�� c�      H   , ,� ܺ ,� �� ,�� �� ,�� ܺ ,� ܺ      H   , ,�� c� ,�� c� ,װ c� ,װ c� ,�� c�      H   , ,�� �� ,�� �l -1� �l -1� �� ,�� ��      H   , ,� )\ ,� )f ,�� )f ,�� )\ ,� )\      H   , -%� [� -%� [� -1� [� -1� [� -%� [�      H   , ,�� � ,�� )\ ,Ÿ )\ ,Ÿ � ,�� �      H   , ,�� �� ,�� �� ,� �� ,� �� ,�� ��      H   , ,� � ,� � ,�� � ,�� � ,� �      H   , ,�� P$ ,�� [� -1� [� -1� P$ ,�� P$      H   , -%� �� -%� �� -1� �� -1� �� -%� ��      H   , -� �� -� �� -� �� -� �� -� ��      H   , ,�� � ,�� �� -1� �� -1� � ,�� �      H   , -%� P -%� P$ -1� P$ -1� P -%� P      H   , -%� �� -%� � -1� � -1� �� -%� ��      H   , ,�� �� ,�� Ԭ -� Ԭ -� �� ,�� ��      H   , -� Vl -� Vv -� Vv -� Vl -� Vl      H   , -� �� -� �� -� �� -� �� -� ��      H   , ,� ^z ,� ^� ,�� ^� ,�� ^z ,� ^z      H   , ,�� &� ,�� &� ,װ &� ,װ &� ,�� &�      H   , -%� ݜ -%� ݦ -1� ݦ -1� ݜ -%� ݜ      H   , -� �j -� �t -� �t -� �j -� �j      H   , ,�� �� ,�� ݜ -1� ݜ -1� �� ,�� ��      H   , ,� �� ,� � ,�� � ,�� �� ,� ��      H   , -%� �� -%� �� -1� �� -1� �� -%� ��      H   , ,�� �4 ,�� �� -1� �� -1� �4 ,�� �4      H   , -� �L -� �V -� �V -� �L -� �L      H   , ,�� �D ,�� �� ,Ÿ �� ,Ÿ �D ,�� �D      H   , ,�� �� ,�� �L -� �L -� �� ,�� ��      H   , ,�  K� ,�  K� ,Ÿ K� ,Ÿ K� ,�  K�      H   , -� �� -� �� -� �� -� �� -� ��      H   , ,� �: ,� �D ,�� �D ,�� �: ,� �:      H   , ,�� P� ,�� Q ,� Q ,� P� ,�� P�      H   , -� �* -� �4 -� �4 -� �* -� �*      H   , ,�� ED ,�� P� ,� P� ,� ED ,�� ED      H   , -%� _\ -%� _f -1� _f -1� _\ -%� _\      H   , ,�� E: ,�� ED ,� ED ,� E: ,�� E:      H   , ,�� �$ ,�� �� ,� �� ,� �$ ,�� �$      H   , ,�  
� ,�  
� ,Ÿ 
� ,Ÿ 
� ,�  
�      H   , ,�� S� ,�� _\ -1� _\ -1� S� ,�� S�      H   , ,�� �� ,�� 
� ,Ÿ 
� ,Ÿ �� ,�� ��      H   , ,�� x� ,�� x� ,�� x� ,�� x� ,�� x�      H   , ,�  �� ,�  �� ,Ÿ �� ,Ÿ �� ,�  ��      H   , -%� S� -%� S� -1� S� -1� S� -%� S�      H   , -� ~ -� ~ -� ~ -� ~ -� ~      H   , ,�� ?� ,�� K� ,Ÿ K� ,Ÿ ?� ,�� ?�      H   , ,�� rT ,�� ~ -1� ~ -1� rT ,�� rT      H   , ,�� �� ,�� �� ,�� �� ,�� �� ,�� ��      H   , -� rJ -� rT -� rT -� rJ -� rJ      H   , ,�� l� ,�� x� -� x� -� l� ,�� l�      H   , ,�� 7� ,�� 7� ,�� 7� ,�� 7� ,�� 7�      H   , ,�� �$ ,�� �� -� �� -� �$ ,�� �$      H   , ,�� , ,�� 7� -� 7� -� , ,�� ,      H   , ,�� �� ,�� �� ,� �� ,� �� ,�� ��      H   , ,�� +� ,�� , ,�� , ,�� +� ,�� +�      H   , ,�� � ,�� �$ ,�� �$ ,�� � ,�� �      H   , ,�� �l ,�� �v ,װ �v ,װ �l ,�� �l      H   , ,�� l� ,�� l� ,�� l� ,�� l� ,�� l�      H   , ,�� � ,�� �l ,� �l ,� � ,�� �      H   , ,�� �� ,�� �� ,װ �� ,װ �� ,�� ��      H   , ,�� � ,�� � ,װ � ,װ � ,�� �      H   , ,�  ?� ,�  ?� ,Ÿ ?� ,Ÿ ?� ,�  ?�      H   , ,� � ,� �& ,�� �& ,�� � ,� �      H   , ,�� �� ,�� �� ,� �� ,� �� ,�� ��      H   , ,�� �d ,�� � ,Ÿ � ,Ÿ �d ,�� �d      H   , ,�� 2L ,�� 2V ,װ 2V ,װ 2L ,�� 2L      H   , ,� �Z ,� �d ,�� �d ,�� �Z ,� �Z      H   , ,�� �� ,�� �� ,װ �� ,װ �� ,�� ��      H   , -%� | -%� � -1� � -1� | -%� |      H   , ,�� � ,�� �$ ,� �$ ,� � ,�� �      H   , ,�� � ,�� | -1� | -1� � ,�� �      H   , ,� j< ,� jF ,�� jF ,�� j< ,� j<      H   , -%� � -%� � -1� � -1� � -%� �      H   , ,�� &� ,�� 2L ,� 2L ,� &� ,�� &�      H   , -� �, -� �6 -� �6 -� �, -� �,      H   , ,�� ^� ,�� j< ,Ÿ j< ,Ÿ ^� ,�� ^�      H   , ,�� �t ,�� �, -� �, -� �t ,�� �t      H   , �T���� �T���� ����� ����� �T����      H   , Tt���� Tt���� `,���� `,���� Tt����      H   , ����� ����� L���� L���� �����      H   , Ҵ���� Ҵ���� �l���� �l���� Ҵ����      H   , !������ !������ !������ !������ !������      H   , �d��ռ �d���� ����� ���ռ �d��ռ      H   , !K���ռ !K����� !W<���� !W<��ռ !K���ռ      H   , 'd��� 'd��� 3��� 3��� 'd���      H   , ���� ���� �<��� �<��� ����      H   , ����� ����� �\��� �\��� �����      H   , �T���
 �T��� ���� ����
 �T���
      H   , Tt���
 Tt��� `,��� `,���
 Tt���
      H   , ����
 ���� L��� L���
 ����
      H   , Ҵ���
 Ҵ��� �l��� �l���
 Ҵ���
      H   , !�����
 !����� !����� !�����
 !�����
      H   , ������ ������ ������ ������ ������      H   , F���� F���� Q����� Q����� F����      H   , O���� O��� Z���� Z����� O����      H   , $���� $��� ���� ����� $����      H   , �D���� �D��� ����� ������ �D����      H   , ������ ������  �����  ����� ������      H   , ����� ����� ������ ������ �����      H   , s$���� s$���� ~����� ~����� s$����      H   ,  2D����  2D����  =�����  =�����  2D����      H   , �d���� �d��� ���� ����� �d����      H   , !K����� !K���� !W<��� !W<���� !K�����      H   , !4���� !4���� !����� !����� !4����      H   , ������ ������ ������ ������ ������      H   , F���� F���� Q����� Q����� F����      H   , ����� �����  ����  ���� �����      H   , ���� ���� ����� ����� ����      H   , s$��� s$��� ~���� ~���� s$���      H   ,  2D���  2D���  =����  =����  2D���      H   , hD���� hD���� s����� s����� hD����      H   , 'd���� 'd���� 3���� 3���� 'd����      H   , ������ ������ �L���� �L���� ������      H   , m����� m����� yl���� yl���� m�����      H   , ۤ���� ۤ���� �\���� �\���� ۤ����      H   , ������ ������ �|���� �|���� ������      H   , Y����� Y����� e����� e����� Y�����      H   , ���� ���� $����� $����� ����      H   , ,����� ,����� 8����� 8����� ,�����      H   , ������ ������ ������ ������ ������      H   , ����� ����� �<���� �<���� �����      H   , ������ ������ �\���� �\���� ������      H   , !4���� !4���� !����� !����� !4����      H   , ۤ��� ۤ���$ �\���$ �\��� ۤ���      H   , ����� �����$ �|���$ �|��� �����      H   , Y���� Y����$ e����$ e���� Y����      H   , ��� ���$ $����$ $���� ���      H   , ������ ������ ӌ���� ӌ���� ������      H   , ������ ������ ӌ���� ӌ���� ������      H   , ����� ����� �L��� �L��� �����      H   , m���� m���� yl��� yl��� m����      H   , ,���� ,���� 8���� 8���� ,����      H   , ;4��{� ;4��{� F���{� F���{� ;4��{�      H   , �T��{� �T��{� ��{� ��{� �T��{�      H   , �t��{� �t��{� �,��{� �,��{� �t��{�      H   ,  x���{�  x���{�  �L��{�  �L��{�  x���{�      H   , ����� ����� ����� ����� �����      H   , hD��� hD��� s���� s���� hD���      H   , O��ռ O���� Z����� Z���ռ O��ռ      H   , $��ռ $���� ����� ���ռ $��ռ      H   , �D��ռ �D���� ������ ����ռ �D��ռ      H   , ;4��p" ;4��p, F���p, F���p" ;4��p"      H   , �T��p" �T��p, ��p, ��p" �T��p"      H   , �t��p" �t��p, �,��p, �,��p" �t��p"      H   ,  x���p"  x���p,  �L��p,  �L��p"  x���p"      H   , ,�� 
� ,�� 
� ,� 
� ,� 
� ,�� 
�      H   , ,�� 
� ,�� 
� ,� 
� ,� 
� ,�� 
�      H   , ,�  	�L ,�  	�V ,Ÿ 	�V ,Ÿ 	�L ,�  	�L      H   , ,�� 	�� ,�� 	�L ,Ÿ 	�L ,Ÿ 	�� ,�� 	��      H   , ,�� Ҽ ,�� �� ,� �� ,� Ҽ ,�� Ҽ      H   , ,�� � ,�� Ҽ ,� Ҽ ,� � ,�� �      H   , ,�� �� ,�� � ,� � ,� �� ,�� ��      H   , ,�  	�� ,�  	�� ,Ÿ 	�� ,Ÿ 	�� ,�  	��      H   , -� 	@� -� 	@� -� 	@� -� 	@� -� 	@�      H   , ,�  �l ,�  �v ,Ÿ �v ,Ÿ �l ,�  �l      H   , ,�� 	4� ,�� 	@� -1� 	@� -1� 	4� ,�� 	4�      H   , -� 	4� -� 	4� -� 	4� -� 	4� -� 	4�      H   , ,�� �� ,�� �l ,Ÿ �l ,Ÿ �� ,�� ��      H   , ,�� �\ ,�� �f ,�� �f ,�� �\ ,�� �\      H   , ,�  �� ,�  �� ,Ÿ �� ,Ÿ �� ,�  ��      H   , ,�� � ,�� �\ -� �\ -� � ,�� �      H   , ,�� � ,�� � ,�� � ,�� � ,�� �      H   , ,�� � ,�� � ,װ � ,װ � ,�� �      H   , ,�� �T ,�� � ,� � ,� �T ,�� �T      H   , ,�� �J ,�� �T ,װ �T ,װ �J ,�� �J      H   , -� �� -� �� -� �� -� �� -� ��      H   , ,�� � ,�� �� -1� �� -1� � ,�� �      H   , ,� m� ,� m� ,�� m� ,�� m� ,� m�      H   , ,�� b ,�� m� ,Ÿ m� ,Ÿ b ,�� b      H   , -� �
 -� � -� � -� �
 -� �
      H   , ,� a� ,� b ,�� b ,�� a� ,� a�      H   , -%� � -%� �& -1� �& -1� � -%� �      H   , ,�� �| ,�� �� ,�� �� ,�� �| ,�� �|      H   , ,�� �d ,�� � -1� � -1� �d ,�� �d      H   , -%� �Z -%� �d -1� �d -1� �Z -%� �Z      H   , -� �� -� �� -� �� -� �� -� ��      H   , ,�� � ,�� �� -� �� -� � ,�� �      H   , -� �
 -� � -� � -� �
 -� �
      H   , ,�� �� ,�� �| -� �| -� �� ,�� ��      H   , ,�� �� ,�� �� ,�� �� ,�� �� ,�� ��      H   , ,�� T| ,�� T� ,� T� ,� T| ,�� T|      H   , ,�� s, ,�� s6 ,װ s6 ,װ s, ,�� s,      H   , ,�� H� ,�� T| ,� T| ,� H� ,�� H�      H   , ,�� H� ,�� H� ,� H� ,� H� ,�� H�      H   , ,�� gt ,�� s, ,� s, ,� gt ,�� gt      H   , ,�  , ,�  6 ,Ÿ 6 ,Ÿ , ,�  ,      H   , ,�� t ,�� , ,Ÿ , ,Ÿ t ,�� t      H   , ,�� gj ,�� gt ,װ gt ,װ gj ,�� gj      H   , ,�  j ,�  t ,Ÿ t ,Ÿ j ,�  j      H   , -� �� -� �� -� �� -� �� -� ��      H   , ,�� u� ,�� �� -1� �� -1� u� ,�� u�      H   , -� u� -� u� -� u� -� u� -� u�      H   , ,� ,� ,� ,� ,�� ,� ,�� ,� ,� ,�      H   , ,�� !$ ,�� ,� ,Ÿ ,� ,Ÿ !$ ,�� !$      H   , ,� ! ,� !$ ,�� !$ ,�� ! ,� !      H   , -%� 
�< -%� 
�F -1� 
�F -1� 
�< -%� 
�<      H   , ,�� 
�� ,�� 
�< -1� 
�< -1� 
�� ,�� 
��      H   , -�  -�  -�  -�  -�       H   , -%� 
�z -%� 
�� -1� 
�� -1� 
�z -%� 
�z      H   , ,�� T ,��  -�  -� T ,�� T      H   , -� 
Y� -� 
Y� -� 
Y� -� 
Y� -� 
Y�      H   , ,�� 
N4 ,�� 
Y� -� 
Y� -� 
N4 ,�� 
N4      H   , -� J -� T -� T -� J -� J      H   , -� 
N* -� 
N4 -� 
N4 -� 
N* -� 
N*      H   , ,�� 
� ,�� 
� ,� 
� ,� 
� ,�� 
�      H   , '���
 '��� '���� '����
 '���
      H   , "�d��� "�d��� "���� "���� "�d���      H   , %����� %����� %�<��� %�<��� %�����      H   , "d���� "d���� "p|��� "p|��� "d����      H   , &�t���� &�t���� &�,���� &�,���� &�t����      H   , "d����� "d����� "p|���� "p|���� "d�����      H   , %#���� %#���� %/���� %/���� %#����      H   , %#����� %#����� %/����� %/����� %#�����      H   , #�T���� #�T���� #����� #����� #�T����      H   , $P����� $P����� $\����� $\����� $P�����      H   , !�$���� !�$���� !������ !������ !�$����      H   , $�D���� $�D���� $������ $������ $�D����      H   , 'Vd���� 'Vd���� 'b���� 'b���� 'Vd����      H   , '���� '���� '����� '����� '����      H   , "���� "���� "����� "����� "����      H   , %j4��� %j4��� %u���� %u���� %j4���      H   , "�d���� "�d���� "����� "����� "�d����      H   , !�$��� !�$���$ !�����$ !����� !�$���      H   , $�D��� $�D���$ $�����$ $����� $�D���      H   , 'Vd��� 'Vd���$ 'b���$ 'b��� 'Vd���      H   , %������ %������ %�<���� %�<���� %������      H   , $
���ռ $
����� $\���� $\��ռ $
���ռ      H   , &����ռ &������ &�|���� &�|��ռ &����ռ      H   , #7���{� #7���{� #Cl��{� #Cl��{� #7���{�      H   , %����{� %����{� &���{� &���{� %����{�      H   , $
����� $
���� $\��� $\���� $
�����      H   , &������ &����� &�|��� &�|���� &������      H   , #�T���� #�T���� #����� #����� #�T����      H   , "����� "����� "������ "������ "�����      H   , &�t���� &�t���� &�,���� &�,���� &�t����      H   , %j4���� %j4���� %u����� %u����� %j4����      H   , $P����
 $P���� $\���� $\����
 $P����
      H   , #7���p" #7���p, #Cl��p, #Cl��p" #7���p"      H   , %����p" %����p, &���p, &���p" %����p"      H   , ,�� CT ,�� O ,Ÿ O ,Ÿ CT ,�� CT      H   , ,�� 5� ,�� 5� ,װ 5� ,װ 5� ,�� 5�      H   , ,� �| ,� � ,�� � ,�� �| ,� �|      H   , ,�� | ,�� |& ,�� |& ,�� | ,�� |      H   , ,�  O ,�  O ,Ÿ O ,Ÿ O ,�  O      H   , ,�� �\ ,�� �f ,� �f ,� �\ ,�� �\      H   , ,�� ;< ,�� ;F ,�� ;F ,�� ;< ,�� ;<      H   , ,�� �� ,�� �� ,� �� ,� �� ,�� ��      H   , ,�� *
 ,�� * ,װ * ,װ *
 ,�� *
      H   , ,�� /� ,�� ;< -� ;< -� /� ,�� /�      H   , ,�� /z ,�� /� ,�� /� ,�� /z ,�� /z      H   , ,�� �� ,�� �� ,װ �� ,װ �� ,�� ��      H   , ,�� �4 ,�� �� ,� �� ,� �4 ,�� �4      H   , ,�� �� ,�� �| ,Ÿ �| ,Ÿ �� ,�� ��      H   , ,�� �* ,�� �4 ,װ �4 ,װ �* ,�� �*      H   , ,�� pd ,�� | -� | -� pd ,�� pd      H   , -� �� -� �� -� �� -� �� -� ��      H   , ,� � ,� �� ,�� �� ,�� � ,� �      H   , ,�  CJ ,�  CT ,Ÿ CT ,Ÿ CJ ,�  CJ      H   , ,� �� ,� �� ,�� �� ,�� �� ,� ��      H   , ,�� �� ,�� �� ,Ÿ �� ,Ÿ �� ,�� ��      H   , ,�� �� ,�� �l -1� �l -1� �� ,�� ��      H   , ,� �� ,� �� ,�� �� ,�� �� ,� ��      H   , ,�� * ,�� 5� ,� 5� ,� * ,�� *      H   , -%� !� -%� " -1� " -1� !� -%� !�      H   , ,�� pZ ,�� pd ,�� pd ,�� pZ ,�� pZ      H   , -� �l -� �v -� �v -� �l -� �l      H   , ,�� D ,�� !� -1� !� -1� D ,�� D      H   , -%� : -%� D -1� D -1� : -%� :      H   , -� ۬ -� ۶ -� ۶ -� ۬ -� ۬      H   , ,�� �� ,�� ۬ -� ۬ -� �� ,�� ��      H   , -� �� -� �� -� �� -� �� -� ��      H   , ,�� �� ,�� �\ ,� �\ ,� �� ,�� ��      H   , )�4���� )�4���� )������ )������ )�4����      H   , )�4���
 )�4��� )����� )�����
 )�4���
      H   , )����ռ )������ )������ )����ռ )����ռ      H   , )B����� )B����� )NL���� )NL���� )B�����      H   , *���� *����$ *!<���$ *!<��� *����      H   , (����{� (����{� (����{� (����{� (����{�      H   , )������ )����� )����� )������ )������      H   , ()T��� ()T��� (5��� (5��� ()T���      H   , (o����� (o����� ({\���� ({\���� (o�����      H   , '����� '����� '����� '����� '�����      H   , ()T���� ()T���� (5���� (5���� ()T����      H   , (o���� (o���� ({\��� ({\��� (o����      H   , '���� '���� '���� '���� '����      H   , *����� *����� *!<���� *!<���� *�����      H   , )B����� )B����� )NL���� )NL���� )B�����      H   , (����p" (����p, (����p, (����p" (����p"      H   , ,�  �* ,�  �4 ,Ÿ �4 ,Ÿ �* ,�  �*      H   , +.����� +.����� +:|���� +:|���� +.�����      H   , -%� W -%� W$ -1� W$ -1� W -%� W      H   , ,��  j� ,��  j� ,װ  j� ,װ  j� ,��  j�      H   , ,�� W$ ,�� b� -1� b� -1� W$ ,�� W$      H   , ,�� ʄ ,�� �< ,� �< ,� ʄ ,�� ʄ      H   , ,�  $� ,�  $� ,��  $� ,��  $� ,�  $�      H   , ,��  �� ,��  � ,��  � ,��  �� ,��  ��      H   , ,����� ,����� ,������ ,������ ,�����      H   , -� � -� � -� � -� � -� �      H   , -����� -����� -����� -����� -�����      H   , ,��  �D ,��  �� -�  �� -�  �D ,��  �D      H   , +.���� +.���� +:|��� +:|��� +.����      H   , -���� -���� -���� -���� -����      H   , -���� -����$ -����$ -���� -����      H   , *�t���� *�t���� *�,���� *�,���� *�t����      H   , ,�  0\ ,�  0f ,��  0f ,��  0\ ,�  0\      H   , ,�� � ,�� � -� � -� � ,�� �      H   , ,������ ,������ ,������ ,������ ,������      H   , ,������ ,������ ,����� ,����� ,������      H   , ,�  �� ,�  �� ,Ÿ �� ,Ÿ �� ,�  ��      H   , ,��  v� ,��  v� ,װ  v� ,װ  v� ,��  v�      H   , ,H���� ,H��� ,S���� ,S����� ,H����      H   , ,����� ,����� ,l���� ,l���� ,�����      H   , ,����� ,����� ,������ ,������ ,�����      H   , ,H��ռ ,H���� ,S����� ,S���ռ ,H��ռ      H   , ,����ռ ,������ ,װ���� ,װ��ռ ,����ռ      H   , *�$���� *�$���� *������ *������ *�$����      H   , ,�����
 ,����� ,����� ,�����
 ,�����
      H   , ,� ���� ,� ���� ,Ÿ���� ,Ÿ���� ,� ����      H   , ,�� �z ,�� ʄ ,� ʄ ,� �z ,�� �z      H   , +u��{� +u��{� +����{� +����{� +u��{�      H   , -%���{� -%���{� -1���{� -1���{� -%���{�      H   , ,��  �: ,��  �D ,��  �D ,��  �: ,��  �:      H   , ,�� �4 ,�� �� ,Ÿ �� ,Ÿ �4 ,�� �4      H   , -�  �� -�  �� -�  �� -�  �� -�  ��      H   , *�t��� *�t��� *�,��� *�,��� *�t���      H   , ,������ ,����� ,װ��� ,װ���� ,������      H   , ,����� ,����� ,���� ,���� ,�����      H   , -%� b� -%� b� -1� b� -1� b� -%� b�      H   , -� � -� � -� � -� � -� �      H   , -����� -����� -����� -����� -�����      H   , ,����� ,����� ,l���� ,l���� ,�����      H   , ,�� �< ,�� �F ,� �F ,� �< ,�� �<      H   , *�$��� *�$��� *����� *����� *�$���      H   , ,��  �� ,�� L -1� L -1�  �� ,��  ��      H   , -� L -� V -� V -� L -� L      H   , ,� ��� ,� ��� ,Ÿ��� ,Ÿ��� ,� ���      H   , ,��  $� ,��  0\ ,Ÿ  0\ ,Ÿ  $� ,��  $�      H   , ,��  j� ,��  v� ,�  v� ,�  j� ,��  j�      H   , +u��p" +u��p, +����p, +����p" +u��p"      H   , -%���p" -%���p, -1���p, -1���p" -%���p"      Q   , +� @� +� 2t )`� 2t )`� @� +� @�      F   ,���@ ִ���@ �d  	` �d  	` ִ���@ ִ      F   , ,�� 'Ѭ ,�� '�\ ,�  '�\ ,�  'Ѭ ,�� 'Ѭ      F   , ,�� +f ,�� +j� ,�  +j� ,�  +f ,�� +f      F   , ,�� .�| ,�� .�, ,�  .�, ,�  .�| ,�� .�|      F   , ,�� 2�� ,�� 2�� ,�  2�� ,�  2�� ,�� 2��      F   , ,�� $=D ,�� $A� ,�  $A� ,�  $=D ,�� $=D      F   , ,�� t ,�� $ ,�  $ ,�  t ,�� t      F   , ,��  �� ,��  �� ,�   �� ,�   �� ,��  ��      F   , ,�� %!� ,�� %&d ,�  %&d ,�  %!� ,�� %!�      F   , ,�� (�� ,�� (�t ,�  (�t ,�  (�� ,�� (��      F   , ,�� ,M, ,�� ,Q� ,�  ,Q� ,�  ,M, ,�� ,M,      F   , ,�� /� ,�� /�D ,�  /�D ,�  /� ,�� /�      F   , ,�� 3u� ,�� 3z� ,�  3z� ,�  3u� ,�� 3u�      F   , ,�� �� ,�� �� ,�  �� ,�  �� ,�� ��      F   , ,�� !�L ,�� !�� ,�  !�� ,�  !�L ,�� !�L      F   , ,�� &�< ,�� &�� ,�  &�� ,�  &�< ,�� &�<      F   , ,�� *�� ,�� *�T ,�  *�T ,�  *�� ,�� *��      F   , ,�� . ,�� .� ,�  .� ,�  . ,�� .      F   , ,�� 1�t ,�� 1�$ ,�  1�$ ,�  1�t ,�� 1�t      F   , ,�� 5>� ,�� 5C� ,�  5C� ,�  5>� ,�� 5>�      F   , ,�� 0 ,�� 4� ,�  4� ,�  0 ,�� 0      F   , ,�� �l ,�� � ,�  � ,�  �l ,�� �l      F   , ,�� #X� ,�� #]� ,�  #]� ,�  #X� ,�� #X�      F   , ,�� &� ,�� &| ,�  &| ,�  &� ,�� &�      F   , ,�� )�4 ,�� )�� ,�  )�� ,�  )�4 ,�� )�4      F   , ,�� -1� ,�� -6L ,�  -6L ,�  -1� ,�� -1�      F   , ,�� 0� ,�� 0ʴ ,�  0ʴ ,�  0� ,�� 0�      F   , ,�� 4Zl ,�� 4_ ,�  4_ ,�  4Zl ,�� 4Zl      F   , ,�� K� ,�� PD ,�  PD ,�  K� ,�� K�      F   , ,�� �� ,�� � ,�  � ,�  �� ,�� ��      F   , ,�� "td ,�� "y ,�  "y ,�  "td ,�� "td      F   ,���@ 4
����@ 4l  	` 4l  	` 4
����@ 4
�      F   ,���@ 1�D���@ 1��  	` 1��  	` 1�D���@ 1�D      F   ,���@ -v����@ -{\  	` -{\  	` -v����@ -v�      F   ,���@ )����@ )l  	` )l  	` )����@ )�      F   ,���@ $�$���@ $��  	` $��  	` $�$���@ $�$      F   ,���@  Q4���@  U�  	`  U�  	`  Q4���@  Q4      F   ,���@ ����@ �L  	` �L  	` ����@ �      F   ,���@ /�����@ /�|  	` /�|  	` /�����@ /��      F   ,���@ +F4���@ +J�  	` +J�  	` +F4���@ +F4      F   ,���@ &�D���@ &��  	` &��  	` &�D���@ &�D      F   ,���@ "�����@ "�\  	` "�\  	` "�����@ "��      F   ,���@  ����@ %l  	` %l  	`  ����@  �      F   ,���@ ,_����@ ,dt  	` ,dt  	` ,_����@ ,_�      F   ,���@ '�,���@ ( �  	` ( �  	` '�,���@ '�,      F   ,���@ #�<���@ #��  	` #��  	` #�<���@ #�<      F   ,���@ 2�����@ 2��  	` 2��  	` 2�����@ 2��      F   ,���@ .�<���@ .��  	` .��  	` .�<���@ .�<      F   ,���@ */L���@ *3�  	` *3�  	` */L���@ */L      F   ,���@ %˴���@ %�d  	` %�d  	` %˴���@ %˴      F   ,���@ !h���@ !l�  	` !l�  	` !h���@ !h      F   ,���@ ,���@ �  	` �  	` ,���@ ,      F   ,���@ 7����@ <T  	` <T  	` 7����@ 7�      F   ,���@ 5$L���@ 5(�  	` 5(�  	` 5$L���@ 5$L      F   ,���@ 0�����@ 0�d  	` 0�d  	` 0�����@ 0��      F   ,���@ ����@ L  	` L  	` ����@ �      F   ,���@ �����@ �D  	` �D  	` �����@ ��      F   ,���@ �$���@ ��  	` ��  	` �$���@ �$      F   ,���@ s���@ w�  	` w�  	` s���@ s      F   ,���@ )���@ -�  	` -�  	` )���@ )      F   ,���@ ����@ �  	` �  	` ����@ �      F   ,���@ ����@ ��  	` ��  	` ����@ �      F   ,���@ �����@ �\  	` �\  	` �����@ ��      F   ,���@ B����@ GT  	` GT  	` B����@ B�      F   ,���@ �����@ �L  	` �L  	` �����@ ��      F   ,���@ �����@ �D  	` �D  	` �����@ ��      F   ,���@ 
d����@ 
i<  	` 
i<  	` 
d����@ 
d�      F   ,���@ ����@ 4  	` 4  	` ����@ �      F   ,���@ �����@ �D  	` �D  	` �����@ ��      F   ,���@ \4���@ `�  	` `�  	` \4���@ \4      F   ,���@ ,���@ �  	` �  	` ,���@ ,      F   ,���@ �$���@ ��  	` ��  	` �$���@ �$      F   ,���@ ~���@ ��  	` ��  	` ~���@ ~      F   ,���@ 4���@ 8�  	` 8�  	` 4���@ 4      F   ,���@ ����@ �  	` �  	` ����@ �      F   ,���@ ����@ ��  	` ��  	` ����@ �      F   ,���@ �|���@ �,  	` �,  	` �|���@ �|      F   ,���@  ����@  ��  	`  ��  	`  ����@  �      F   ,���@ 	M����@ 	RT  	` 	RT  	` 	M����@ 	M�      F   , ,�� � ,�� � ,�  � ,�  � ,�� �      F   , ,�� : ,�� >� ,�  >� ,�  : ,�� :      F   , ,�� �� ,�� �� ,�  �� ,�  �� ,�� ��      F   , ,�� � ,�� �� ,�  �� ,�  � ,�� �      F   , ,�� � ,�� 
L ,�  
L ,�  � ,�� �      F   , ,�� � ,�� �� ,�  �� ,�  � ,�� �      F   , ,�� U� ,�� ZT ,�  ZT ,�  U� ,�� U�      F   , ,�� �| ,�� �, ,�  �, ,�  �| ,�� �|      F   , ,�� � ,�� � ,�  � ,�  � ,�� �      F   , ,�� �D ,�� �� ,�  �� ,�  �D ,�� �D      F   , ,�� 
GT ,�� 
L ,�  
L ,�  
GT ,�� 
GT      F   , ,�� ;� ,�� @\ ,�  @\ ,�  ;� ,�� ;�      F   , ,�� � ,�� �� ,�  �� ,�  � ,�� �      F   , ,�� d| ,�� i, ,�  i, ,�  d| ,�� d|      F   , ,�� 	b� ,�� 	g� ,�  	g� ,�  	b� ,�� 	b�      F   , ,��  q4 ,��  u� ,�   u� ,�   q4 ,��  q4      F   , ,�� .l ,�� 3 ,�  3 ,�  .l ,�� .l      F   , ,�� � ,�� #4 ,�  #4 ,�  � ,�� �      F   , ,�� ~t ,�� �$ ,�  �$ ,�  ~t ,�� ~t      F   , ,�� �� ,�� Ǆ ,�  Ǆ ,�  �� ,�� ��      F   , ,�� �d ,�� � ,�  � ,�  �d ,�� �d      F   , ,�� r� ,�� w| ,�  w| ,�  r� ,�� r�      F   , ,�� 4 ,�� � ,�  � ,�  4 ,�� 4      F   , ,�� �L ,�� �� ,�  �� ,�  �L ,�� �L      F   , ,�� �� ,�� �d ,�  �d ,�  �� ,�� ��      F   , ,��   ,�� $� ,�  $� ,�    ,��        F   , ,�� �� ,�� �4 ,�  �4 ,�  �� ,�� ��      F   , ,�� �� ,�� �L ,�  �L ,�  �� ,�� ��      F   , ,�� W< ,�� [� ,�  [� ,�  W< ,�� W<      F   , ,�� � ,�� �T ,�  �T ,�  � ,�� �      F    ,�� $?� analog_io[10]       F    ,�� '� analog_io[11]       F    ,�� +hl analog_io[12]       F    ,�� .�� analog_io[13]       F    ,�� 2�< analog_io[14]       F    ,�� � analog_io[8]      F    ,��  �4 analog_io[9]      F    ,�� %$ io_in[10]       F    ,�� (� io_in[11]       F    ,�� ,O� io_in[12]       F    ,�� /�� io_in[13]       F    ,�� 3xT io_in[14]       F    ,�� �< io_in[8]      F    ,�� !�� io_in[9]      F    ,�� &� io_oeb[10]      F    ,�� *�� io_oeb[11]      F    ,�� .d io_oeb[12]      F    ,�� 1�� io_oeb[13]      F    ,�� 5A4 io_oeb[14]      F    ,�� 2\ io_oeb[7]       F    ,�� �� io_oeb[8]       F    ,�� #[, io_oeb[9]       F    ,�� &$ io_out[10]      F    ,�� )�� io_out[11]      F    ,�� -3� io_out[12]      F    ,�� 0�\ io_out[13]      F    ,�� 4\� io_out[14]      F    ,�� M� io_out[7]       F    ,�� �T io_out[8]       F    ,�� "v� io_out[9]       F   ���P 4 io_in[24]       F   ���P 1ܜ io_oeb[24]      F   ���P -y io_oeb[25]      F   ���P ) io_oeb[26]      F   ���P $�| io_oeb[27]      F   ���P  S� io_oeb[28]      F   ���P �� io_oeb[29]      F   ���P /�$ io_in[25]       F   ���P +H� io_in[26]       F   ���P &� io_in[27]       F   ���P "� io_in[28]       F   ���P # io_in[29]       F   ���P 0� analog_io[25]       F   ���P ,b analog_io[26]       F   ���P '�� analog_io[27]       F   ���P 2�, io_out[24]      F   ���P .�� io_out[25]      F   ���P *1� io_out[26]      F   ���P %� io_out[27]      F   ���P !jt io_out[28]      F   ���P 	� io_out[29]      F   ���P #�� analog_io[28]       F   ���P 9� analog_io[29]       F   ���P 5&� analog_io[24]       F   ���P �d io_in[33]       F   ���P �\ io_in[34]       F   ���P 	O� io_in[35]       F   ���P � io_in[36]       F   ���P �� io_in[37]       F   ���P � analog_io[30]       F   ���P �| io_in[30]       F   ���P ut io_in[31]       F   ���P +l io_in[32]       F   ���P � io_oeb[30]      F   ���P D� io_oeb[31]      F   ���P �� io_oeb[32]      F   ���P �� io_oeb[33]      F   ���P 
f� io_oeb[34]      F   ���P �� io_out[30]      F   ���P ^� io_out[31]      F   ���P � io_out[32]      F   ���P �| io_out[33]      F   ���P �t io_out[34]      F   ���P 6l io_out[35]      F   ���P �d io_out[36]      F   ���P �\ io_out[37]      F   ���P � io_oeb[35]      F   ���P �� io_oeb[36]      F   ���P  �t io_oeb[37]      F    ,�� �d io_in[1]      F    ,�� <l io_out[0]       F    ,�� �D io_oeb[1]       F    ,�� �d analog_io[7]      F    ,�� � analog_io[1]      F    ,�� �\ analog_io[2]      F    ,�� W� io_in[0]      F    ,�� �� io_out[1]       F    ,�� 4 io_in[3]      F    ,�� �� io_in[4]      F    ,�� 
I� io_oeb[2]       F    ,�� > io_in[5]      F    ,�� �l io_in[6]      F    ,�� f� io_in[7]      F    ,�� 	e< io_out[2]       F    ,��  s� analog_io[0]      F    ,�� 0� analog_io[3]      F    ,��  � io_oeb[0]       F    ,�� �� io_in[2]      F    ,�� �, analog_io[4]      F    ,�� � io_oeb[3]       F    ,�� u$ io_oeb[4]       F    ,�� 	� io_oeb[5]       F    ,�� �� io_out[3]       F    ,�� � io_out[4]       F    ,�� "t io_out[5]       F    ,�� �� io_out[6]       F    ,�� �� io_oeb[6]       F    ,�� Y� analog_io[5]      F    ,�� �� analog_io[6]      E   , EJ���@ EJ  	` Gz  	` Gz���@ EJ���@      E   , &�� 5�� &�� 5�� &�� 5�� &�� 5�� &�� 5��      E   , "� 5�� "� 5�� "
 5�� "
 5�� "� 5��      E   , B 5�� B 5�� r 5�� r 5�� B 5��      E   , !v 5�� !v 5�� #� 5�� #� 5�� !v 5��      E   , *�2 5�� *�2 5�� *�b 5�� *�b 5�� *�2 5��      E   , %�f 5�� %�f 5�� %�� 5�� %�� 5�� %�f 5��      E   ,  �� 5��  �� 5��  �� 5��  �� 5��  �� 5��      E   , � 5�� � 5�� �2 5�� �2 5�� � 5��      E   , �6 5�� �6 5�� �f 5�� �f 5�� �6 5��      E   , (7� 5�� (7� 5�� (: 5�� (: 5�� (7� 5��      E   , #E 5�� #E 5�� #GJ 5�� #GJ 5�� #E 5��      E   , RN 5�� RN 5�� T~ 5�� T~ 5�� RN 5��      E   , ]� 5�� ]� 5�� _� 5�� _� 5�� ]� 5��      E   , )u� 5�� )u� 5�� )x" 5�� )x" 5�� )u� 5��      E   , $�Z 5�� $�Z 5�� $�� 5�� $�� 5�� $�Z 5��      E   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      E   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      E   , +�r 5�� +�r 5�� +� 5�� +� 5�� +�r 5��      E   , 	GF 5�� 	GF 5�� 	Iv 5�� 	Iv 5�� 	GF 5��      E   , Tz 5�� Tz 5�� V� 5�� V� 5�� Tz 5��      E   , .� 5�� .� 5�� 0� 5�� 0� 5�� .� 5��      E   , j� 5�� j� 5�� m 5�� m 5�� j� 5��      E   , x 5�� x 5�� zN 5�� zN 5�� x 5��      E   , 
�� 5�� 
�� 5�� 
�� 5�� 
�� 5�� 
�� 5��      E   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      E   ,  �� 5��  �� 5��  � 5��  � 5��  �� 5��      E   , � 5�� � 5�� �� 5�� �� 5�� � 5��      E   , �� 5�� �� 5��   5��   5�� �� 5��      E   ,  5��  5�� 6 5�� 6 5��  5��      E   , n 5�� n 5�� � 5�� � 5�� n 5��      E   , �* 5�� �* 5�� �Z 5�� �Z 5�� �* 5��      E   , �^ 5�� �^ 5�� �� 5�� �� 5�� �^ 5��      E   , �� 5�� �� 5�� �� 5�� �� 5�� �� 5��      E   , �� 5�� �� 5�� �* 5�� �* 5�� �� 5��      E   , �. 5�� �. 5�� �^ 5�� �^ 5�� �. 5��      E   , : 5�� : 5�� <B 5�� <B 5�� : 5��      E   ,  
����@  
�  	`  �  	`  ����@  
����@      E   ,   &���@   &  	`  "V  	`  "V���@   &���@      E   ,  7����@  7�  	`  9�  	`  9����@  7����@      E   ,  �����@  ��  	`  �"  	`  �"���@  �����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �
  	` �
���@ �����@      E   , 5����@ 5�  	` 8  	` 8���@ 5����@      E   , |���@ |  	` ~2  	` ~2���@ |���@      E   , ����@ �  	` �F  	` �F���@ ����@      E   , *���@ *  	` 
Z  	` 
Z���@ *���@      E   , Lr���@ Lr  	` N�  	` N����@ Lr���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   ,  �b���@  �b  	`  ��  	`  �����@  �b���@      E   , O����@ O�  	` R  	` R���@ O����@      E   , �v���@ �v  	` ��  	` �����@ �v���@      E   , ����@ �  	`   	` ���@ ����@      E   , N����@ N�  	` Q*  	` Q*���@ N����@      E   , ����@ �  	` �>  	` �>���@ ����@      E   , �V���@ �V  	` ۆ  	` ۆ���@ �V���@      E   , j���@ j  	` !�  	` !����@ j���@      E   , e~���@ e~  	` g�  	` g����@ e~���@      E   ,  N����@  N�  	`  Q  	`  Q���@  N����@      E   ,  �N���@  �N  	`  �~  	`  �~���@  �N���@      E   , �����@ ��  	` �  	` ����@ �����@      E   , 6���@ 6  	` 	f  	` 	f���@ 6���@      E   , MJ���@ MJ  	` Oz  	` Oz���@ MJ���@      E   , �^���@ �^  	` ��  	` �����@ �^���@      E   , �r���@ �r  	` ۢ  	` ۢ���@ �r���@      E   , ����@ �  	` !�  	` !����@ ����@      E   , c����@ c�  	` e�  	` e����@ c����@      E   , 	����@ 	�  	` �  	` ����@ 	����@      E   , eb���@ eb  	` g�  	` g����@ eb���@      E   , �����@ ��  	` �  	` ����@ �����@      E   ,  B���@  B  	` "r  	` "r���@  B���@      E   , fV���@ fV  	` h�  	` h����@ fV���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` ��  	` �����@ ����@      E   , 6����@ 6�  	` 8�  	` 8����@ 6����@      E   , |����@ |�  	` 
  	` 
���@ |����@      E   ,  ê���@  ê  	`  ��  	`  �����@  ê���@      E   , �J���@ �J  	` �z  	` �z���@ �J���@      E   , ����@ �  	`  �  	`  ����@ ����@      E   , d����@ d�  	` f�  	` f����@ d����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , 5���@ 5  	` 7F  	` 7F���@ 5���@      E   , {*���@ {*  	` }Z  	` }Z���@ {*���@      E   , !���@ !  	` #J  	` #J���@ !���@      E   , |����@ |�  	` ~�  	` ~����@ |����@      E   , �.���@ �.  	` �^  	` �^���@ �.���@      E   , 7����@ 7�  	` 9�  	` 9����@ 7����@      E   , }����@ }�  	` �  	` ����@ }����@      E   , �����@ ��  	` �*  	` �*���@ �����@      E   , ���@   	` 
>  	` 
>���@ ���@      E   , N"���@ N"  	` PR  	` PR���@ N"���@      E   , �6���@ �6  	` �f  	` �f���@ �6���@      E   ,  ����@  �  	`  �6  	`  �6���@  ����@      E   , 8v���@ 8v  	` :�  	` :����@ 8v���@      E   , ����@ �  	` �J  	` �J���@ ����@      E   , ����@ �  	` �  	` ����@ ����@      E   ,  f:���@  f:  	`  hj  	`  hj���@  f:���@      E   ,  }����@  }�  	`  �  	`  ����@  }����@      E   , �����@ ��  	` �&  	` �&���@ �����@      E   , 6
���@ 6
  	` 8:  	` 8:���@ 6
���@      E   , ����@ �  	`  �  	`  ����@ ����@      E   , zR���@ zR  	` |�  	` |����@ zR���@      E   , �f���@ �f  	`   	` ���@ �f���@      E   , z���@ z  	` �  	` ����@ z���@      E   , L����@ L�  	` N�  	` N����@ L����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , ����@ �  	` .  	` .���@ ����@      E   , c���@ c  	` eB  	` eB���@ c���@      E   , �&���@ �&  	` �V  	` �V���@ �&���@      E   , �:���@ �:  	` �j  	` �j���@ �:���@      E   , 	����@ 	�  	` 	�6  	` 	�6���@ 	����@      E   , 	3����@ 	3�  	` 	5�  	` 	5����@ 	3����@      E   , 	y����@ 	y�  	` 	{�  	` 	{����@ 	y����@      E   , d����@ d�  	` f�  	` f����@ d����@      E   , �
���@ �
  	` �:  	` �:���@ �
���@      E   , ����@ �  	` �N  	` �N���@ ����@      E   , 52���@ 52  	` 7b  	` 7b���@ 52���@      E   , {F���@ {F  	` }v  	` }v���@ {F���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �  	` ����@ ����@      E   , K����@ K�  	` M�  	` M����@ K����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , 
���@ 
  	` 
J  	` 
J���@ 
���@      E   , 	&���@ 	&  	` 	V  	` 	V���@ 	&���@      E   , 	b:���@ 	b:  	` 	dj  	` 	dj���@ 	b:���@      E   , 
ab���@ 
ab  	` 
c�  	` 
c����@ 
ab���@      E   , 
�v���@ 
�v  	` 
��  	` 
�����@ 
�v���@      E   , �>���@ �>  	` �n  	` �n���@ �>���@      E   , R���@ R  	` 	�  	` 	����@ R���@      E   , Mf���@ Mf  	` O�  	` O����@ Mf���@      E   , 
����@ 
�  	` 
�  	` 
����@ 
����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	`    	`  ���@ ����@      E   , c����@ c�  	` f  	` f���@ c����@      E   , �����@ ��  	` �.  	` �.���@ �����@      E   , �F���@ �F  	` �v  	` �v���@ �F���@      E   , 4Z���@ 4Z  	` 6�  	` 6����@ 4Z���@      E   , zn���@ zn  	` |�  	` |����@ zn���@      E   , �����@ ��  	` ²  	` ²���@ �����@      E   , 	����@ 	�  	` 	�  	` 	����@ 	����@      E   , 	�b���@ 	�b  	` 	�  	` 	����@ 	�b���@      E   , 	J����@ 	J�  	` 	M  	` 	M���@ 	J����@      E   , 	�����@ 	��  	` 	�"  	` 	�"���@ 	�����@      E   , 
4v���@ 
4v  	` 
6�  	` 
6����@ 
4v���@      E   , 
x����@ 
x�  	` 
z�  	` 
z����@ 
x����@      E   , 
�����@ 
��  	` 
�  	` 
����@ 
�����@      E   , ����@ �  	`   	` ���@ ����@      E   , 	�����@ 	��  	` 	��  	` 	�����@ 	�����@      E   , 
����@ 
�  	` 
�  	` 
����@ 
����@      E   , 
J���@ 
J  	` 
L6  	` 
L6���@ 
J���@      E   , 
����@ 
�  	` 
�J  	` 
�J���@ 
����@      E   , 	�N���@ 	�N  	` 	�~  	` 	�~���@ 	�N���@      E   , 
�.���@ 
�.  	` 
�^  	` 
�^���@ 
�.���@      E   , B���@ B  	` r  	` r���@ B���@      E   , ؚ���@ ؚ  	` ��  	` �����@ ؚ���@      E   , �����@ ��  	` �  	` ����@ �����@      E   , 12���@ 12  	` 3b  	` 3b���@ 12���@      E   , wF���@ wF  	` yv  	` yv���@ wF���@      E   , 3����@ 3�  	` 5�  	` 5����@ 3����@      E   , y����@ y�  	` {�  	` {����@ y����@      E   , �����@ ��  	` �*  	` �*���@ �����@      E   , ���@   	` >  	` >���@ ���@      E   , J"���@ J"  	` LR  	` LR���@ J"���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �
  	` �
���@ �����@      E   , 1����@ 1�  	` 4  	` 4���@ 1����@      E   , x���@ x  	` z2  	` z2���@ x���@      E   , J����@ J�  	` M*  	` M*���@ J����@      E   , �B���@ �B  	` �r  	` �r���@ �B���@      E   , �V���@ �V  	` ׆  	` ׆���@ �V���@      E   , j���@ j  	` �  	` ����@ j���@      E   , ����@ �  	` �F  	` �F���@ ����@      E   , x����@ x�  	` {
  	` {
���@ x����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , 6���@ 6  	` f  	` f���@ 6���@      E   , IJ���@ IJ  	` Kz  	` Kz���@ IJ���@      E   , �^���@ �^  	` ��  	` �����@ �^���@      E   , �r���@ �r  	` ע  	` ע���@ �r���@      E   , ����@ �  	` �  	` ����@ ����@      E   , _����@ _�  	` a�  	` a����@ _����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �����@ ��  	` �&  	` �&���@ �����@      E   , *���@ *  	` Z  	` Z���@ *���@      E   , 2
���@ 2
  	` 4:  	` 4:���@ 2
���@      E   , vR���@ vR  	` x�  	` x����@ vR���@      E   , �f���@ �f  	` ��  	` �����@ �f���@      E   , z���@ z  	` �  	` ����@ z���@      E   , H����@ H�  	` J�  	` J����@ H����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , Hr���@ Hr  	` J�  	` J����@ Hr���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , Ԛ���@ Ԛ  	` ��  	` �����@ Ԛ���@      E   , a~���@ a~  	` c�  	` c����@ a~���@      E   , ����@ �  	` �  	` ����@ ����@      E   , bV���@ bV  	` d�  	` d����@ bV���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` ��  	` �����@ ����@      E   , 2����@ 2�  	` 4�  	` 4����@ 2����@      E   , ^����@ ^�  	` a&  	` a&���@ ^����@      E   , �6���@ �6  	` �f  	` �f���@ �6���@      E   , �~���@ �~  	` ֮  	` ֮���@ �~���@      E   , ����@ �  	` �  	` ����@ ����@      E   , `����@ `�  	` b�  	` b����@ `����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , 1���@ 1  	` 3F  	` 3F���@ 1���@      E   , w*���@ w*  	` yZ  	` yZ���@ w*���@      E   , �>���@ �>  	` �n  	` �n���@ �>���@      E   , R���@ R  	` �  	` ����@ R���@      E   , �
���@ �
  	` �:  	` �:���@ �
���@      E   , If���@ If  	` K�  	` K����@ If���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	`   	` ���@ ����@      E   , _����@ _�  	` b  	` b���@ _����@      E   , �2���@ �2  	` �b  	` �b���@ �2���@      E   , ����@ �  	` �N  	` �N���@ ����@      E   , �~���@ �~  	` Ү  	` Ү���@ �~���@      E   , �B���@ �B  	` �r  	` �r���@ �B���@      E   , �����@ ��  	` �  	` ����@ �����@      E   , ����@ �  	` .  	` .���@ ����@      E   , _���@ _  	` aB  	` aB���@ _���@      E   , �&���@ �&  	` �V  	` �V���@ �&���@      E   , �V���@ �V  	` ӆ  	` ӆ���@ �V���@      E   , �n���@ �n  	` �  	` ����@ �n���@      E   , /����@ /�  	` 1�  	` 1����@ /����@      E   , u����@ u�  	` w�  	` w����@ u����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �  	` ����@ ����@      E   , F���@ F  	` H6  	` H6���@ F���@      E   , ����@ �  	` �J  	` �J���@ ����@      E   , �.���@ �.  	` �^  	` �^���@ �.���@      E   , B���@ B  	` r  	` r���@ B���@      E   , ^V���@ ^V  	` `�  	` `����@ ^V���@      E   , j���@ j  	` �  	` ����@ j���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` ��  	` �����@ ����@      E   , .����@ .�  	` 0�  	` 0����@ .����@      E   , t����@ t�  	` w
  	` w
���@ t����@      E   , �"���@ �"  	` �R  	` �R���@ �"���@      E   , �6���@ �6  	` f  	` f���@ �6���@      E   , ]~���@ ]~  	` _�  	` _����@ ]~���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �
  	` �
���@ �����@      E   , -����@ -�  	` 0  	` 0���@ -����@      E   , ����@ �  	` �  	` ����@ ����@      E   , /����@ /�  	` 1�  	` 1����@ /����@      E   , s����@ s�  	` v  	` v���@ s����@      E   , ����@ �  	` �  	` ����@ ����@      E   , �����@ ��  	` �*  	` �*���@ �����@      E   ,  ���@    	` >  	` >���@  ���@      E   , F"���@ F"  	` HR  	` HR���@ F"���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �  	` ����@ ����@      E   , G����@ G�  	` I�  	` I����@ G����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �6���@ �6  	` �f  	` �f���@ �6���@      E   , �����@ ��  	` �  	` ����@ �����@      E   , &���@ &  	` V  	` V���@ &���@      E   , ^:���@ ^:  	` `j  	` `j���@ ^:���@      E   , �N���@ �N  	` �~  	` �~���@ �N���@      E   , �b���@ �b  	` �  	` ����@ �b���@      E   , .����@ .�  	` 0�  	` 0����@ .����@      E   , t����@ t�  	` v�  	` v����@ t����@      E   , �����@ ��  	` �  	` ����@ �����@      E   ,  ����@  �  	`   	` ���@  ����@      E   , �F���@ �F  	` �v  	` �v���@ �F���@      E   , 0Z���@ 0Z  	` 2�  	` 2����@ 0Z���@      E   , vn���@ vn  	` x�  	` x����@ vn���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , F����@ F�  	` I*  	` I*���@ F����@      E   ,  ����@  �  	` �  	` ����@  ����@      E   , F����@ F�  	` I  	` I���@ F����@      E   , �����@ ��  	` �"  	` �"���@ �����@      E   , ����@ �  	` �6  	` �6���@ ����@      E   , ���@   	` J  	` J���@ ���@      E   , ]b���@ ]b  	` _�  	` _����@ ]b���@      E   , �v���@ �v  	` ��  	` �����@ �v���@      E   , \����@ \�  	` ^�  	` ^����@ \����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , -���@ -  	` /F  	` /F���@ -���@      E   , s*���@ s*  	` uZ  	` uZ���@ s*���@      E   , �>���@ �>  	` �n  	` �n���@ �>���@      E   , �R���@ �R  	` �  	` ����@ �R���@      E   , C����@ C�  	` E�  	` E����@ C����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	`   	` ���@ ����@      E   , [����@ [�  	` ^  	` ^���@ [����@      E   , �2���@ �2  	` �b  	` �b���@ �2���@      E   , �F���@ �F  	` �v  	` �v���@ �F���@      E   , ,Z���@ ,Z  	` .�  	` .����@ ,Z���@      E   , rn���@ rn  	` t�  	` t����@ rn���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , B����@ B�  	` E  	` E���@ B����@      E   , �����@ ��  	` �"  	` �"���@ �����@      E   , ����@ �  	` �6  	` �6���@ ����@      E   , t���@ t  	` v2  	` v2���@ t���@      E   , ����@ �  	` �F  	` �F���@ ����@      E   , �^���@ �^  	`  �  	`  ����@ �^���@      E   , Dr���@ Dr  	` F�  	` F����@ Dr���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , К���@ К  	` ��  	` �����@ К���@      E   , ����@ �  	` �  	` ����@ ����@      E   , Z����@ Z�  	` ]&  	` ]&���@ Z����@      E   , �
���@ �
  	` �:  	` �:���@ �
���@      E   , ����@ �  	` �N  	` �N���@ ����@      E   , -2���@ -2  	` /b  	` /b���@ -2���@      E   , sF���@ sF  	` uv  	` uv���@ sF���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , C����@ C�  	` E�  	` E����@ C����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �B  	` �B���@ ����@      E   , �^���@ �^  	` ��  	` �����@ �^���@      E   , �r���@ �r  	` Ӣ  	` Ӣ���@ �r���@      E   , ����@ �  	` �  	` ����@ ����@      E   , &���@ &  	` V  	` V���@ &���@      E   , [����@ [�  	` ]�  	` ]����@ [����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �����@ ��  	` �&  	` �&���@ �����@      E   , .
���@ .
  	` 0:  	` 0:���@ .
���@      E   , rR���@ rR  	` t�  	` t����@ rR���@      E   , �f���@ �f  	` ��  	` �����@ �f���@      E   , �z���@ �z  	`  �  	`  ����@ �z���@      E   , D����@ D�  	` F�  	` F����@ D����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , Z:���@ Z:  	` \j  	` \j���@ Z:���@      E   , ����@ �  	` .  	` .���@ ����@      E   , [���@ [  	` ]B  	` ]B���@ [���@      E   , �&���@ �&  	` �V  	` �V���@ �&���@      E   , �n���@ �n  	` �  	` ����@ �n���@      E   , +����@ +�  	` -�  	` -����@ +����@      E   , q����@ q�  	` s�  	` s����@ q����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �N���@ �N  	` �~  	` �~���@ �N���@      E   , B����@ B�  	` E*  	` E*���@ B����@      E   , �B���@ �B  	` �r  	` �r���@ �B���@      E   , �V���@ �V  	` φ  	` φ���@ �V���@      E   , j���@ j  	` �  	` ����@ j���@      E   , Y~���@ Y~  	` [�  	` [����@ Y~���@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , �����@ ��  	` �
  	` �
���@ �����@      E   , )����@ )�  	` ,  	` ,���@ )����@      E   , p���@ p  	` r2  	` r2���@ p���@      E   , ����@ �  	` �F  	` �F���@ ����@      E   , �^���@ �^  	` ��  	` �����@ �^���@      E   ,  @r���@  @r  	`  B�  	`  B����@  @r���@      E   ,  �����@  ��  	`  ��  	`  �����@  �����@      E   ,  ̚���@  ̚  	`  ��  	`  �����@  ̚���@      E   , !����@ !�  	` !�  	` !����@ !����@      E   , !V����@ !V�  	` !Y&  	` !Y&���@ !V����@      E   , p����@ p�  	` r�  	` r����@ p����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , N���@ N  	` ~  	` ~���@ N���@      E   , Yb���@ Yb  	` [�  	` [����@ Yb���@      E   , �v���@ �v  	` ��  	` �����@ �v���@      E   , ����@ �  	` �  	` ����@ ����@      E   , +����@ +�  	` -�  	` -����@ +����@      E   , o����@ o�  	` r  	` r���@ o����@      E   , �����@ ��  	` �*  	` �*���@ �����@      E   , ����@ �  	` �>  	` �>���@ ����@      E   , B"���@ B"  	` DR  	` DR���@ B"���@      E   , �6���@ �6  	` �f  	` �f���@ �6���@      E   , �~���@ �~  	` ή  	` ή���@ �~���@      E   , ����@ �  	` �  	` ����@ ����@      E   , X����@ X�  	` Z�  	` Z����@ X����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` �2  	` �2���@ ����@      E   ,  )���@  )  	`  +F  	`  +F���@  )���@      E   ,  o*���@  o*  	`  qZ  	`  qZ���@  o*���@      E   ,  �>���@  �>  	`  �n  	`  �n���@  �>���@      E   ,  �R���@  �R  	`  ��  	`  �����@  �R���@      E   , !?����@ !?�  	` !A�  	` !A����@ !?����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , B���@ B  	` D6  	` D6���@ B���@      E   , ����@ �  	` �J  	` �J���@ ����@      E   , �����@ ��  	` �  	` ����@ �����@      E   , �.���@ �.  	` �^  	` �^���@ �.���@      E   , B���@ B  	` r  	` r���@ B���@      E   , X����@ X�  	` Z�  	` Z����@ X����@      E   , �����@ ��  	` ��  	` �����@ �����@      E   , ����@ �  	` ��  	` �����@ ����@      E   , *����@ *�  	` ,�  	` ,����@ *����@      E   , p����@ p�  	` s
  	` s
���@ p����@      E   , �"���@ �"  	` �R  	` �R���@ �"���@      E   , �6���@ �6  	` �f  	` �f���@ �6���@      E   , AJ���@ AJ  	` Cz  	` Cz���@ AJ���@      E   , �b���@ �b  	` �  	` ����@ �b���@      E   , �^���@ �^  	` ��  	` �����@ �^���@      E   , �r���@ �r  	` Ϣ  	` Ϣ���@ �r���@      E   ,  ����@  �  	`  �  	`  ����@  ����@      E   ,  W����@  W�  	`  Y�  	`  Y����@  W����@      E   ,  �����@  ��  	`  �  	`  ����@  �����@      E   ,  �����@  ��  	`  �&  	`  �&���@  �����@      E   , !(>���@ !(>  	` !*n  	` !*n���@ !(>���@      E   , *����@ *�  	` ,�  	` ,����@ *����@      E   , !����@ !�  	` !�N  	` !�N���@ !����@      E   , !�����@ !��  	` !��  	` !�����@ !�����@      E   , !�����@ !��  	` !��  	` !�����@ !�����@      E   , "����@ "�  	` "  	` "���@ "����@      E   , "W����@ "W�  	` "Z  	` "Z���@ "W����@      E   , "�2���@ "�2  	` "�b  	` "�b���@ "�2���@      E   , "�F���@ "�F  	` "�v  	` "�v���@ "�F���@      E   , #(Z���@ #(Z  	` #*�  	` #*����@ #(Z���@      E   , #nn���@ #nn  	` #p�  	` #p����@ #nn���@      E   , #�����@ #��  	` #��  	` #�����@ #�����@      E   , #�����@ #��  	` #��  	` #�����@ #�����@      E   , $>����@ $>�  	` $A  	` $A���@ $>����@      E   , $�����@ $��  	` $�"  	` $�"���@ $�����@      E   , $����@ $�  	` $�6  	` $�6���@ $����@      E   , %&����@ %&�  	` %(�  	` %(����@ %&����@      E   , %l����@ %l�  	` %n�  	` %n����@ %l����@      E   , %�����@ %��  	` %�  	` %����@ %�����@      E   , %�����@ %��  	` %�  	` %����@ %�����@      E   , &=.���@ &=.  	` &?^  	` &?^���@ &=.���@      E   , &�B���@ &�B  	` &�r  	` &�r���@ &�B���@      E   , &�V���@ &�V  	` &ˆ  	` &ˆ���@ &�V���@      E   , $�b���@ $�b  	` $�  	` $����@ $�b���@      E   , ")2���@ ")2  	` "+b  	` "+b���@ ")2���@      E   , "mz���@ "mz  	` "o�  	` "o����@ "mz���@      E   , "�����@ "��  	` "��  	` "�����@ "�����@      E   , "�����@ "��  	` "��  	` "�����@ "�����@      E   , #?����@ #?�  	` #A�  	` #A����@ #?����@      E   , #�����@ #��  	` #��  	` #�����@ #�����@      E   , #����@ #�  	` #�B  	` #�B���@ #����@      E   , $&���@ $&  	` $V  	` $V���@ $&���@      E   , $V:���@ $V:  	` $Xj  	` $Xj���@ $V:���@      E   , $�N���@ $�N  	` $�~  	` $�~���@ $�N���@      E   , $�����@ $��  	` $�"  	` $�"���@ $�����@      E   , %>���@ %>  	` %@6  	` %@6���@ %>���@      E   , %����@ %�  	` %�J  	` %�J���@ %����@      E   , %�.���@ %�.  	` %�^  	` %�^���@ %�.���@      E   , &B���@ &B  	` &r  	` &r���@ &B���@      E   , "�����@ "��  	` "�  	` "����@ "�����@      E   , &T����@ &T�  	` &V�  	` &V����@ &T����@      E   , #����@ #�  	` #.  	` #.���@ #����@      E   , &�����@ &��  	` &��  	` &�����@ &�����@      E   , #W���@ #W  	` #YB  	` #YB���@ #W���@      E   , #�&���@ #�&  	` #�V  	` #�V���@ #�&���@      E   , &����@ &�  	` &��  	` &�����@ &����@      E   , #�n���@ #�n  	` #�  	` #����@ #�n���@      E   , $'����@ $'�  	` $)�  	` $)����@ $'����@      E   , $m����@ $m�  	` $o�  	` $o����@ $m����@      E   , $�����@ $��  	` $��  	` $�����@ $�����@      E   , "�����@ "��  	` "�  	` "����@ "�����@      E   , %N���@ %N  	` %~  	` %~���@ %N���@      E   , %Ub���@ %Ub  	` %W�  	` %W����@ %Ub���@      E   , %�v���@ %�v  	` %��  	` %�����@ %�v���@      E   , %����@ %�  	` %�  	` %����@ %����@      E   , &'����@ &'�  	` &)�  	` &)����@ &'����@      E   , &k����@ &k�  	` &n  	` &n���@ &k����@      E   , &�����@ &��  	` &�*  	` &�*���@ &�����@      E   , !nR���@ !nR  	` !p�  	` !p����@ !nR���@      E   , !�f���@ !�f  	` !��  	` !�����@ !�f���@      E   , !�z���@ !�z  	` !��  	` !�����@ !�z���@      E   , !�
���@ !�
  	` !�:  	` !�:���@ !�
���@      E   , "@����@ "@�  	` "B�  	` "B����@ "@����@      E   , *$>���@ *$>  	` *&n  	` *&n���@ *$>���@      E   , *����@ *�  	` *  	` *���@ *����@      E   , *jR���@ *jR  	` *l�  	` *l����@ *jR���@      E   , *�f���@ *�f  	` *��  	` *�����@ *�f���@      E   , *�z���@ *�z  	` *��  	` *�����@ *�z���@      E   , +<����@ +<�  	` +>�  	` +>����@ +<����@      E   , )<r���@ )<r  	` )>�  	` )>����@ )<r���@      E   , )�����@ )��  	` )��  	` )�����@ )�����@      E   , (%����@ (%�  	` ((  	` ((���@ (%����@      E   , +�����@ +��  	` +�  	` +����@ +�����@      E   , +�����@ +��  	` +�  	` +����@ +�����@      E   , ,����@ ,�  	` ,.  	` ,.���@ ,����@      E   , ,S���@ ,S  	` ,UB  	` ,UB���@ ,S���@      E   , 'l����@ 'l�  	` 'o
  	` 'o
���@ 'l����@      E   , '>"���@ '>"  	` '@R  	` '@R���@ '>"���@      E   , '�j���@ '�j  	` '��  	` '�����@ '�j���@      E   , *R����@ *R�  	` *U&  	` *U&���@ *R����@      E   , '�~���@ '�~  	` 'ʮ  	` 'ʮ���@ '�~���@      E   , *�
���@ *�
  	` *�:  	` *�:���@ *�
���@      E   , (����@ (�  	` (�  	` (����@ (����@      E   , (T����@ (T�  	` (V�  	` (V����@ (T����@      E   , (�����@ (��  	` (��  	` (�����@ (�����@      E   , (����@ (�  	` (�2  	` (�2���@ (����@      E   , )%���@ )%  	` )'F  	` )'F���@ )%���@      E   , )k*���@ )k*  	` )mZ  	` )mZ���@ )k*���@      E   , )�>���@ )�>  	` )�n  	` )�n���@ )�>���@      E   , )�R���@ )�R  	` )��  	` )�����@ )�R���@      E   , *;����@ *;�  	` *=�  	` *=����@ *;����@      E   , *����@ *�  	` *�N  	` *�N���@ *����@      E   , +%2���@ +%2  	` +'b  	` +'b���@ +%2���@      E   , *�����@ *��  	` *��  	` *�����@ *�����@      E   , *�����@ *��  	` *��  	` *�����@ *�����@      E   , +����@ +�  	` +  	` +���@ +����@      E   , +R���@ +R  	` +TN  	` +TN���@ +R���@      E   , +�2���@ +�2  	` +�b  	` +�b���@ +�2���@      E   , +�F���@ +�F  	` +�v  	` +�v���@ +�F���@      E   , ,$Z���@ ,$Z  	` ,&�  	` ,&����@ ,$Z���@      E   , ,jn���@ ,jn  	` ,l�  	` ,l����@ ,jn���@      E   , +iz���@ +iz  	` +k�  	` +k����@ +iz���@      E   , +�����@ +��  	` +��  	` +�����@ +�����@      E   , +�����@ +��  	` +��  	` +�����@ +�����@      E   , ,;����@ ,;�  	` ,=�  	` ,=����@ ,;����@      E   , )Ț���@ )Ț  	` )��  	` )�����@ )Ț���@      E   , ,�����@ ,��  	` ,��  	` ,�����@ ,�����@      E   , '�"���@ '�"  	` '�R  	` '�R���@ '�"���@      E   , '�6���@ '�6  	` '�f  	` '�f���@ '�6���@      E   , (l���@ (l  	` (n2  	` (n2���@ (l���@      E   , (����@ (�  	` (�F  	` (�F���@ (����@      E   , (=J���@ (=J  	` (?z  	` (?z���@ (=J���@      E   , (�^���@ (�^  	` (��  	` (�����@ (�^���@      E   , 'j���@ 'j  	` '�  	` '����@ 'j���@      E   , '&����@ '&�  	` '(�  	` '(����@ '&����@      E   , 'U~���@ 'U~  	` 'W�  	` 'W����@ 'U~���@      E   , (Ǧ���@ (Ǧ  	` (��  	` (�����@ (Ǧ���@      E   , '�����@ '��  	` '��  	` '�����@ '�����@      E   , (�^���@ (�^  	` (��  	` (�����@ (�^���@      E   , &����@ &�  	` &�>  	` &�>���@ &����@      E   , )����@ )�  	` )�  	` )����@ )����@      E   , )S����@ )S�  	` )U�  	` )U����@ )S����@      E   , '�����@ '��  	` '�
  	` '�
���@ '�����@      E   , )�����@ )��  	` )�  	` )����@ )�����@      E   , )�����@ )��  	` )�&  	` )�&���@ )�����@      E    +� 5�� analog_io[15]       E    &�� 5�� analog_io[16]       E    "	� 5�� analog_io[17]       E    Z 5�� analog_io[18]       E    "� 5�� analog_io[19]       E    *�J 5�� io_in[15]       E    %�~ 5�� io_in[16]       E     �� 5�� io_in[17]       E    � 5�� io_in[18]       E    �N 5�� io_in[19]       E    (8� 5�� io_oeb[15]      E    #F2 5�� io_oeb[16]      E    Sf 5�� io_oeb[17]      E    ^� 5�� io_oeb[18]      E    )w
 5�� io_out[15]      E    $�r 5�� io_out[16]      E    �� 5�� io_out[17]      E    �� 5�� io_out[18]      E    ;* 5�� analog_io[21]       E    	H^ 5�� analog_io[22]       E    U� 5�� analog_io[23]       E    /� 5�� analog_io[20]       E    l 5�� io_oeb[19]      E    y6 5�� io_oeb[20]      E    
�� 5�� io_oeb[21]      E    �� 5�� io_oeb[22]      E     � 5�� io_oeb[23]      E    � 5�� io_in[20]       E    �� 5�� io_in[21]       E     5�� io_in[22]       E    � 5�� io_in[23]       E    �B 5�� io_out[19]      E    �v 5�� io_out[20]      E    ª 5�� io_out[21]      E    � 5�� io_out[22]      E    �F 5�� io_out[23]      E     ����P wb_clk_i      E     !>���P wb_rst_i      E     8����P wbs_ack_o       E     �
���P wbs_adr_i[0]      E    �����P wbs_adr_i[10]       E    �����P wbs_adr_i[11]       E    7���P wbs_adr_i[12]       E    }���P wbs_adr_i[13]       E    �.���P wbs_adr_i[14]       E    	B���P wbs_adr_i[15]       E    M����P wbs_adr_i[16]       E    �����P wbs_adr_i[17]       E     �z���P wbs_adr_i[1]      E    P����P wbs_adr_i[2]      E    �����P wbs_adr_i[3]      E    	����P wbs_adr_i[4]      E    P���P wbs_adr_i[5]      E    �&���P wbs_adr_i[6]      E    �n���P wbs_adr_i[7]      E     ����P wbs_adr_i[8]      E    f����P wbs_adr_i[9]      E     O����P wbs_cyc_i       E     �f���P wbs_dat_i[0]      E    ����P wbs_dat_i[10]       E    N���P wbs_dat_i[11]       E    Nb���P wbs_dat_i[12]       E    �v���P wbs_dat_i[13]       E    ڊ���P wbs_dat_i[14]       E     ����P wbs_dat_i[15]       E    d����P wbs_dat_i[16]       E    
����P wbs_dat_i[1]      E    fz���P wbs_dat_i[2]      E    �����P wbs_dat_i[3]      E    !Z���P wbs_dat_i[4]      E    gn���P wbs_dat_i[5]      E    �����P wbs_dat_i[6]      E    �����P wbs_dat_i[7]      E    7����P wbs_dat_i[8]      E    }����P wbs_dat_i[9]      E     �����P wbs_dat_o[0]      E    �b���P wbs_dat_o[10]       E    ����P wbs_dat_o[11]       E    e����P wbs_dat_o[12]       E    �����P wbs_dat_o[13]       E    �����P wbs_dat_o[14]       E    6.���P wbs_dat_o[15]       E    |B���P wbs_dat_o[16]       E    "2���P wbs_dat_o[1]      E    }����P wbs_dat_o[2]      E    �F���P wbs_dat_o[3]      E    8����P wbs_dat_o[4]      E    ~����P wbs_dat_o[5]      E    ����P wbs_dat_o[6]      E    	&���P wbs_dat_o[7]      E    O:���P wbs_dat_o[8]      E    �N���P wbs_dat_o[9]      E     ����P wbs_sel_i[0]      E    9����P wbs_sel_i[1]      E    �2���P wbs_sel_i[2]      E    ����P wbs_sel_i[3]      E     gR���P wbs_stb_i       E     ~����P wbs_we_i      E    ����P wbs_dat_i[18]       E    7"���P wbs_dat_i[19]       E    ����P wbs_adr_i[19]       E    {j���P wbs_dat_i[20]       E    �~���P wbs_dat_i[21]       E    ����P wbs_dat_i[22]       E    M����P wbs_dat_i[23]       E    �����P wbs_dat_i[24]       E    ����P wbs_dat_i[25]       E    ���P wbs_dat_i[26]       E    d*���P wbs_dat_i[27]       E    �>���P wbs_dat_i[28]       E    �R���P wbs_dat_i[29]       E    	����P la_oen[0]       E    	4����P wbs_dat_i[30]       E    	z����P wbs_dat_i[31]       E    e����P wbs_adr_i[20]       E    �"���P wbs_adr_i[21]       E    �6���P wbs_adr_i[22]       E    6J���P wbs_adr_i[23]       E    |^���P wbs_adr_i[24]       E    �����P wbs_adr_i[25]       E    ����P wbs_adr_i[26]       E    L����P wbs_adr_i[27]       E    �����P wbs_adr_i[28]       E    �����P wbs_adr_i[29]       E    
2���P la_oen[1]       E    	>���P wbs_adr_i[30]       E    	cR���P wbs_adr_i[31]       E    
bz���P la_oen[2]       E    
�����P la_oen[3]       E    �V���P wbs_dat_o[17]       E    j���P wbs_dat_o[18]       E    N~���P wbs_dat_o[19]       E    
����P la_oen[4]       E    �����P wbs_dat_o[20]       E    �����P wbs_dat_o[21]       E    ����P wbs_dat_o[22]       E    e���P wbs_dat_o[23]       E    ����P wbs_dat_o[24]       E    �^���P wbs_dat_o[25]       E    5r���P wbs_dat_o[26]       E    {����P wbs_dat_o[27]       E    �����P wbs_dat_o[28]       E    	����P wbs_dat_o[29]       E    	�f���P la_data_in[0]       E    	K����P wbs_dat_o[30]       E    	�
���P wbs_dat_o[31]       E    	�z���P la_data_in[1]       E    
5����P la_data_in[2]       E    
y����P la_data_in[3]       E    
�����P la_data_in[4]       E    ����P la_data_in[5]       E    	�����P la_data_out[0]      E    
����P la_data_out[1]      E    
K���P la_data_out[2]      E    
�2���P la_data_out[3]      E    
�F���P la_data_out[4]      E    Z���P la_data_out[5]      E    ٲ���P wbs_adr_i[18]       E    �����P wbs_dat_i[17]       E    �6���P la_data_in[23]      E    2J���P la_data_in[24]      E    4����P la_oen[5]       E    z����P la_oen[6]       E    ����P la_oen[7]       E    &���P la_oen[8]       E    K:���P la_oen[9]       E    x^���P la_data_in[25]      E    �����P la_data_in[11]      E    �����P la_data_in[12]      E    3���P la_data_in[13]      E    y���P la_data_in[14]      E    L���P la_data_in[6]       E    �Z���P la_data_in[7]       E    �n���P la_data_in[8]       E    ����P la_data_in[9]       E    �.���P la_data_in[15]      E    y����P la_data_out[10]       E    ����P la_data_out[11]       E    N���P la_data_out[12]       E    Jb���P la_data_out[13]       E    �v���P la_data_out[14]       E    ֊���P la_data_out[15]       E    ����P la_data_out[16]       E    `����P la_data_out[17]       E    �����P la_data_out[18]       E    ����P la_data_out[19]       E    B���P la_data_in[16]      E    3"���P la_data_out[20]       E    wj���P la_data_out[21]       E    �~���P la_data_out[22]       E    ����P la_data_out[23]       E    I����P la_data_out[24]       E    �����P la_data_out[25]       E    I����P la_data_in[17]      E    �����P la_data_in[18]      E    ղ���P la_data_in[19]      E    b����P la_data_in[10]      E    cn���P la_data_out[6]      E    �����P la_data_out[7]      E    �����P la_data_out[8]      E    3����P la_data_out[9]      E    ����P la_data_in[20]      E    �N���P la_oen[10]      E    Ֆ���P la_oen[11]      E    ����P la_oen[12]      E    a����P la_oen[13]      E    �����P la_oen[14]      E    �����P la_oen[15]      E    2.���P la_oen[16]      E    xB���P la_oen[17]      E    �V���P la_oen[18]      E    j���P la_oen[19]      E    `���P la_data_in[21]      E    J~���P la_oen[20]      E    �����P la_oen[21]      E    �����P la_oen[22]      E    ����P la_oen[23]      E    a���P la_oen[24]      E    �J���P la_oen[25]      E    �"���P la_data_in[22]      E    �����P la_data_in[37]      E    ����P la_data_in[38]      E    H���P la_data_in[39]      E    і���P la_oen[44]      E    ����P la_data_out[26]       E    ���P la_data_out[27]       E    `*���P la_data_out[28]       E    �>���P la_data_out[29]       E    �Z���P la_data_in[40]      E    ����P la_data_out[30]       E    0����P la_data_out[31]       E    v����P la_data_out[32]       E    �����P la_data_out[33]       E    ����P la_data_out[34]       E    G���P la_data_out[35]       E    �2���P la_data_out[36]       E    �F���P la_data_out[37]       E    Z���P la_data_out[38]       E    _n���P la_data_out[39]       E    �n���P la_data_in[41]      E    �����P la_data_out[40]       E    �����P la_data_out[41]       E    /����P la_data_out[42]       E    u����P la_data_out[43]       E    �:���P la_data_out[44]       E     N���P la_data_out[45]       E    Fb���P la_data_out[46]       E    ����P la_data_in[42]      E    ^����P la_data_in[43]      E    �����P la_data_in[44]      E    �����P la_data_in[45]      E    /���P la_data_in[46]      E    ����P la_oen[45]      E    ����P la_oen[37]      E    0����P la_oen[38]      E    t����P la_oen[39]      E    �����P la_oen[36]      E    ����P la_oen[40]      E    &���P la_oen[41]      E    G:���P la_oen[42]      E    �����P la_data_in[26]      E    ����P la_data_in[27]      E    H����P la_data_in[28]      E    �����P la_data_in[29]      E    �N���P la_oen[43]      E    �����P la_data_in[30]      E    >���P la_data_in[31]      E    _R���P la_data_in[32]      E    �f���P la_data_in[33]      E    �z���P la_data_in[34]      E    /����P la_data_in[35]      E    �^���P la_oen[26]      E    1r���P la_oen[27]      E    w����P la_oen[28]      E    �����P la_oen[29]      E    u����P la_data_in[36]      E    ����P la_oen[30]      E    G����P la_oen[31]      E    �
���P la_oen[32]      E    ����P la_oen[33]      E    2���P la_oen[34]      E    ^z���P la_oen[35]      E    ]����P la_oen[46]      E    �����P la_oen[47]      E    �����P la_oen[48]      E    ..���P la_oen[49]      E    tB���P la_oen[50]      E    �V���P la_oen[51]      E     j���P la_oen[52]      E    D����P la_oen[53]      E    �����P la_oen[54]      E    �����P la_oen[55]      E    ����P la_oen[56]      E    ]���P la_oen[57]      E    �J���P la_oen[58]      E    �^���P la_oen[59]      E    -r���P la_oen[60]      E    s����P la_oen[61]      E    �����P la_oen[62]      E    �����P la_oen[63]      E    C����P la_oen[64]      E    �
���P la_oen[65]      E    ����P la_oen[66]      E    u���P la_data_in[47]      E    �.���P la_data_in[48]      E    �v���P la_data_in[49]      E    E����P la_data_in[50]      E    �����P la_data_in[51]      E    Ѳ���P la_data_in[52]      E    ����P la_data_in[53]      E    \���P la_data_in[54]      E    �"���P la_data_in[55]      E    �6���P la_data_in[56]      E    .J���P la_data_in[57]      E    t^���P la_data_in[58]      E    �����P la_data_in[59]      E    �����P la_data_in[60]      E    D����P la_data_in[61]      E    �����P la_data_in[62]      E    �*���P la_data_in[63]      E    �v���P la_data_out[47]       E    Ҋ���P la_data_out[48]       E    ����P la_data_out[49]       E    >���P la_data_in[64]      E    \����P la_data_out[50]       E    �����P la_data_out[51]       E    ����P la_data_out[52]       E    /"���P la_data_out[53]       E    sj���P la_data_out[54]       E    �~���P la_data_out[55]       E    �����P la_data_out[56]       E    E����P la_data_out[57]       E    �����P la_data_out[58]       E    ����P la_data_out[59]       E    [R���P la_data_in[65]      E    ���P la_data_out[60]       E    \*���P la_data_out[61]       E    �>���P la_data_out[62]       E    ����P la_data_out[63]       E    ,����P la_data_out[64]       E    r����P la_data_out[65]       E    �����P la_data_out[66]       E    �f���P la_data_in[66]      E    D���P la_data_in[72]      E    �Z���P la_data_in[73]      E    �n���P la_data_in[74]      E    ����P la_data_in[75]      E    Z����P la_data_in[76]      E    �����P la_data_in[77]      E    �����P la_data_in[78]      E    +���P la_data_in[79]      E    q���P la_data_in[80]      E    �.���P la_data_in[81]      E    �v���P la_data_in[82]      E     A����P la_data_in[83]      E     �����P la_data_in[84]      E     Ͳ���P la_data_in[85]      E    !����P la_data_in[86]      E    !X���P la_data_in[87]      E    q����P la_data_in[69]      E    �����P la_data_in[70]      E    f���P la_oen[67]      E    Zz���P la_oen[68]      E    �����P la_oen[69]      E    ����P la_oen[70]      E    ,����P la_oen[71]      E    p����P la_oen[72]      E    ����P la_oen[73]      E    �&���P la_oen[74]      E    C:���P la_oen[75]      E    �N���P la_oen[76]      E    ͖���P la_oen[77]      E    ����P la_oen[78]      E    Y����P la_oen[79]      E    �����P la_oen[80]      E    ����P la_oen[81]      E     *.���P la_oen[82]      E     pB���P la_oen[83]      E     �V���P la_oen[84]      E     �j���P la_oen[85]      E    !@����P la_oen[86]      E    �����P la_data_out[67]       E    C���P la_data_out[68]       E    �2���P la_data_out[69]       E    �����P la_data_in[71]      E    �F���P la_data_out[70]       E    Z���P la_data_out[71]       E    Y����P la_data_out[72]       E    �����P la_data_out[73]       E    �����P la_data_out[74]       E    +����P la_data_out[75]       E    q����P la_data_out[76]       E    �:���P la_data_out[77]       E    �N���P la_data_out[78]       E    Bb���P la_data_out[79]       E    �z���P la_data_in[67]      E    �v���P la_data_out[80]       E    Ί���P la_data_out[81]       E     ����P la_data_out[82]       E     X����P la_data_out[83]       E     �����P la_data_out[84]       E     ����P la_data_out[85]       E    !)V���P la_data_out[86]       E    +����P la_data_in[68]      E    !�6���P la_data_in[89]      E    !�����P la_oen[87]      E    !�����P la_oen[88]      E    "����P la_oen[89]      E    "Y���P la_oen[90]      E    "�J���P la_oen[91]      E    "�^���P la_oen[92]      E    #)r���P la_oen[93]      E    #o����P la_oen[94]      E    #�����P la_oen[95]      E    #�����P la_oen[96]      E    $?����P la_oen[97]      E    $�
���P la_oen[98]      E    $����P la_oen[99]      E    %'����P la_data_in[101]       E    %m����P la_data_in[102]       E    %�����P la_data_in[103]       E    %�����P la_data_in[104]       E    &>F���P la_data_in[105]       E    &�Z���P la_data_in[106]       E    &�n���P la_data_in[107]       E    $�z���P la_data_in[100]       E    "*J���P la_data_in[90]      E    "n����P la_data_in[91]      E    "�����P la_data_in[92]      E    "�����P la_data_in[93]      E    #@����P la_data_in[94]      E    #�����P la_data_in[95]      E    #�*���P la_data_in[96]      E    $>���P la_data_in[97]      E    $WR���P la_data_in[98]      E    $�f���P la_data_in[99]      E    $�
���P la_data_out[100]      E    %?���P la_data_out[101]      E    %�2���P la_data_out[102]      E    %�F���P la_data_out[103]      E    &Z���P la_data_out[104]      E    "����P la_data_out[92]       E    &U����P la_data_out[105]      E    #���P la_data_out[93]       E    &�����P la_data_out[106]      E    #X*���P la_data_out[94]       E    #�>���P la_data_out[95]       E    &�����P la_data_out[107]      E    #����P la_data_out[96]       E    $(����P la_data_out[97]       E    $n����P la_data_out[98]       E    $�����P la_data_out[99]       E    "�����P la_data_out[91]       E    %f���P la_oen[100]       E    %Vz���P la_oen[101]       E    %�����P la_oen[102]       E    %����P la_oen[103]       E    &(����P la_oen[104]       E    &l����P la_oen[105]       E    &����P la_oen[106]       E    !oj���P la_data_out[87]       E    !�~���P la_data_out[88]       E    !�����P la_data_out[89]       E    !�"���P la_data_in[88]      E    "A����P la_data_out[90]       E    *%V���P la_data_out[119]      E    *����P la_data_in[119]       E    *kj���P la_data_out[120]      E    *�~���P la_data_out[121]      E    *�����P la_data_out[122]      E    +=����P la_data_out[123]      E    )=����P la_data_in[116]       E    )�����P la_data_in[117]       E    ('���P la_data_in[112]       E    +�����P la_data_out[124]      E    +����P la_data_out[125]      E    ,���P la_data_out[126]      E    ,T*���P la_data_out[127]      E    'm����P la_data_out[109]      E    '?:���P la_oen[108]       E    '�����P la_oen[109]       E    *T���P la_data_in[120]       E    'ɖ���P la_oen[110]       E    *�"���P la_data_in[121]       E    (����P la_oen[111]       E    (U����P la_oen[112]       E    (�����P la_oen[113]       E    (����P la_oen[114]       E    )&.���P la_oen[115]       E    )lB���P la_oen[116]       E    )�V���P la_oen[117]       E    )�j���P la_oen[118]       E    *<����P la_oen[119]       E    *�6���P la_data_in[122]       E    +&J���P la_data_in[123]       E    *�����P la_oen[120]       E    *�����P la_oen[121]       E    +����P la_oen[122]       E    +S6���P la_oen[123]       E    +�J���P la_oen[124]       E    +�^���P la_oen[125]       E    ,%r���P la_oen[126]       E    ,k����P la_oen[127]       E    +j����P la_data_in[124]       E    +�����P la_data_in[125]       E    +�����P la_data_in[126]       E    ,<����P la_data_in[127]       E    )ɲ���P la_data_in[118]       E    ,�����P user_clock2       E    '�:���P la_data_out[110]      E    '�N���P la_data_out[111]      E    (m���P la_data_in[113]       E    (�.���P la_data_in[114]       E    (>b���P la_data_out[112]      E    (�v���P la_data_out[113]      E    '����P la_data_in[108]       E    ''����P la_data_out[108]      E    'V����P la_data_in[109]       E    (Ⱦ���P la_data_out[114]      E    '�����P la_data_in[110]       E    (�v���P la_data_in[115]       E    &�&���P la_oen[107]       E    )����P la_data_out[115]      E    )T����P la_data_out[116]      E    '�����P la_data_in[111]       E    )�����P la_data_out[117]      E    )����P la_data_out[118]      H   ,�������������� ,������ ,�������������      H   ,������������� ,Ÿ��� ,Ÿ�����������      H   ,�����������ռ ,װ��ռ ,װ���������      H   ,������������� ,����� ,����������      H   ,���$������$���� ,������ ,��������$���      H   ,��,�����,���� -����� -������,���      H   ,��m4���$��m4���� -����� -����$��m4���$      H   ,��[<��p,��[<��{� -1���{� -1���p,��[<��p,      H    Fb���� 
vccd1       H    Fb���� 
vssd1       H    Fb���� 
vccd2       H    Fb���� 
vssd2       H    Fb���� 
vdda1       H    Fb���� 
vssa1       H    Fb���  
vdda2       H    Fb��v 
vssa2    	   B   !        *�� + *�� 5 *�� 5   	   B   !        +|; �� +�� ��      B  , , *�p 0 *�p � *� � *� 0 *�p 0      B  , , *�� 0 *�� � *�� � *�� 0 *�� 0      B  , , *�p 0 *�p � *� � *� 0 *�p 0      B  , , *��  *�� � *�� � *��  *��       B  , , *�p  *�p � *� � *�  *�p       B  , , *�� � *�� � *�� � *�� � *�� �      B  , , *�p � *�p � *� � *� � *�p �      B  , , +�& �` +�& �
 +�� �
 +�� �` +�& �`      B  , , +�� �` +�� �
 +�= �
 +�= �` +�� �`      B  , , +�& �` +�& �
 +�� �
 +�� �` +�& �`      B  , , +�� �2 +�� �� +�= �� +�= �2 +�� �2      B  , , +�& �2 +�& �� +�� �� +�� �2 +�& �2      B  , , +�� � +�� �� +�= �� +�= � +�� �      B  , , +�& � +�& �� +�� �� +�� � +�& �      E  , , +8� �
 +8� �� +9x �� +9x �
 +8� �
      E  , , +j( G +j( � +j� � +j� G +j( G      E  , , +k� � +k� M +lO M +lO � +k� �      E  , , +k� G +k� � +lO � +lO G +k� G      E  , , +j' � +j' K +j� K +j� � +j' �      E  , , +:s �z +:s � +;	 � +;	 �z +:s �z      E  , , +:s �
 +:s �� +;	 �� +;	 �
 +:s �
      E  , , +8� �x +8� � +9w � +9w �x +8� �x      E  , , *�� 1h *�� 1� *�Z 1� *�Z 1h *�� 1h      E  , , *�U /� *�U 0n *�� 0n *�� /� *�U /�      E  , , *�U 1h *�U 1� *�� 1� *�� 1h *�U 1h      E  , , *�� /� *�� 0l *�Y 0l *�Y /� *�� /�      