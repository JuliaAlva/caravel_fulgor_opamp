* NGSPICE file created from opamp_v1.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_YT7TV5 a_n1268_n718# a_1147_n815# VSUBS a_n269_21#
+ a_1210_n718# a_85_21# a_n859_n815# a_793_n815# a_1210_118# a_n977_21# a_n505_n815#
+ a_974_118# a_n442_118# a_148_n718# a_n859_21# a_n151_n815# a_n1386_n718# a_1265_n815#
+ a_n1032_n718# a_911_n815# a_n1032_118# a_n88_n718# a_n796_118# a_502_118# a_n977_n815#
+ a_n623_n815# a_266_118# a_n88_118# a_266_n718# a_n1504_n718# a_n1386_118# a_1383_21#
+ a_1383_n815# a_856_118# a_n1150_n718# a_1265_21# a_n324_118# a_n206_n718# a_738_n718#
+ a_1147_21# a_30_n718# a_n741_n815# a_1029_21# a_384_n718# a_1446_118# a_n914_118#
+ a_n33_21# a_n678_118# a_321_21# a_n1449_n815# a_148_118# a_n678_n718# a_203_21#
+ a_439_n815# a_n324_n718# a_85_n815# a_856_n718# a_n1095_n815# a_502_n718# a_n1504_118#
+ a_793_21# a_n1268_118# a_911_21# a_738_118# a_675_21# a_n206_118# a_n1331_21# a_1328_n718#
+ a_557_21# a_n1095_21# a_n1213_21# a_n1213_n815# a_439_21# a_n796_n718# a_557_n815#
+ a_n442_n718# a_974_n718# a_203_n815# a_30_118# a_1328_118# a_620_n718# a_n269_n815#
+ a_1092_118# a_n560_118# a_n151_21# a_1029_n815# a_1446_n718# a_n914_n718# a_n1449_21#
+ a_n1331_n815# a_1092_n718# a_675_n815# a_n560_n718# a_321_n815# a_n741_21# a_n33_n815#
+ a_n1150_118# a_n387_n815# a_620_118# a_n623_21# w_n1642_n937# a_384_118# a_n387_21#
+ a_n505_21#
X0 a_n796_118# a_n859_21# a_n914_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X1 a_266_118# a_203_21# a_148_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X2 a_1092_118# a_1029_21# a_974_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X3 a_n442_n718# a_n505_n815# a_n560_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X4 a_n678_118# a_n741_21# a_n796_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X5 a_856_118# a_793_21# a_738_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X6 a_148_n718# a_85_n815# a_30_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X7 a_1210_n718# a_1147_n815# a_1092_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X8 a_n1386_118# a_n1449_21# a_n1504_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X9 a_n560_118# a_n623_21# a_n678_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X10 a_738_118# a_675_21# a_620_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X11 a_1092_n718# a_1029_n815# a_974_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X12 a_n1268_118# a_n1331_21# a_n1386_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X13 a_n1150_118# a_n1213_21# a_n1268_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X14 a_1446_118# a_1383_21# a_1328_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X15 a_n324_118# a_n387_21# a_n442_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X16 a_1328_118# a_1265_21# a_1210_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X17 a_n914_n718# a_n977_n815# a_n1032_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X18 a_n324_n718# a_n387_n815# a_n442_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X19 a_n796_n718# a_n859_n815# a_n914_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X20 a_n206_n718# a_n269_n815# a_n324_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X21 a_n1032_118# a_n1095_21# a_n1150_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X22 a_n206_118# a_n269_21# a_n324_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X23 a_n88_n718# a_n151_n815# a_n206_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X24 a_n678_n718# a_n741_n815# a_n796_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X25 a_620_n718# a_557_n815# a_502_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X26 a_n88_118# a_n151_21# a_n206_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X27 a_n560_n718# a_n623_n815# a_n678_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X28 a_148_118# a_85_21# a_30_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X29 a_974_118# a_911_21# a_856_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X30 a_n1032_n718# a_n1095_n815# a_n1150_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X31 a_502_n718# a_439_n815# a_384_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X32 a_384_n718# a_321_n815# a_266_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X33 a_1446_n718# a_1383_n815# a_1328_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X34 a_974_n718# a_911_n815# a_856_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X35 a_1328_n718# a_1265_n815# a_1210_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X36 a_n1386_n718# a_n1449_n815# a_n1504_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X37 a_266_n718# a_203_n815# a_148_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X38 a_n1268_n718# a_n1331_n815# a_n1386_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X39 a_30_n718# a_n33_n815# a_n88_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X40 a_30_118# a_n33_21# a_n88_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X41 a_n1150_n718# a_n1213_n815# a_n1268_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X42 a_n442_118# a_n505_21# a_n560_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X43 a_620_118# a_557_21# a_502_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X44 a_502_118# a_439_21# a_384_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X45 a_856_n718# a_793_n815# a_738_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X46 a_n914_118# a_n977_21# a_n1032_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X47 a_738_n718# a_675_n815# a_620_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X48 a_384_118# a_321_21# a_266_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X49 a_1210_118# a_1147_21# a_1092_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
.ends

.subckt sky130_fd_pr__nfet_01v8_8HUREQ VSUBS a_n269_21# a_n914_109# a_n678_109# a_n269_n797#
+ a_85_21# a_148_109# a_n678_n709# a_n324_n709# a_856_n709# a_n859_21# a_502_n709#
+ a_738_109# a_675_n797# a_n206_109# a_n33_n797# a_321_n797# a_n387_n797# a_n796_n709#
+ a_30_109# a_n442_n709# a_620_n709# a_n560_109# a_n859_n797# a_n505_n797# a_793_n797#
+ a_n914_n709# a_n151_n797# a_n560_n709# a_n33_21# a_384_109# a_620_109# a_321_21#
+ a_n623_n797# a_203_21# a_793_21# a_n442_109# a_675_21# a_148_n709# a_557_21# a_n741_n797#
+ w_n1052_n919# a_439_21# a_n796_109# a_502_109# a_n88_n709# a_266_109# a_n88_109#
+ a_439_n797# a_266_n709# a_n151_21# a_85_n797# a_856_109# a_n324_109# a_n741_21#
+ a_n206_n709# a_738_n709# a_n623_21# a_30_n709# a_n505_21# a_n387_21# a_203_n797#
+ a_557_n797# a_384_n709#
X0 a_30_109# a_n33_21# a_n88_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X1 a_n442_109# a_n505_21# a_n560_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X2 a_620_109# a_557_21# a_502_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X3 a_502_109# a_439_21# a_384_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X4 a_856_n709# a_793_n797# a_738_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X5 a_738_n709# a_675_n797# a_620_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X6 a_384_109# a_321_21# a_266_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X7 a_n796_109# a_n859_21# a_n914_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X8 a_266_109# a_203_21# a_148_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X9 a_n442_n709# a_n505_n797# a_n560_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X10 a_n678_109# a_n741_21# a_n796_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X11 a_856_109# a_793_21# a_738_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X12 a_148_n709# a_85_n797# a_30_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X13 a_n560_109# a_n623_21# a_n678_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X14 a_738_109# a_675_21# a_620_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X15 a_n324_n709# a_n387_n797# a_n442_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X16 a_n324_109# a_n387_21# a_n442_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X17 a_n796_n709# a_n859_n797# a_n914_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X18 a_n206_n709# a_n269_n797# a_n324_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X19 a_n206_109# a_n269_21# a_n324_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X20 a_n88_n709# a_n151_n797# a_n206_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X21 a_n678_n709# a_n741_n797# a_n796_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X22 a_620_n709# a_557_n797# a_502_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X23 a_n88_109# a_n151_21# a_n206_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X24 a_148_109# a_85_21# a_30_109# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X25 a_n560_n709# a_n623_n797# a_n678_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X26 a_502_n709# a_439_n797# a_384_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X27 a_384_n709# a_321_n797# a_266_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X28 a_266_n709# a_203_n797# a_148_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X29 a_30_n709# a_n33_n797# a_n88_n709# VSUBS sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_BLS9H9 VSUBS c1_n1841_n1500# m3_n1941_n1600#
X0 c1_n1841_n1500# m3_n1941_n1600# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.755e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_YC9MKB VSUBS a_502_n300# a_n151_n397# a_n623_n397#
+ a_n796_n300# a_n442_n300# a_620_n300# a_n914_n300# a_n741_n397# a_n560_n300# w_n1052_n519#
+ a_85_n397# a_439_n397# a_148_n300# a_557_n397# a_203_n397# a_n88_n300# a_n269_n397#
+ a_266_n300# a_675_n397# a_n206_n300# a_738_n300# a_n33_n397# a_321_n397# a_30_n300#
+ a_n387_n397# a_384_n300# a_n859_n397# a_793_n397# a_n678_n300# a_n505_n397# a_n324_n300#
+ a_856_n300#
X0 a_266_n300# a_203_n397# a_148_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X1 a_30_n300# a_n33_n397# a_n88_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X2 a_856_n300# a_793_n397# a_738_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X3 a_738_n300# a_675_n397# a_620_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X4 a_n442_n300# a_n505_n397# a_n560_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X5 a_148_n300# a_85_n397# a_30_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X6 a_n324_n300# a_n387_n397# a_n442_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X7 a_n796_n300# a_n859_n397# a_n914_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X8 a_n206_n300# a_n269_n397# a_n324_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X9 a_n88_n300# a_n151_n397# a_n206_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X10 a_n678_n300# a_n741_n397# a_n796_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X11 a_620_n300# a_557_n397# a_502_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X12 a_n560_n300# a_n623_n397# a_n678_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X13 a_502_n300# a_439_n397# a_384_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X14 a_384_n300# a_321_n397# a_266_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
.ends

.subckt sky130_fd_pr__nfet_01v8_THKFL3 VSUBS a_n73_n150# w_n211_n360# a_15_n150#
X0 a_15_n150# a_n33_n238# a_n73_n150# VSUBS sky130_fd_pr__nfet_01v8 w=1.5e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_YCMRKB a_262_21# a_679_118# a_2803_118# VSUBS a_2567_118#
+ a_n446_n815# a_n2924_21# a_n2035_118# a_n147_118# a_380_n815# a_n92_n815# a_144_21#
+ a_2858_n815# a_n2688_21# a_n2979_n718# a_n2806_21# a_970_21# a_1977_n718# a_1206_n815#
+ a_n1327_n718# a_n2625_n718# a_2504_n815# a_n1799_118# a_1623_n718# a_2921_n718#
+ a_852_21# a_1505_118# a_n1862_n815# a_1269_118# a_n29_n718# a_n2625_118# a_n737_118#
+ a_2150_n815# a_n918_n815# a_n1390_21# a_n2271_n718# a_852_n815# a_734_21# a_n2389_118#
+ a_207_118# a_498_21# a_n29_118# a_n1272_21# a_n2098_n815# a_616_21# a_207_n718#
+ a_n564_n815# a_n210_n815# a_n1154_21# a_n1799_n718# a_1678_n815# a_n1980_21# a_n1327_118#
+ a_1859_118# a_1324_n815# a_n1445_n718# a_n2743_n718# a_2622_n815# a_n1036_21# a_n2979_118#
+ a_1741_n718# a_n1862_21# a_n1980_n815# a_2449_118# a_n1091_118# a_n1091_n718# a_n1744_21#
+ a_970_n815# a_n2216_n815# a_561_118# a_n147_n718# a_n210_21# a_n1917_118# a_679_n718#
+ a_n1626_21# a_325_n718# a_n1917_n718# a_n682_n815# a_n1508_21# a_1796_n815# a_n2507_118#
+ a_n682_21# a_n1681_118# a_n619_118# a_1442_n815# a_n1563_n718# a_n2861_n718# a_2740_n815#
+ a_n800_21# a_2150_21# a_2449_n718# a_n619_n718# a_n564_21# a_1151_118# a_26_n815#
+ a_2032_21# a_n2688_n815# a_n2271_118# a_n383_118# a_n1036_n815# a_n2334_n815# a_n446_21#
+ a_2095_n718# a_n265_n718# a_n800_n815# a_n1209_118# a_797_n718# a_2740_21# a_n328_21#
+ a_443_n718# a_1914_n815# a_1741_118# a_2622_21# a_n2861_118# a_n973_118# a_1560_n815#
+ a_26_21# a_2386_21# a_n1681_n718# a_n1508_n815# a_2504_21# a_n2806_n815# a_443_118#
+ a_1269_n718# a_2567_n718# a_n737_n718# a_2331_118# a_n918_21# a_2268_21# a_2213_n718#
+ a_2095_118# a_915_n718# a_n1154_n815# a_n2452_n815# a_498_n815# a_n383_n718# a_n1563_118#
+ a_144_n815# a_561_n718# a_2858_21# a_1033_118# a_2921_118# a_n501_118# a_797_118#
+ a_n2153_118# a_n265_118# a_2685_118# a_n1626_n815# a_n2924_n815# a_n2389_n718# a_2268_n815#
+ a_1387_n718# a_2685_n718# a_n855_n718# a_89_118# a_n2035_n718# a_616_n815# a_1560_21#
+ a_2331_n718# a_1033_n718# a_n501_n718# a_n1272_n815# a_n2570_n815# a_1623_118# a_1442_21#
+ a_1387_118# a_n328_n815# a_n2570_21# a_n2743_118# a_n855_118# a_262_n815# a_1324_21#
+ a_325_118# a_n2452_21# a_2213_118# a_1859_n718# a_1088_21# a_n1209_n718# a_n2507_n718#
+ a_1505_n718# a_1206_21# a_2803_n718# w_n3117_n937# a_n2334_21# a_1088_n815# a_n1744_n815#
+ a_2386_n815# a_n92_21# a_1977_118# a_1796_21# a_n1445_118# a_n973_n718# a_2032_n815#
+ a_n2098_21# a_380_21# a_n2153_n718# a_734_n815# a_n2216_21# a_1914_21# a_1151_n718#
+ a_915_118# a_1678_21# a_89_n718# a_n1390_n815#
X0 a_n1445_n718# a_n1508_n815# a_n1563_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X1 a_2567_118# a_2504_21# a_2449_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X2 a_n501_118# a_n564_21# a_n619_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X3 a_1269_n718# a_1206_n815# a_1151_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X4 a_n1917_118# a_n1980_21# a_n2035_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X5 a_n737_n718# a_n800_n815# a_n855_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X6 a_1387_118# a_1324_21# a_1269_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X7 a_n383_118# a_n446_21# a_n501_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X8 a_n2271_118# a_n2334_21# a_n2389_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X9 a_n619_n718# a_n682_n815# a_n737_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X10 a_n1799_118# a_n1862_21# a_n1917_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X11 a_1269_118# a_1206_21# a_1151_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X12 a_n265_118# a_n328_21# a_n383_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X13 a_n1091_118# a_n1154_21# a_n1209_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X14 a_2331_n718# a_2268_n815# a_2213_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X15 a_n2153_118# a_n2216_21# a_n2271_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X16 a_443_n718# a_380_n815# a_325_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X17 a_2921_n718# a_2858_n815# a_2803_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X18 a_1033_n718# a_970_n815# a_915_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X19 a_443_118# a_380_21# a_325_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X20 a_2331_118# a_2268_21# a_2213_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X21 a_n147_118# a_n210_21# a_n265_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X22 a_2213_n718# a_2150_n815# a_2095_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X23 a_n973_118# a_n1036_21# a_n1091_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X24 a_325_n718# a_262_n815# a_207_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X25 a_2803_n718# a_2740_n815# a_2685_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X26 a_1859_118# a_1796_21# a_1741_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X27 a_915_n718# a_852_n815# a_797_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X28 a_n2271_n718# a_n2334_n815# a_n2389_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X29 a_325_118# a_262_21# a_207_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X30 a_n2861_n718# a_n2924_n815# a_n2979_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X31 a_1151_118# a_1088_21# a_1033_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X32 a_2095_n718# a_2032_n815# a_1977_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X33 a_1859_n718# a_1796_n815# a_1741_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X34 a_207_n718# a_144_n815# a_89_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X35 a_2213_118# a_2150_21# a_2095_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X36 a_2685_n718# a_2622_n815# a_2567_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X37 a_797_n718# a_734_n815# a_679_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X38 a_n1327_n718# a_n1390_n815# a_n1445_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X39 a_89_118# a_26_21# a_n29_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X40 a_n1917_n718# a_n1980_n815# a_n2035_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X41 a_n2153_n718# a_n2216_n815# a_n2271_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X42 a_n29_n718# a_n92_n815# a_n147_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X43 a_n2743_n718# a_n2806_n815# a_n2861_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X44 a_n737_118# a_n800_21# a_n855_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X45 a_207_118# a_144_21# a_89_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X46 a_n2625_118# a_n2688_21# a_n2743_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X47 a_2567_n718# a_2504_n815# a_2449_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X48 a_679_n718# a_616_n815# a_561_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X49 a_n1209_n718# a_n1272_n815# a_n1327_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X50 a_2095_118# a_2032_21# a_1977_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X51 a_n1799_n718# a_n1862_n815# a_n1917_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X52 a_n619_118# a_n682_21# a_n737_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X53 a_n2507_118# a_n2570_21# a_n2625_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X54 a_n1327_118# a_n1390_21# a_n1445_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X55 a_n2389_118# a_n2452_21# a_n2507_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X56 a_n1209_118# a_n1272_21# a_n1327_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X57 a_89_n718# a_26_n815# a_n29_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X58 a_n2035_n718# a_n2098_n815# a_n2153_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X59 a_2449_118# a_2386_21# a_2331_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X60 a_561_118# a_498_21# a_443_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X61 a_n2625_n718# a_n2688_n815# a_n2743_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X62 a_2449_n718# a_2386_n815# a_2331_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X63 a_n501_n718# a_n564_n815# a_n619_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X64 a_1977_118# a_1914_21# a_1859_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X65 a_n2507_n718# a_n2570_n815# a_n2625_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X66 a_n2861_118# a_n2924_21# a_n2979_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X67 a_n383_n718# a_n446_n815# a_n501_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X68 a_n2389_n718# a_n2452_n815# a_n2507_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X69 a_n855_118# a_n918_21# a_n973_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X70 a_n1681_118# a_n1744_21# a_n1799_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X71 a_n2743_118# a_n2806_21# a_n2861_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X72 a_n2035_118# a_n2098_21# a_n2153_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X73 a_n265_n718# a_n328_n815# a_n383_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X74 a_n855_n718# a_n918_n815# a_n973_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X75 a_1033_118# a_970_21# a_915_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X76 a_1151_n718# a_1088_n815# a_1033_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X77 a_1741_n718# a_1678_n815# a_1623_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X78 a_2921_118# a_2858_21# a_2803_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X79 a_n1563_118# a_n1626_21# a_n1681_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X80 a_n147_n718# a_n210_n815# a_n265_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X81 a_915_118# a_852_21# a_797_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X82 a_1623_n718# a_1560_n815# a_1505_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X83 a_1741_118# a_1678_21# a_1623_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X84 a_2803_118# a_2740_21# a_2685_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X85 a_n1445_118# a_n1508_21# a_n1563_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X86 a_561_n718# a_498_n815# a_443_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X87 a_n1091_n718# a_n1154_n815# a_n1209_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X88 a_n1681_n718# a_n1744_n815# a_n1799_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X89 a_1505_n718# a_1442_n815# a_1387_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X90 a_797_118# a_734_21# a_679_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X91 a_1623_118# a_1560_21# a_1505_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X92 a_n973_n718# a_n1036_n815# a_n1091_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X93 a_2685_118# a_2622_21# a_2567_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X94 a_n1563_n718# a_n1626_n815# a_n1681_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X95 a_1387_n718# a_1324_n815# a_1269_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X96 a_1977_n718# a_1914_n815# a_1859_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X97 a_679_118# a_616_21# a_561_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X98 a_1505_118# a_1442_21# a_1387_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X99 a_n29_118# a_n92_21# a_n147_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
.ends

.subckt sky130_fd_pr__nfet_01v8_8JUMX6 a_n341_n1097# VSUBS a_n4041_21# a_3951_21#
+ a_695_21# a_4543_21# a_n843_109# a_5135_21# a_n3951_109# a_933_109# a_4041_109#
+ a_n341_21# a_2027_n1097# a_4691_21# a_n2767_109# a_n5431_n1009# a_n1969_21# a_5283_21#
+ a_4929_n1009# a_3063_n1097# a_n3507_n1009# a_843_21# a_1139_21# a_n399_109# a_2857_109#
+ a_n489_n1097# a_1139_n1097# a_547_n1097# a_n4543_n1009# a_n4691_109# a_n1081_n1097#
+ a_n1583_109# a_489_109# a_2175_n1097# a_991_21# a_1287_21# a_n1731_n1009# a_n2619_n1009#
+ a_4099_n1097# a_4781_109# a_193_n1009# a_n3655_n1009# a_5431_21# a_1673_109# a_3597_109#
+ a_1287_n1097# a_695_n1097# a_n5579_n1009# a_n2709_21# a_n5521_n1097# a_n4691_n1009#
+ a_3301_n1009# a_n2767_n1009# a_n2915_109# a_3005_109# a_n2857_21# a_1435_21# a_n4839_109#
+ a_5225_n1009# a_3803_n1097# a_n4633_n1097# a_n3449_21# a_n1081_21# a_2027_21# a_2413_n1009#
+ a_n547_109# a_n2709_n1097# a_n1879_n1009# a_1583_21# a_4929_109# a_n1821_n1097#
+ a_4337_n1009# a_n3597_21# a_2915_n1097# a_2175_21# a_n1731_109# a_637_109# a_n3745_n1097#
+ a_n4189_21# a_n5579_109# a_n3655_109# a_5373_n1009# a_4839_n1097# a_3951_n1097#
+ a_n4781_n1097# a_1525_n1009# a_933_n1009# a_3449_n1009# a_1821_109# a_n2857_n1097#
+ a_2561_n1009# a_n547_n1009# a_3745_109# a_n2027_n1009# a_4485_n1009# a_n489_21#
+ a_n3893_n1097# a_n3063_n1009# a_1731_21# a_n4395_109# a_n2471_109# a_4987_n1097#
+ a_n3745_21# a_n1287_109# a_1673_n1009# a_2323_21# a_n1969_n1097# a_n4337_21# a_3597_n1009#
+ a_45_n1009# a_n1139_n1009# a_n695_n1009# a_4839_21# a_2561_109# a_4485_109# a_n2175_n1009#
+ a_n3893_21# a_2471_21# a_1377_109# a_n3005_n1097# a_n4099_n1009# a_3211_n1097# a_n4485_21#
+ a_3063_21# a_193_109# a_n4041_n1097# a_n637_21# a_5135_n1097# a_n5077_21# a_4987_21#
+ a_n3803_109# a_n637_n1097# a_n1287_n1009# a_n2117_n1097# a_n2619_109# a_2323_n1097#
+ a_n785_21# a_n3153_n1097# a_4247_n1097# a_n5077_n1097# a_n1229_n1097# a_341_n1009#
+ a_2709_109# a_n3803_n1009# a_5283_n1097# a_n4633_21# a_3211_21# a_n785_n1097# a_1435_n1097#
+ a_n4543_109# a_n2265_n1097# a_843_n1097# a_n5225_21# a_n3359_109# a_n1435_109# a_2471_n1097#
+ a_3359_n1097# a_n4189_n1097# a_n4781_21# a_n2915_n1009# a_4395_n1097# a_n251_109#
+ a_n5373_21# a_n933_21# a_4633_109# a_1081_n1009# a_n4839_n1009# a_1525_109# a_3449_109#
+ a_n1377_n1097# a_n3951_n1009# a_341_109# a_1583_n1097# a_n1229_21# a_n45_21# a_n5283_109#
+ a_991_n1097# a_n2175_109# a_n4099_109# a_103_21# a_489_n1009# a_n1377_21# a_5373_109#
+ a_5521_n1009# a_2265_109# a_n4987_n1009# a_251_21# a_1879_21# a_4189_109# a_103_n1097#
+ a_n5521_21# a_n991_109# a_4633_n1009# a_n4929_n1097# a_n3507_109# a_n3211_n1009#
+ a_1081_109# a_n193_n1097# a_2709_n1009# a_45_109# a_251_n1097# a_1821_n1009# a_n5135_n1009#
+ a_n1525_21# a_n45_n1097# a_3745_n1009# a_n2117_21# a_n843_n1009# a_4781_n1009# a_n2323_n1009#
+ a_n1673_21# a_2619_21# a_n5431_109# a_n4247_109# a_n2323_109# a_n4247_n1009# a_n2265_21#
+ a_n1139_109# a_2857_n1009# a_n5283_n1009# a_2767_21# a_n1435_n1009# a_5521_109#
+ a_3893_n1009# a_3359_21# a_2413_109# a_4337_109# a_n991_n1009# a_n3359_n1009# a_1229_109#
+ a_n2471_n1009# a_n3301_n1097# a_399_n1097# a_1969_n1009# a_n3063_109# a_n4395_n1009#
+ a_n5225_n1097# a_n1821_21# a_5431_n1097# a_n933_n1097# a_3005_n1009# a_n2413_21#
+ a_4099_21# a_n2413_n1097# a_n103_n1009# a_n1583_n1009# a_3153_109# a_4041_n1009#
+ a_3507_n1097# a_n3005_21# a_2915_21# a_n4987_109# a_5077_109# a_n4337_n1097# a_n1879_109#
+ a_n4929_21# a_n2561_21# a_3507_21# a_4543_n1097# a_n5373_n1097# a_2117_n1009# a_n3153_21#
+ a_n695_109# a_n1525_n1097# a_3153_n1009# a_2619_n1097# a_1969_109# a_n3449_n1097#
+ a_1731_n1097# a_n251_n1009# a_399_21# a_3655_21# a_785_109# a_n2561_n1097# a_5077_n1009#
+ a_3655_n1097# a_1229_n1009# a_4247_21# a_n4485_n1097# a_637_n1009# a_n103_109# a_4691_n1097#
+ a_2265_n1009# a_n1673_n1097# a_4395_21# a_3893_109# a_4189_n1009# a_2767_n1097#
+ a_n5135_109# a_n3211_109# a_n3597_n1097# a_n3301_21# a_n2027_109# a_n193_21# a_1377_n1009#
+ a_785_n1009# a_547_21# a_3803_21# a_3301_109# a_5225_109# a_1879_n1097# a_n399_n1009#
+ a_2117_109#
X0 a_2413_n1009# a_2323_n1097# a_2265_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X1 a_4485_109# a_4395_21# a_4337_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X2 a_n1287_109# a_n1377_21# a_n1435_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X3 a_n1731_n1009# a_n1821_n1097# a_n1879_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X4 a_n103_109# a_n193_21# a_n251_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X5 a_4337_109# a_4247_21# a_4189_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X6 a_4485_n1009# a_4395_n1097# a_4337_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X7 a_785_n1009# a_695_n1097# a_637_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X8 a_45_n1009# a_n45_n1097# a_n103_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X9 a_3745_109# a_3655_21# a_3597_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X10 a_4337_n1009# a_4247_n1097# a_4189_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X11 a_n1139_109# a_n1229_21# a_n1287_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X12 a_1969_n1009# a_1879_n1097# a_1821_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X13 a_n4839_n1009# a_n4929_n1097# a_n4987_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X14 a_637_n1009# a_547_n1097# a_489_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X15 a_n843_n1009# a_n933_n1097# a_n991_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X16 a_n3803_n1009# a_n3893_n1097# a_n3951_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X17 a_3153_n1009# a_3063_n1097# a_3005_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X18 a_n3655_n1009# a_n3745_n1097# a_n3803_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X19 a_n3951_109# a_n4041_21# a_n4099_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X20 a_3597_109# a_3507_21# a_3449_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X21 a_1377_109# a_1287_21# a_1229_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X22 a_3005_109# a_2915_21# a_2857_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X23 a_n2471_n1009# a_n2561_n1097# a_n2619_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X24 a_n4839_109# a_n4929_21# a_n4987_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X25 a_n2323_n1009# a_n2413_n1097# a_n2471_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X26 a_1229_109# a_1139_21# a_1081_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X27 a_n3211_109# a_n3301_21# a_n3359_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X28 a_n991_109# a_n1081_21# a_n1139_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X29 a_5077_109# a_4987_21# a_4929_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X30 a_n4395_n1009# a_n4485_n1097# a_n4543_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X31 a_n4247_n1009# a_n4337_n1097# a_n4395_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X32 a_n1879_109# a_n1969_21# a_n2027_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X33 a_1377_n1009# a_1287_n1097# a_1229_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X34 a_n1879_n1009# a_n1969_n1097# a_n2027_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X35 a_4041_n1009# a_3951_n1097# a_3893_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X36 a_n251_n1009# a_n341_n1097# a_n399_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X37 a_n695_109# a_n785_21# a_n843_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X38 a_1229_n1009# a_1139_n1097# a_1081_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X39 a_4929_109# a_4839_21# a_4781_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X40 a_n5283_109# a_n5373_21# a_n5431_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X41 a_3893_n1009# a_3803_n1097# a_3745_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X42 a_n3063_n1009# a_n3153_n1097# a_n3211_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X43 a_n4691_109# a_n4781_21# a_n4839_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X44 a_3301_109# a_3211_21# a_3153_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X45 a_45_109# a_n45_21# a_n103_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X46 a_n2915_n1009# a_n3005_n1097# a_n3063_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X47 a_n547_109# a_n637_21# a_n695_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X48 a_n5135_109# a_n5225_21# a_n5283_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X49 a_n4543_109# a_n4633_21# a_n4691_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X50 a_1969_109# a_1879_21# a_1821_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X51 a_n4987_n1009# a_n5077_n1097# a_n5135_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X52 a_785_109# a_695_21# a_637_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X53 a_4781_n1009# a_4691_n1097# a_4633_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X54 a_5373_109# a_5283_21# a_5225_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X55 a_1081_n1009# a_991_n1097# a_933_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X56 a_4633_n1009# a_4543_n1097# a_4485_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X57 a_933_n1009# a_843_n1097# a_785_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X58 a_4781_109# a_4691_21# a_4633_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X59 a_n2175_109# a_n2265_21# a_n2323_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X60 a_637_109# a_547_21# a_489_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X61 a_n1287_n1009# a_n1377_n1097# a_n1435_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X62 a_5225_109# a_5135_21# a_5077_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X63 a_n1583_109# a_n1673_21# a_n1731_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X64 a_n1139_n1009# a_n1229_n1097# a_n1287_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X65 a_3301_n1009# a_3211_n1097# a_3153_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X66 a_4633_109# a_4543_21# a_4485_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X67 a_n2027_109# a_n2117_21# a_n2175_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X68 a_4041_109# a_3951_21# a_3893_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X69 a_n1435_109# a_n1525_21# a_n1583_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X70 a_n399_n1009# a_n489_n1097# a_n547_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X71 a_n251_109# a_n341_21# a_n399_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X72 a_5373_n1009# a_5283_n1097# a_5225_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X73 a_2265_109# a_2175_21# a_2117_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X74 a_3893_109# a_3803_21# a_3745_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X75 a_1673_109# a_1583_21# a_1525_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X76 a_5225_n1009# a_5135_n1097# a_5077_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X77 a_n4099_109# a_n4189_21# a_n4247_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X78 a_2857_n1009# a_2767_n1097# a_2709_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X79 a_n4691_n1009# a_n4781_n1097# a_n4839_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X80 a_2709_n1009# a_2619_n1097# a_2561_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X81 a_n3507_109# a_n3597_21# a_n3655_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X82 a_2117_109# a_2027_21# a_1969_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X83 a_n4543_n1009# a_n4633_n1097# a_n4691_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X84 a_1673_n1009# a_1583_n1097# a_1525_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X85 a_341_n1009# a_251_n1097# a_193_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X86 a_1525_109# a_1435_21# a_1377_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X87 a_1525_n1009# a_1435_n1097# a_1377_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X88 a_193_n1009# a_103_n1097# a_45_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X89 a_341_109# a_251_21# a_193_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X90 a_n3359_109# a_n3449_21# a_n3507_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X91 a_n3211_n1009# a_n3301_n1097# a_n3359_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X92 a_n2767_109# a_n2857_21# a_n2915_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X93 a_4189_109# a_4099_21# a_4041_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X94 a_193_109# a_103_21# a_45_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X95 a_3449_n1009# a_3359_n1097# a_3301_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X96 a_n5283_n1009# a_n5373_n1097# a_n5431_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X97 a_n2619_109# a_n2709_21# a_n2767_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X98 a_2265_n1009# a_2175_n1097# a_2117_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X99 a_n5135_n1009# a_n5225_n1097# a_n5283_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X100 a_n2767_n1009# a_n2857_n1097# a_n2915_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X101 a_3449_109# a_3359_21# a_3301_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X102 a_n843_109# a_n933_21# a_n991_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X103 a_n5431_109# a_n5521_21# a_n5579_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X104 a_2117_n1009# a_2027_n1097# a_1969_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X105 a_n2619_n1009# a_n2709_n1097# a_n2767_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X106 a_n3951_n1009# a_n4041_n1097# a_n4099_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X107 a_2857_109# a_2767_21# a_2709_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X108 a_n1583_n1009# a_n1673_n1097# a_n1731_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X109 a_n1435_n1009# a_n1525_n1097# a_n1583_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X110 a_1081_109# a_991_21# a_933_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X111 a_4189_n1009# a_4099_n1097# a_4041_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X112 a_2709_109# a_2619_21# a_2561_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X113 a_n3063_109# a_n3153_21# a_n3211_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X114 a_489_n1009# a_399_n1097# a_341_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X115 a_n695_n1009# a_n785_n1097# a_n843_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X116 a_n2471_109# a_n2561_21# a_n2619_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X117 a_n547_n1009# a_n637_n1097# a_n695_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X118 a_933_109# a_843_21# a_785_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X119 a_n3507_n1009# a_n3597_n1097# a_n3655_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X120 a_5521_109# a_5431_21# a_5373_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X121 a_n2915_109# a_n3005_21# a_n3063_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X122 a_n3359_n1009# a_n3449_n1097# a_n3507_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X123 a_5521_n1009# a_5431_n1097# a_5373_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X124 a_n2323_109# a_n2413_21# a_n2471_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X125 a_3005_n1009# a_2915_n1097# a_2857_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X126 a_n2175_n1009# a_n2265_n1097# a_n2323_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X127 a_n1731_109# a_n1821_21# a_n1879_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X128 a_3153_109# a_3063_21# a_3005_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X129 a_n2027_n1009# a_n2117_n1097# a_n2175_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X130 a_1821_n1009# a_1731_n1097# a_1673_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X131 a_n991_n1009# a_n1081_n1097# a_n1139_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X132 a_n399_109# a_n489_21# a_n547_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X133 a_2561_109# a_2471_21# a_2413_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X134 a_n4987_109# a_n5077_21# a_n5135_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X135 a_5077_n1009# a_4987_n1097# a_4929_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X136 a_n4395_109# a_n4485_21# a_n4543_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X137 a_4929_n1009# a_4839_n1097# a_4781_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X138 a_n4099_n1009# a_n4189_n1097# a_n4247_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X139 a_n3803_109# a_n3893_21# a_n3951_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X140 a_2413_109# a_2323_21# a_2265_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X141 a_n103_n1009# a_n193_n1097# a_n251_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X142 a_1821_109# a_1731_21# a_1673_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X143 a_n4247_109# a_n4337_21# a_n4395_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X144 a_3745_n1009# a_3655_n1097# a_3597_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X145 a_3597_n1009# a_3507_n1097# a_3449_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X146 a_n3655_109# a_n3745_21# a_n3803_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X147 a_489_109# a_399_21# a_341_109# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X148 a_2561_n1009# a_2471_n1097# a_2413_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
X149 a_n5431_n1009# a_n5521_n1097# a_n5579_n1009# VSUBS sky130_fd_pr__nfet_01v8 w=4.5e+06u l=450000u
.ends


* Top level circuit opamp_v1

Xsky130_fd_pr__pfet_01v8_YT7TV5_0[0] vdd iref vss iref vout iref iref iref vout iref
+ iref vout vout vdd iref iref vout iref vdd iref vdd vdd vdd vout iref iref vout
+ vdd vout vdd vout iref iref vdd vout iref vdd vout vout iref vout iref iref vdd
+ vout vout iref vout iref iref vdd vout iref iref vdd iref vdd iref vout vdd iref
+ vdd iref vout iref vout iref vdd iref iref iref iref iref vdd iref vout vout iref
+ vout vdd vdd iref vdd vdd iref iref vout vout iref iref vdd iref vdd iref iref iref
+ vout iref vdd iref vdd vdd iref iref sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[1] vdd iref vss iref vout iref iref iref vout iref
+ iref vout vout vdd iref iref vout iref vdd iref vdd vdd vdd vout iref iref vout
+ vdd vout vdd vout iref iref vdd vout iref vdd vout vout iref vout iref iref vdd
+ vout vout iref vout iref iref vdd vout iref iref vdd iref vdd iref vout vdd iref
+ vdd iref vout iref vout iref vdd iref iref iref iref iref vdd iref vout vout iref
+ vout vdd vdd iref vdd vdd iref iref vout vout iref iref vdd iref vdd iref iref iref
+ vout iref vdd iref vdd vdd iref iref sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[2] vdd iref vss iref vout iref iref iref vout iref
+ iref vout vout vdd iref iref vout iref vdd iref vdd vdd vdd vout iref iref vout
+ vdd vout vdd vout iref iref vdd vout iref vdd vout vout iref vout iref iref vdd
+ vout vout iref vout iref iref vdd vout iref iref vdd iref vdd iref vout vdd iref
+ vdd iref vout iref vout iref vdd iref iref iref iref iref vdd iref vout vout iref
+ vout vdd vdd iref vdd vdd iref iref vout vout iref iref vdd iref vdd iref iref iref
+ vout iref vdd iref vdd vdd iref iref sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__nfet_01v8_8HUREQ_0 vss vbn vss vss vbn vbn vbn vss vbn vbn vbn vss
+ vss vbn vss vbn vbn vbn vbn vss vss vbn vbn vbn vbn vbn vss vbn vbn vbn vbn vbn
+ vbn vbn vbn vbn vss vbn vbn vbn vbn vss vbn vbn vss vbn vss vbn vbn vss vbn vbn
+ vbn vbn vbn vss vss vbn vss vbn vbn vbn vbn vbn sky130_fd_pr__nfet_01v8_8HUREQ
Xsky130_fd_pr__nfet_01v8_8HUREQ_1 vss vbn vss vss vbn vbn voe1 vss voe1 voe1 vbn vss
+ vss vbn vss vbn vbn vbn voe1 vss vss voe1 voe1 vbn vbn vbn vss vbn voe1 vbn voe1
+ voe1 vbn vbn vbn vbn vss vbn voe1 vbn vbn vss vbn voe1 vss voe1 vss voe1 vbn vss
+ vbn vbn voe1 voe1 vbn vss vss vbn vss vbn vbn vbn vbn voe1 sky130_fd_pr__nfet_01v8_8HUREQ
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_0 vss vout m3_11697_n3158# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_1 vss vout m3_11697_n3158# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_2 vss vout m3_11697_n3158# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__pfet_01v8_YC9MKB_1 vss vdd iref iref li_4703_1515# vdd li_4703_1515#
+ vdd iref li_4703_1515# vdd iref iref li_4703_1515# iref iref li_4703_1515# iref
+ vdd iref vdd vdd iref iref vdd iref li_4703_1515# iref iref vdd iref li_4703_1515#
+ li_4703_1515# sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__pfet_01v8_YC9MKB_0 vss vdd iref iref iref vdd iref vdd iref iref vdd
+ iref iref iref iref iref iref iref vdd iref vdd vdd iref iref vdd iref iref iref
+ iref vdd iref iref iref sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_3 vss vout m3_11697_n3158# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__pfet_01v8_YC9MKB_2 vss vdd iref iref li_4703_1515# vdd li_4703_1515#
+ vdd iref li_4703_1515# vdd iref iref li_4703_1515# iref iref li_4703_1515# iref
+ vdd iref vdd vdd iref iref vdd iref li_4703_1515# iref iref vdd iref li_4703_1515#
+ li_4703_1515# sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_4 vss vout m3_11697_n3158# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_5 vss vout m3_11697_n3158# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__nfet_01v8_THKFL3_0[0] vss voe1 vss m3_11697_n3158# sky130_fd_pr__nfet_01v8_THKFL3
Xsky130_fd_pr__nfet_01v8_THKFL3_0[1] vss voe1 vss m3_11697_n3158# sky130_fd_pr__nfet_01v8_THKFL3
Xsky130_fd_pr__pfet_01v8_YCMRKB_0 vin_p voe1 voe1 vss voe1 vin_p vin_p li_4703_1515#
+ li_4703_1515# vin_p vin_p vin_p vin_p vin_p li_4703_1515# vin_p vin_p li_4703_1515#
+ vin_p li_4703_1515# voe1 vin_p li_4703_1515# voe1 li_4703_1515# vin_p li_4703_1515#
+ vin_p li_4703_1515# voe1 voe1 voe1 vin_p vin_p vin_p li_4703_1515# vin_p vin_p voe1
+ voe1 vin_p voe1 vin_p vin_p vin_p voe1 vin_p vin_p vin_p li_4703_1515# vin_p vin_p
+ li_4703_1515# voe1 vin_p voe1 li_4703_1515# vin_p vin_p li_4703_1515# li_4703_1515#
+ vin_p vin_p li_4703_1515# li_4703_1515# li_4703_1515# vin_p vin_p vin_p li_4703_1515#
+ li_4703_1515# vin_p voe1 voe1 vin_p li_4703_1515# voe1 vin_p vin_p vin_p li_4703_1515#
+ vin_p voe1 li_4703_1515# vin_p li_4703_1515# voe1 vin_p vin_p vin_p li_4703_1515#
+ li_4703_1515# vin_p voe1 vin_p vin_p vin_p li_4703_1515# li_4703_1515# vin_p vin_p
+ vin_p voe1 voe1 vin_p voe1 li_4703_1515# vin_p vin_p voe1 vin_p li_4703_1515# vin_p
+ voe1 voe1 vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 li_4703_1515# voe1 voe1
+ voe1 vin_p vin_p li_4703_1515# voe1 voe1 vin_p vin_p vin_p li_4703_1515# li_4703_1515#
+ vin_p li_4703_1515# vin_p li_4703_1515# li_4703_1515# voe1 li_4703_1515# voe1 voe1
+ li_4703_1515# vin_p vin_p voe1 vin_p voe1 li_4703_1515# li_4703_1515# li_4703_1515#
+ li_4703_1515# vin_p vin_p voe1 li_4703_1515# voe1 vin_p vin_p voe1 vin_p voe1 vin_p
+ vin_p li_4703_1515# li_4703_1515# vin_p vin_p li_4703_1515# vin_p li_4703_1515#
+ voe1 vin_p voe1 li_4703_1515# li_4703_1515# vin_p voe1 li_4703_1515# vin_p vin_p
+ vin_p vin_p vin_p li_4703_1515# vin_p voe1 voe1 vin_p vin_p vin_p voe1 vin_p vin_p
+ vin_p voe1 voe1 vin_p li_4703_1515# vin_p sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__pfet_01v8_YCMRKB_1 vin_n vbn vbn vss vbn vin_n vin_n li_4703_1515#
+ li_4703_1515# vin_n vin_n vin_n vin_n vin_n li_4703_1515# vin_n vin_n li_4703_1515#
+ vin_n li_4703_1515# vbn vin_n li_4703_1515# vbn li_4703_1515# vin_n li_4703_1515#
+ vin_n li_4703_1515# vbn vbn vbn vin_n vin_n vin_n li_4703_1515# vin_n vin_n vbn
+ vbn vin_n vbn vin_n vin_n vin_n vbn vin_n vin_n vin_n li_4703_1515# vin_n vin_n
+ li_4703_1515# vbn vin_n vbn li_4703_1515# vin_n vin_n li_4703_1515# li_4703_1515#
+ vin_n vin_n li_4703_1515# li_4703_1515# li_4703_1515# vin_n vin_n vin_n li_4703_1515#
+ li_4703_1515# vin_n vbn vbn vin_n li_4703_1515# vbn vin_n vin_n vin_n li_4703_1515#
+ vin_n vbn li_4703_1515# vin_n li_4703_1515# vbn vin_n vin_n vin_n li_4703_1515#
+ li_4703_1515# vin_n vbn vin_n vin_n vin_n li_4703_1515# li_4703_1515# vin_n vin_n
+ vin_n vbn vbn vin_n vbn li_4703_1515# vin_n vin_n vbn vin_n li_4703_1515# vin_n
+ vbn vbn vin_n vin_n vin_n vbn vin_n vin_n vin_n vbn li_4703_1515# vbn vbn vbn vin_n
+ vin_n li_4703_1515# vbn vbn vin_n vin_n vin_n li_4703_1515# li_4703_1515# vin_n
+ li_4703_1515# vin_n li_4703_1515# li_4703_1515# vbn li_4703_1515# vbn vbn li_4703_1515#
+ vin_n vin_n vbn vin_n vbn li_4703_1515# li_4703_1515# li_4703_1515# li_4703_1515#
+ vin_n vin_n vbn li_4703_1515# vbn vin_n vin_n vbn vin_n vbn vin_n vin_n li_4703_1515#
+ li_4703_1515# vin_n vin_n li_4703_1515# vin_n li_4703_1515# vbn vin_n vbn li_4703_1515#
+ li_4703_1515# vin_n vbn li_4703_1515# vin_n vin_n vin_n vin_n vin_n li_4703_1515#
+ vin_n vbn vbn vin_n vin_n vin_n vbn vin_n vin_n vin_n vbn vbn vin_n li_4703_1515#
+ vin_n sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__pfet_01v8_YCMRKB_2 vin_n vbn vbn vss vbn vin_n vin_n li_4703_1515#
+ li_4703_1515# vin_n vin_n vin_n vin_n vin_n li_4703_1515# vin_n vin_n li_4703_1515#
+ vin_n li_4703_1515# vbn vin_n li_4703_1515# vbn li_4703_1515# vin_n li_4703_1515#
+ vin_n li_4703_1515# vbn vbn vbn vin_n vin_n vin_n li_4703_1515# vin_n vin_n vbn
+ vbn vin_n vbn vin_n vin_n vin_n vbn vin_n vin_n vin_n li_4703_1515# vin_n vin_n
+ li_4703_1515# vbn vin_n vbn li_4703_1515# vin_n vin_n li_4703_1515# li_4703_1515#
+ vin_n vin_n li_4703_1515# li_4703_1515# li_4703_1515# vin_n vin_n vin_n li_4703_1515#
+ li_4703_1515# vin_n vbn vbn vin_n li_4703_1515# vbn vin_n vin_n vin_n li_4703_1515#
+ vin_n vbn li_4703_1515# vin_n li_4703_1515# vbn vin_n vin_n vin_n li_4703_1515#
+ li_4703_1515# vin_n vbn vin_n vin_n vin_n li_4703_1515# li_4703_1515# vin_n vin_n
+ vin_n vbn vbn vin_n vbn li_4703_1515# vin_n vin_n vbn vin_n li_4703_1515# vin_n
+ vbn vbn vin_n vin_n vin_n vbn vin_n vin_n vin_n vbn li_4703_1515# vbn vbn vbn vin_n
+ vin_n li_4703_1515# vbn vbn vin_n vin_n vin_n li_4703_1515# li_4703_1515# vin_n
+ li_4703_1515# vin_n li_4703_1515# li_4703_1515# vbn li_4703_1515# vbn vbn li_4703_1515#
+ vin_n vin_n vbn vin_n vbn li_4703_1515# li_4703_1515# li_4703_1515# li_4703_1515#
+ vin_n vin_n vbn li_4703_1515# vbn vin_n vin_n vbn vin_n vbn vin_n vin_n li_4703_1515#
+ li_4703_1515# vin_n vin_n li_4703_1515# vin_n li_4703_1515# vbn vin_n vbn li_4703_1515#
+ li_4703_1515# vin_n vbn li_4703_1515# vin_n vin_n vin_n vin_n vin_n li_4703_1515#
+ vin_n vbn vbn vin_n vin_n vin_n vbn vin_n vin_n vin_n vbn vbn vin_n li_4703_1515#
+ vin_n sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__nfet_01v8_8JUMX6_0 voe1 vss voe1 voe1 voe1 voe1 vss voe1 vout vss vout
+ voe1 voe1 voe1 vout vout voe1 voe1 vout voe1 vss voe1 voe1 vout vout voe1 voe1 voe1
+ vout vss voe1 vout vout voe1 voe1 voe1 vss vss voe1 vss vout vout voe1 vout vss
+ voe1 voe1 vss voe1 voe1 vss vss vout vss vss voe1 voe1 vout vout voe1 voe1 voe1
+ voe1 voe1 vss vss voe1 vout voe1 vout voe1 vout voe1 voe1 voe1 vss vss voe1 voe1
+ vss vout vss voe1 voe1 voe1 vss vss vout vss voe1 vout vss vout vss vss voe1 voe1
+ vout voe1 vss vout voe1 voe1 vout vout voe1 voe1 voe1 vss vss vss vout voe1 vout
+ vss vout voe1 voe1 vout voe1 vss voe1 voe1 voe1 vout voe1 voe1 voe1 voe1 voe1 vss
+ voe1 vout voe1 vss voe1 voe1 voe1 voe1 voe1 voe1 vss vss vss voe1 voe1 voe1 voe1
+ voe1 vout voe1 voe1 voe1 vout vss voe1 voe1 voe1 voe1 vss voe1 vss voe1 voe1 vout
+ vout vout vss vout voe1 vout vss voe1 voe1 voe1 vss voe1 vout vss voe1 vout voe1
+ vss vout vout vss voe1 voe1 vss voe1 voe1 vout vout voe1 vss vss vout voe1 vss vss
+ voe1 vss vout voe1 voe1 vout voe1 vss vss vss voe1 voe1 vout vout vss vout voe1
+ vss vout vss voe1 vss vout vss voe1 vss vout vout vout vss vout voe1 voe1 vout vout
+ vss voe1 voe1 voe1 voe1 vss voe1 voe1 voe1 vout vout vout vout voe1 voe1 voe1 vss
+ vss voe1 vout voe1 voe1 voe1 voe1 voe1 vss voe1 vout voe1 vout voe1 vout voe1 voe1
+ vss voe1 voe1 vout voe1 vss voe1 vss voe1 voe1 vss vout voe1 vout voe1 voe1 vss
+ vss voe1 vout vss voe1 voe1 vss voe1 vout vout voe1 voe1 vss vout voe1 vout vss
+ sky130_fd_pr__nfet_01v8_8JUMX6
Xsky130_fd_pr__pfet_01v8_YCMRKB_3 vin_p voe1 voe1 vss voe1 vin_p vin_p li_4703_1515#
+ li_4703_1515# vin_p vin_p vin_p vin_p vin_p li_4703_1515# vin_p vin_p li_4703_1515#
+ vin_p li_4703_1515# voe1 vin_p li_4703_1515# voe1 li_4703_1515# vin_p li_4703_1515#
+ vin_p li_4703_1515# voe1 voe1 voe1 vin_p vin_p vin_p li_4703_1515# vin_p vin_p voe1
+ voe1 vin_p voe1 vin_p vin_p vin_p voe1 vin_p vin_p vin_p li_4703_1515# vin_p vin_p
+ li_4703_1515# voe1 vin_p voe1 li_4703_1515# vin_p vin_p li_4703_1515# li_4703_1515#
+ vin_p vin_p li_4703_1515# li_4703_1515# li_4703_1515# vin_p vin_p vin_p li_4703_1515#
+ li_4703_1515# vin_p voe1 voe1 vin_p li_4703_1515# voe1 vin_p vin_p vin_p li_4703_1515#
+ vin_p voe1 li_4703_1515# vin_p li_4703_1515# voe1 vin_p vin_p vin_p li_4703_1515#
+ li_4703_1515# vin_p voe1 vin_p vin_p vin_p li_4703_1515# li_4703_1515# vin_p vin_p
+ vin_p voe1 voe1 vin_p voe1 li_4703_1515# vin_p vin_p voe1 vin_p li_4703_1515# vin_p
+ voe1 voe1 vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 li_4703_1515# voe1 voe1
+ voe1 vin_p vin_p li_4703_1515# voe1 voe1 vin_p vin_p vin_p li_4703_1515# li_4703_1515#
+ vin_p li_4703_1515# vin_p li_4703_1515# li_4703_1515# voe1 li_4703_1515# voe1 voe1
+ li_4703_1515# vin_p vin_p voe1 vin_p voe1 li_4703_1515# li_4703_1515# li_4703_1515#
+ li_4703_1515# vin_p vin_p voe1 li_4703_1515# voe1 vin_p vin_p voe1 vin_p voe1 vin_p
+ vin_p li_4703_1515# li_4703_1515# vin_p vin_p li_4703_1515# vin_p li_4703_1515#
+ voe1 vin_p voe1 li_4703_1515# li_4703_1515# vin_p voe1 li_4703_1515# vin_p vin_p
+ vin_p vin_p vin_p li_4703_1515# vin_p voe1 voe1 vin_p vin_p vin_p voe1 vin_p vin_p
+ vin_p voe1 voe1 vin_p li_4703_1515# vin_p sky130_fd_pr__pfet_01v8_YCMRKB
.end

